��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P��v�"<ߞ��&'��k%P碶�R�ӣ�sĞ����tBtᆉi���5F�[��� JL�5�C2g] >�Qv'�{ɷ��2�͞��0�
��+��o)H#irw�����D�؀Lz}��#��}2�C�=\�>���aꥋ�Zv���_��1�0zvV���v��GJ���A	���p�sf���n{"v���Ҝ&K<�PG�e`_�#��`+�w=�)�6��h���s0�AT�!��%�����G�")l,��?��xp-z�Y��W0��7���t)|���9W %̦a"D�%�GTh�{m�P\�̂Ʋ��Dm �H��;Z{���ze�r��m�f$ԫ]M%���¢|����lAԙ!~�z���]w������x&o.aO�|��}���]MF��:����N4"{�һ��X`/i�F���d�[�.j���V�w1���E�aU�K�!IT��v��F���t�Ē��8zo=ߜH�Wk�*�SK�@�?��8���Ϗ�L�FJ���Էt�kgC:zkV�'��~�-5�z�{�e���V�UHf�����tެh�I[�k	������~�R�[�jC<�KӅ]0�G�Yjwb!���Q��tIj�6�C
rcO.�����KR�7`f��L�=p4�$.z���,�P8��>��v��ｫF\��hM�5e0^O�V�&��/J�o����p�ސ��O�������)ϨN>;:_.���e�<W����)ϋ��EW�/˝@&͙g3@�H�;��P��m���oۍ���F@�N�B�M�{1�s�"_F���e�En������/Q�H�4n����e~m�h����;�XO�nH2G��ď�p�A\5f�f���e��<�4�ݝg��#L�V_wq`��FR)�OM���8F�}��>ғ!�e�8РsN`����PA�eђ���vʁ�� 3i�v�X�H֎�����J=��Va��-���m@�z�������(������gnQ�����(���8)�!�T���s��mٕ��&��qki�z�})#���>��'Z���d�7-P�I?~Zu��]2w՟�7��̶S�WOv��$?�.&����ac�Σ\����	Q��qC$ �I-��jI\��27ү	�5gԣ=^n�Jy��M��X#��6��u����+h���/�-�i�L����kg�7�qhv֧Ti_��~��΅����k��?7�z]�`^�+PX]��	-��3�]�.X�[���(�W�}<����Pr��k�]M��:�����wb�y;?��n�o��`h���ֆ�&gm�刟6f#�0T�$X���ym�3|=J"���\�
\�X@��:{���BH��-�� Ô���N���q��"�f~?
�h���畩��=���F�;����4�4{�����3�"�;�qv��B@oB���h
�j�H(�8�`�T/�LQzkڵ�k�j������`�8m�)J�j<ϴ^���K�-/��/�(��N�t�7��Sw�K�3e?�:��}`d_���;�3�B���VN`��^���Ap�h&�K��+��E��-QbXo�j]?x^[f2���Q��j%a�<װ.MߖR��\h!�ha�k��+6}_y�d�C W�q<-/Ö�Ġȑ������X�I�#~`��}q?�A��Gb ��v�餒�����k$�u��o�a�CS���˄��Q�_��#�ADLD��H��'��_�/nِ���X�<�*��P��ksu2�D���:�	�!!��C�*E�����'�fc�{���r =�v��TR�21ó�/'(�AЋ�/o��a�@9���&Na���h�������QH)��}!�yo����H��b{�UJ�,9���O�it>�����e��<��g��JXaHf���+�]�"P�d���m�}M����I����n '-��Գ;Kt����~�H�_$y5E7�j`���L�X������
(m狱��f�^a���F�w|�2/̡�a�y���[�2C{P���
j�?�TI����3�s�~�kz�i/��K,s�j !.�_����s����O�@Uf>T�Ok�1l��T�ay�MA����X�ɤ�@x�K��5r����1q��ϊ��� Ex��9�����:�~�+(�¢��w;D��"PYO�v`NĻzF�P�CAe��ꁼ��]i(3�n6�C�$<kĪ18S��l!�v��j��=6���v��KǕl� ĵ*+p)"A�^~}� W������窓���(*��	X��*w�t�#���>V��h+I 2[|ZT�O���R-z���OR-��{�hp�k�����~*�. �����9\�m�� ��@k*	L��<#c��˷�%��sIe���@�'>!��o��
_�G�_���p��fx)�;$���y�r�g�iVk�Śf ���˟�=��_X��AFvy�u�ش�q`���AF(M*����8�-������A�ʧ&�)��N.s8s�d����CW�Nlk�7dz���V}'���cS�nE��,�� E<
���9-�@J�z����QU=ծ|��N�K�C"L�J�&�nUׄ�Ӗ��/A������,PH��[�h�h˦�DG��3U��V�X>�@\�N�!ya�����������^F�"��\�&��5�I��2V�*���%�n���Ԟ��XE�R۠=@�M7lz�a?�P[2{��u��ԗ,6�7�GQ��z�����Ŭ\��D��ɝczp���WyG���r����l�m3b�֟TJ�'�GU�F���d�~��3� ��������\�2w{M�n�\Z;'�צm����A9"����n�k��i ��r >ş#�V���m���-a5-W@㾹)�d��m�z��Օ�rd��ҷ�C�YĎѲ)�Wte�g�M��g5Hu
��&�}�n���<��6���a�J�Ҿ܅vg��4���c�X�돝�ͱ���A�)����^�\�Ջ�%Iy��}0j�X<�rt��P ]�٨V�H��5�keU��tz�����@�1V��>w�����W�� �[kϸɫ_�3��ܤ�D���!9�@?(�-��0�'�n,/�9Q��-y�_�W�ѽ�r����۵�#,Pǫ=͠S��}�)�W�� 2#��m�����g��Ӱ�ux3��紪	�o�
�G)���K��Q�W�U�<��A� Y��:M�Adk�BAΣ�������4M���只o�1b�Y&�pF�T�|��%�ӟx�eM�/��L�����h굀���R?�aĴp��q���R<g����jud� ���BC��
�C��r���`� �#��K3֌`rFg��\��(.���o!p�Ri��x�O�~��� ��k�rk��Ƒ�����M[߬@R�6��z�P3�Z�����O��0��A㠌���_������T���� �� 뙺�*�v$��&�3{�h���8�p���_���l���Û�;,u��;X�����zϣW�:����k8�$�jq5=zVv,'�~�+*�Ԁ������4$X�E�Kݕ0v�4����ms٫(��o�lQ%x�ک�m�� ����H�:Q��E�1EH���ֹ9G����և�_��%R}
�Vj
�_�BsGs��i�D0%࣡��>ِ��t����m�/�i�h��;+��Ji�c�P���2N9@DfW���hֆ��:����Z������7��dLE +`>Dg`��B_\>���Z6�\��ｵh\����LI�ۙ~?��(�-����	�
�=&��<y.�T蠕���A9B�j�rqT|�M"Y]	#%�
!�p_��%G�/���.Ե'����PZ�P��=���|F.�μst��X�$��t�I�k�D� u<�>r˵:��׭a��Ό���EqNa&�p�[����7�-ճ�p%�d�iT��s��`�m��*s�^eP��Z� ����9֎������w0[��fm� ��@�FIFYϢ)z��;�"�H���0q�i",-ucA^�B"�#�jzA��R��<����(�Y�\�_ �N;ϲ�j���+��,���ӆ���ߏI�_\�'e�;~�̽�m��ۆ���1?k0�9��(����O�;2.iQ��?��=�fU�g��{��9���5E5;AB�D5G���\ -ZBsр|��7�3��o/n�}~B(�80[Y�R��(�8��܁)~r�,e
'����\W,�sg���:w�ӻjT�awYm[M_Ϭ!c��*���|$����>����R٠s��d&*4����Ak�v�I΋�Up��۠7ژ�"��H�[/e�PS?k�GPǳ��`�B�^��|���������cl�g���WlKN�FR��	D��"�� �	����� �W�SKpXd��PaM�A$M��=K�b��
���4i�?���G�k�S@�Ͼ/?�}���O܍�r���Pz{�i����\�w�����&���y�生����b�z5hj�X�zE���g�o����g��� K)C�o?��LΑu�ζz�������|�����x �4f\� �묽�#U����fH�_M��q:q�ؘK�?*k�B�:���'v������l�A硇���j��Q$Z1.�_��c8� L�Y���OꞛLV�Ӆ%���8Qu�~{�^�_�v�����Z�<�7���8��^�%B�FkI0���Y��&�)HNX�^`��&N�m��<���
�̾��wv�`6}��ui����f��ˠu�d��
��$K���:��o>fJ:o:��MOoT���`��W�i��_��{95�Ve&�cx"Q�U����W��eKOT���l1��.�H�o甄/����13x��)�&?�K�#s=���R������5T�0�Ն�쿙 -���	#%����[�d�z
O�a��W:pU{�߆ ^���;_��O�{�S85�-F�qu�>�֡5r�}V`�?�j���߯���.��/o�g���i*25 ��[��$]*Z��'���֡`��˅ަ����!P��]��c�<��-x��#E��_����V��e�f�Ɛ�
RH�{Y8L7rb�P��e�3�?�ߋ��Ϙk�U}����`%���WR��2�:8 ��G<���������9�]�<+�	�PU |;VH����������t��[�P)ŵ�-bjNH�q&$s��Q�ϕ�D��3
�aN��=�����M����:��[k�'ִ!��E�;������0!��4Gߔ� r�%���o�o�U߈~��7߱
������z�I�[��o�;I����y�����@�@��\����@R)�t1�� F�1�y����U�)]b���(҃]���y�t�8�i[Z�&�r�LX��FV"�Q����Q�XUQ�0{�p��B�y��7�*2�t���M����IY{��yJ�
��t/��T
K�_�л��3K=x���S�W�W�������g���Xj�ܹq����޿^�1���S���c��Ȅg���<����uC��A���6������U߉L�z���ÿvm�K�֎F�mg���b���]~f����z��u��54N?��c�خ���:;9��������ſ��������@*X����f����sS��+�21yF�^��4~۸�=��
F<T�}0m�j�}{E���!�*@�O*��e�'A�9F|��66��\8ˑ��"�F�F'��J��և�A�"��E+`�М�*Pk�c%��y�8��?��9�z%E��,IwgƆ��@�ش<���|��4:�:�ͻԉd�S1m�)������ΐ��na����q����ߖ<����� x��[�?^�_�[��`���̊����0d2kW��yU �l�'}1��Da�Rq�di3�	�&N�Q񊐷h�'�<�1ii�Gm�Qc���*e3�l�Ͳ�>(s$��s�<�,z ����2f����!*f;j�}��	�\��-��$�l�Q�L�N�yF /'��(2[u��\&Vt[�A@���F���K�PX`5ɃF����y�6�Z�p��p���Y�{�����瓎'W�0�q]䠗Vt����������q
����?�Գy����2_OM�H{5z@U�߹;b�5�j�i� b�A9�u@�jX�rh�����}�ۙt v��`����!�=�����X��K%�v>�UzE�5�����D�Rs;�������������=U��/z@r�o|�"�l}�Jw�Ԫ�25~ʕcL�����]���}���1��೶�s��H���g�%�$B�B?� mXZ!���,R�8K��b�6k����Gn�����j�F}�g�� P�^8ڄ0\Xv���\^DۃsX@|�����}�h_�?���<C��O�T���6>�s.?m����KD|Ul�f����%9�n�"���rFC�h2�+Pn�|�4?���~�.���AO�&p�W�V��S������X��;�M���_���'����*���㰥��1?j.X5#��&�J�C_�L��kU�NG��$c��i-�U/	쇰i�"F`w&Q������r�
������G�|�c2=��ւ��!�N�v�a���,�8�0��=[�C�ł�E3s�� 9�A�t�o�/��<Q��uN.���;c��EGx�O��#��"�������Sp���c�Z�Pײl�)��q�錕���a�M.Q%��Z@s�ѢDd�@�MhZ�k8��0�{T:R�����_ZNW*
�HM
ܲ����K��IWQ�:Y	6�&�)�|��C�8���y&(^?
����˵M}����8,b��^�h\���!��)��S�'�]��o�kՀFN0�C�M�_3X�<���P�����\��Ee$���I����DI����B������������,)�M��%0�V���o/�C��_V>8���|���|���g�o��^���{�Q�B6y,��݆ rA��DY�p㯫p�)L�D�˄�M#{�2g�[�F�b��T���
�E=�'IINv��׫WL0}�th � 2ML����M��9P��EH��es���?����Yy�Z�ݏ_���9���ƌ�w�kq���"�bu��p��5�cΝ7���ja���č�@����y�����)o�m��C�r�|qm5I�l��Nh0�`�IPhe�6������;i�KN�21�.�G/e�M�s)%���X)�����aE�8�n{���\��0C����2�YЈc����� ���[1/:l�r�&�q�vN赙��O�+��}�� ɮ+���g5�N�Mƽ�e�
Վ��q~^p�Ǖ��ǸQ�X%���+�l����}��`�U8E�kh&p��5��ޘZ�Ӟ4V��nt������D݄���ϟs����]�M��oa>�dGə����0�%��;WB7��n`mV7	�5�Y]�������SI��	�1:�y咔�uK5���:��+m�#a����rH�i�b�魀2T��&�{;���G�Bc&Y�Sx��3q�
���ӡ�;�*<�d���%U�N��+"�W��pj�����F���V��j��������K�'�z��W~ϴm��ƞ��?^�v�h�Yפ����\�1%��ґiN9���8a��QE_I�y]�"w�i=�
#e�g�֌�~�_�}�.ᦈ��8�ɳa��x�v������������F)�"�VM �n�o�I�����$�gZe�`,G���ce��+�����sE��o9�x5c�*���?UQ�ڏ8��
�K�k��$���gr/�$�}��O.��X4S%�����"�j|P����v�ܺRI����t]6��ER&�T��qj0�|�\����I`(S��4ZR�#S�˯�V��h�`��Y��ˣ�̸��Q�Z�3I?ukN(W���y�BLw�/^s�?F*<cO��1 ����Z�S�b����%?�/��K��ѲPV�IL�NǎW��#���X�e�j���a�0�Edɋ��;h5Rq���Zf�����隔P�@�����#:��y�~�����pa��"8v�m=�2��8���fa ����'�
�+�,KGA���� &��V�N���a��Nst�j�~5/T�v��/Yw�%��I*3�� ��pG�S���D��ٛ��U(߇��U�}2�����X�:�d��3����]U��40�}��vV���M%/�%hjk��LHH����rqsm�D8%Z&G@����e�vVf2�2k�uq�Okl�0� \��,yv.���p�7%(��Y�m&�3��� ]�I��}ra4'�;�����6�P���K�x并���F/� e�l��jd�	�e�|��q	i�s�����Z���
��Am���9���^�^Y�����R�{��@��Ow�S#��p5��9
H���faSjO0�ry������rCw@3�B7�5���X��]�k�y�����Otzn=el[^��^z�o.K0��f�([����Ӥ(�\Kn���jӄAN�6�MP����*�1�!���(�r�d�:�rwy����-4����tE�KD,Oqh뚣\�qB�Ԗ}�p�K�Q���J�6��hn��{O�+�����������u3!�[�3x[��O����r��Vعy�h#��ۇ�.�.����x������! �Ι�t�D]�~SFr�D���:n�������AJ;�0��� �Qm��-K&�*W3����s�e�D��D6|%�}�F��V�r���3<d�uq �f^����{m����Ompt?��"�|^W�`/�z�Έ�3�..���'�����j٨i�o:�Pi���I���$]wG�-'o���Lw�&P����Gy�K�\�I�T���i!@�b�D�_ē<7
U�V��Z�2ۃ�����?^�N��^�d��j@�8�&���V�|:���.��n�����(lX��\F��jM�]oW�b�s�#C��s��ʮ�CÃ�K��a(�:�p�M���O�^��o����އ�9=nn��-\y<I�6y�� �v��ԥ����%��h��o�R�iI(d~�)4*i�VЎ	)��U��<Z˹�Ҩ�T������3G�����g�0Dm���e�� �t�`|�H����(���D�Y�E�O���۔?��%'�~����O
g0{�x����|%���u�/Yh�ehX
g����V1��-�Mv�}ob�	���y�N�)1r\9>I��CԦA";��
i��4�� �-�|-����0�|���i��ioDϝ�t��������D��|��r�8>��"��|�r��~m��?f�(M��ĒĊ��rɍc����[�Г|��\��������_��V��)^ݴצur��k������˩����x�7�}�/ؠ�]	l�#��t�.Zy=E�G4 G	�ؠ-�LA�l,�y��*hc��S�Fx�pĲ0��d�lD���|�a@<w��#�g����jvU����O!���_��?�m��
��Y&G���"��`\���S��fQ�<���敏���zt~��V6��V?0aш���L�����\�S�M�i��T���Oa}0h���#s�t���;u�.yC��qQx�_�"]OX���u�4й��w�=j7\#��V�jY"j�����K|�f�c<N�d`U7:�p�:����m�)A���s��I����ݪPB�5H�[e��Y����i[e�|,t��kMNW[3�߁&�Ov�F�C��p�;�.��~�(H��I��Z$���2L{ڦ4��ޅ;�F�M��F�ZHϯ��,VvA�_���t�'��.���IS�����Ñ���˱�8��"�v�3S���*�, Lk
��yYz ���z�\�ton���#����w��P�� ��h��0\������9���0�]��J�I�؀��܏��R�"�����YR��}Ko俯��O �pʉ?���]Mzz�?�	�=��$Xu8xe�.��=H����������4���Gra?Y|h�u���U�@���k��^�
M��^��`}��de�'���ӡ�/8g�n�7M��_���sv&1`��v�����#��F[�b0�����+b��ʱ��֬x�r��צ�o\������K�|/��ex%�}a֠��X��bF́�ʹ�b��17 �xK�����a
�G3 B�IH�8G� �)�iK.��?�Y��D��=��A�zb|OѺF���KAȳk��뷣� '���2XqO��T�lgn����A������'�﵁-.���Q����5��"ȤT#��Bȶ��zQ(�����{�6B��ǘ�P7x��P_�'&�f�,GzlRC���N@�7����p����3֑mm�m�:�@g���ڙ�A�s氉�z?�;���h�����$0T���,;���	�#e«o1�m���3�������hP�4,�	r��F\hܤ�&}��Q�w����޾|2��=��/�8)+�\�{�傱��	��&����iST;G�	��	�ݓkߞ�!(^���,G���N���Hb���� �}�V���fZ(z%�GE�m�yG�� ����2�4����:��.ϡ�Ğ�����3�yN]&�>�j��92�o�&j�ca�	��@���O^ȸ������ ��^��}J�� Ŝ|���;4���&�:�  �r�'�����I����,U��ag6�h��E�~*#��q_�d+�s
Ч�6��?�JAQ�Ȇ�X����٢��>H�Eه�~�ݏ����ժt �4��Cć��'�'-Km�w�zW۹Kn�F��ol��iB	�(X��"�H��\
�}�6�T�(k �9h(�>�*I:w9ߥG@����
e*�VJ1G�f�ci�#�;�׾�/�;��Z�E��2�nK}=iU�~U�*�7��+���_R�'�Y>�^��3M����Lbo6Yk��=�w����q�g#���]\���>N�G�;���u~&����"������|���;Vf|z*>�NyCOD�6��]��� ��$����F͍j��c?JZA�0s�B�GŊ˘D4��2���U���N$�����H�S��S��4:����f���7}��#� &啂h[��D���xÔ�'���O�����1����s��Mq�Л����c	�^��/k��˿�؟�L�ڞx�LĲ#�������+u��y��`�M[�>��dR��� ��-��#�&蚨�x�y|X(Z�ج�5R��b�~�4DA�	_���K|�r><�}�������z[� 6Õc��r�a9�	�6P�mVE�Fu��t���/�v "]2��0�������y�"��d��	��q,��HlnF�ԥ���*������ScK�(����ؾ+�H���ٺ�-��hQV/:W���~H���N��?������)S��W�鈃%���H�"`�,S����'����R��M���xl�EqWN����F�ҏ�?��GJ�\8�#~���e��4�:����3�Y%��]������^%'�B�H�􇩗�����D[���v{6}�6�v���z 3�E�c�O��Z|�����cr�n� m���sb�.wJ�0��s2�o9��i����,�'(_�~n���Q�}^�yy�@�P%iM��U������5�>���z	 E\���z�T�Z�s_a#��ҁs2��.Uz��l�m��<:h�a�S�pZ�-�>�/)�{:�9��i=�Ӟ�ߝ�C��bۿ�E|%뎗\�? "L�o��x\���2
) �~T�����Y��Px���|Ga�jW��dk��F�j]>^� ���U�>�f�h^
`�D�~��*E�=�����f|ޕq��p�7ݥ �3q}Oո�~�PL��s���5<z��_��>���4Y�-̾�ۨѵ�JCD�G�p�m�B��GM�N8�S�>x�	C���+`ϫ`��Q�_����ㄬFC�4.¥�A��!(��}�v��ߝ��u�<�Q4}}c1�g����cq���c�fG��|_��Y�c��	��"�۸ �� �0_2�T�~.�g��'���ڣ��7���s���QWN�#��^��O���r2����[�ǖ�W������M|�2��b��8���l4rP���`N���x&�#�������c��Ew��D��c����,7(�x`���V����IrOH�mc�ᬍCB�������~���y����� ?��&)|�ܗ`AH�])$�@�хc>��v���k�'b���e�,M��=�.<���>���5�?5O�`;�.�T�,OQ6c󎪗|�|aԙ�Z�	���Ï��T�;�p�N��О�Ql7�&Ы���/\��#�����n�2�4��&~��;V���V�u?x=s�DC|�UkzW��kn�������u:1�M�_c<�?�0@3ܳ+BH�=M"&����1qɨy��/|wW�p����-���'�B�x}��3;h�TAq����O'�uBwCb�D!�V	�4�S��iM|�3�C3N���ߘ���{	q'*�Z�V�ժ��a)!�+�I���b�7��/�+�;���͌Y\Г-:�Mm���@Oa�	ɰ��|��%2o�!�éB�&�0���w��B-|s�!ٓ��eB����g�kF�(��@�
�W���I_���b������Xzb�h���p���U4���})���V�n�,v �8 ��6 GݸX����	�n=B�������
%Rˢ�&���.�H�=�^����Ɍu58o��`�_{�o�Gy�P�0:� S�����y|�ڭI3fv�r^�"M��ñn��g6�G�5,���]������l��vjU*�m35Q����:�_����D5}N6�o���c&A#+:�`�|]㗉��  }Bp�0�h�[���)�ZJ�@V���1���LUlȤ��%���C7ݰc6�Y4��'w��ZTwgN�i�*���jc��Q�|(!;����0��|��K�ߕ� P�R�e����,&�@n�G7��F���q~7Ę����&ؒ��jE"]��:渢���1S_8��K���o��y���NU~��������4���������|� K
��n� �,�S�P��S�I�ږPS�_�g��a���,��y*� s]�՟�S\ƒx�����p�HP�}f���έ,�g�6"��L��rG�WT�А��/����E?B2�b�o��(�Yb�Ȑ��5���YM�E|�t灲Ec��l����U�DF������˚+�N�A�ĸ�FLP&N�i�w����d�Q Ç9�OQ�SjF`���5MX�Y�SH��uo}�b)�����_��z�*��W����0��!
G�V�ӿ�[%��Twd��&��o��i�M͵l~, �i7iq�L�_����������(��H%'���+]�;�¢�J�Мv�C@�.�4�>�915H��7ɍ\ ��B�VL�L�5�VJ�8��\a��}JYtp.��߲Tr[fՒ(���]X 2��c2�	[s~�[�_n�ӻU��q�K�Q��$�b��7��8C���
�_B볥I������4ZI:����3^��|�{c�F�<��m ����}�ce�N�zoU�^J
�n�W*��{�������q˲|;���z.(G/k(����酡O����P��n�e��Z3��-��:\?���/��t�C�POa�t�W�d���q���A� ]��N�?S4�c^5@��ؗ+>:a�*��x�M��c|{T��}N��s[*GB���Lp��K��=&U�O˜K���?��@�� ���`������5pI�kx=}cL�+2~����p����a�Y�ξ���ax��p�~��f(V��8g�^a���	-�Pz�̘j>�
��X�w�aơ?l�TF��.]�Y�5�-t޻.���?�9myl����y.MB�
����s�%ml �fDL�"���O,�7��>1�5P��dA���T�����ΦB�狭KU�Vn���8�Й���ίbV��� �:*�lV����M��8$�R�`ӗO��+�CxH�,σ�����}�J��oש��ƾ	_�(�
�>%�;>,�x	�#lq#N�� OӰk�ZND݂p��%��IZs%�u�In���s����yz�LJ� �P1�g�i$���7�߻n�à��?�#E.H�w@�̫���Wg�(#s*��w����)��?�*�x	%MA�2����>�k0[�'��ɯfDH	E��+��	���ȁ��}��,�jFW�fd�'�=-H�BELM�[!al@"���]�C����=��rl����u\�fԈ��	��sM.��P��_�/�ש�K}�~ܺV������,��+)\���-r�1E�=�w�0�i��'&����[�@�r]���4F��~�!y�
@m�q����K��K�=�${ش����X���=H�>����=tX�L�YQ����,��P�ؑuI���43����a	c�Y �Bl�2_��C�gK�+o iB��1&�6��a����;s.#S���ػ���Es@�yI�'�q!,�Eb�0��jT_��Nk�zh��ȿ���͂�Z?�Uz�n�� �?i_�.8�.}{�ީC�vl�Ã�FiWh�%I��n�݊�X̡Ђ��.�f�c�C����(����=lY��
�`@̂�<��ۊ����4s	��hE�[�p��vّ��
����?����b_o$�M�m�!��Ȩ�?�sFg�V���˯�=qaXL��vVd�å���k�+�E@K��.W9��@��g?��~�O3�9T�֊&����ϐ���
ܿ��H�_�X�o��g�]�-)/J7�O%��A%�tg5��kU��^�߀��`
��:<7>}��4�#}���(=Hn��Y�j��������ʻcoW�O���c�i�'=�=��}
��_-v�¥ڵ���~G\[p���h��ʕeA$i�ܾ�D�@�ف�	�j3,�[T�A�Zs����!CY���t���
L�2�_&g�hf��+DV�X���>��,`�1�~���<��R�h����-�e�q����P��r���jo��W߼T��Vh	���;��<*�/�Y��l��wqRB�ç��XI_����]S�]��Fh�4E-'V����Ƙ�͚x?�/���筹 R��m��X���p�C[_��X<��	�7�^;�[uR(��~UhIȘlƻ<��ꓠ��5d��JVW��}�}�52����͑.���v<��x�[an`Q��[b�7XܥW��K�7��#�¬����Ɇ��uX��@<Xm~�ӂ
�֞�a}�O��p.�r
C\�-h������@Ĩ�آ��A� �jmB�|�UK�O��^��V��A�P�
F���i����m���w^�p�TLip�k��}�f�4��E�880�R�Y�x��cq�`�z���(4��9�|/��y7RG%�\�w���Z;�(� =q^x�_ԇ�;���!g�
ݐ�\��K��s=1� ^�:�!���dY���A�^�D���q�m�����k^mW�aI_�x�2_��N蔍��h���ρݥ�0���6V��V@�D�P#q��.J|w����}���К� �o�A�|���� ������r�k/��t"!"c<�-����#0f�,ߜ���8�ע�Љe��臆�v1�'�$�b
(��*@���zo�0uS[RfR�ȳ=C�B�m�0-xssx(=��ѷ�B�JGfPH�S�<�c6QY˚�Y�;�������|r�����5p'Y��g�kkOԶY(�ڜ�"�*:�[�U�]Q}� k�b1i/�\הv�P!��<���G���0j�w&�[A?�'BT���	��uᏐӊ�JU��'�/�x�+�)��WPdu��D5-��(#�Mn���6G����B���h�D�L�o
��MX���#,�����j@ �p2v�\+�_~I�UsB��Z<�}`�Tc�Q�W�X�������S'ZE�����*O�$�&� �d��������zr�� �m� ����T��q��p��]�&͇	����eAw�S|ݻ�u4�����
�J�Qx����5�Ι.�X'-�p!�ԁ�lYJ�,�>E��} �6=`p���,�-�
ӈ9~�Sh��I�l��Raf� �A�*�7`��*����9;w}�f;o�ў�۔����L�	Bz&	���l�����kB@�k�t³́lQ'.�4�))�O�;Gni�UG�ڽ�n��Z^N��^�{��>Q�2���C�4�Q�,xv�l�h"�$c��ӕ��N͠Z�/�ls���H�T�\.�1)��>���W�W�a� AIZ���7�?wϋ�v��Ǌ�wf�CU&�_�X�9 ���}q�%ep."7�pis;ט�^��H����-3G�O��n��ᢷ0Kf�B�_�6AKWA�[�o����TX��m7�������&�)���P1�?b�9L���;��0N���z~� ��=|v:��!f�#t�Zާ�b�3d
�1�tWL�bv��h���g$�p��i�k@:�Q0;�����I�,�)�Tf���>��P$�M����4z|~K��td<m�Vxp5�LWhxk���m�J�4��Pe]�T��ﴬ��y�m%�ji>��A��0s+�PA�y6.�?BS��E�FD��Yt'�)&g	敇)��'�F9��]��C�������%�&p���2��^�܌4�H�b�I� d{��5m2F�ߓ(��p�x7�R�}@�:a���fg�'����y�����1�;J��[��1Թ��%����LBz]e��+���R��ONҹӜ�!�xw�8&�¢�TY}H�V ��Q�� �1/T99~��=�Ƭ����smn�	%%|����x�y��v So�����bu��bb�&��b���FMI���>��Fx�ă5��`,ΰcYdJ���?�i0�߰��]��`�\�6���X�2\����%2��i�P��T���h�JH�2c���*w��F)B"�"�_T+��=�0w��=�5xa�ٞ���_P0�b�~d<y|�i�'����3���~����k2K�vח!���"jT��=��_�H+L:y����-�隆��*8]���=o��m��44��Zh�<tOb��a���e��(+��vI���ww��k4�����S�r?k�O�m46	��]�I��}�?�0_��D�/x\Mv�v���G��iթ�`�k�xt��;�Z�۵z�3��;ɜ����<R��>������4+N`�׋�������=��3,��e��$�#!ѬZ,b�ߍ�Ǖ�tV��=u
�V 4��nx�������#��-��*=�̥�h@�A�#���[��4���u��3������;�5����UW�R��P
q�(��+���3�c�$v�[��z3;v��T7Y�O�8��˿�nnu��7�2y ��'�?�񇩝����}�w)�*�*��mȓ'�@l�L����>��l�%�j8�6t/-�����?9�s��iH�qsim���T/��t�S�-��K�`����J���駌U��� �f��1�;T�&���-�V\��**��}�Z��V�
��@7�O��nw�}l����ް���=Kw�s@5W�'������|���o�Uw���-�dл���r��Y�@�)��J�_���7�cB�����~ǲ�	��w�Ex���y<>��)yFT��њY_�=�S�J���w���M�,H����4J��r�f]$u��8�L7��O�I���st��u�m7�<�c�~ֹv	��cL�(��Aϟ���":�^�@��_[��A��D�"X���0��A���H�j���H�~G�3)�tLvQ�w��?��j���`�uJ@(�Qe�N3�Ll��+�\ ��y�*9�v��d����$*d���S1�Ʒ���5}�s�Ǝje�����y�ɏ�[q�N�3`��	��wluS�J�.N�}A��OU���%��k��g;yۣ|��ߍw{&���Q�g_�.=�a������u]����"�"�[ʛ���K���H�ԊTR��V]b6�/ ��h8��[�S�Ez�%Ϧ�s�n�9Ì
�I�h􊅞ٍLw��FqA�x�o�F�l+�/2��J�i�M�9��kv��E�']W ]@�����+Q��b�N��XF���0�-����'nE���(v�p���7�����B�[�9��J`WQ�61�C݀�h<�nKƹ�V�͊g�QL '
xo��#Q��=E�=1���Yx́�il��ߍ�аQTR>{�qf�A�)A�G$�n�Ů5�p&�7��g�*0]�t"l��f޳�i(i3��ޣ��^&/��jM���H��@����oߧ,���M�Ќ$�j�7���&��t��P��S&��B�(^�N�@ �nfU�P0�[�q���P��%�p�Fx㈁l7AF����xL4�?�#�n�Ŋ�_�˲�
���ܜ7Y��9��Z�e����w]T�f������`J�f�ѓ��6�<RE 6)����_�T�N�l�<&]�'̊c;���șM�b�9jx����fi����ͦ&5��`L��4�3tBB2.T�	 �M8�m�������h�[���(�Q*�����W����#p\|_0�����=C�Ө#��T�,�a^&]b��0��P���y�,�^AjYȌ=n�ج;�W܂M�:�B��G���٫�U1��5�?�R��A�IZq���
(}$��^��b����{�,?'�'1�x�ނ1��τ�b |�Zun�y	�\���"2�Ȟ~���NRag�h���IքW�ҶNt�B�L��x^�U���Y.�v�5ma_�UfB�GN�PR�G�������ht�LU9`V�x;XY`k�ɏޜ<��ʲ��E�wa�sx�uR%�f�w��O���Σ!�g�!e8|�+N5*T!K�~{5P(D�\��� 0�o��A�2hiK�f)������惷gH�|8IB��O.�z�x%�Z�/�FH���'��:��\<j>,Hyn��#4d���r�g	t�ĽC֕��^�i#/�&�_n5��߄1�4���}�%�C.�4K')tKI#$�~���1v�F*�Z \��W:rtd��=�cJߤB/�=f�2q����H�2�2��J`͓=%[w6g���lLK�A��S�''���h������I{vt5���]���[� ��3vP,=�]'*M͝ԷU�]b���/���XGoq6{�p={w������(r��X֟ �}���8��y}]K�Zb�1�-rt	C�T�����4�>)M*�L8�[�:=�K2iS��B������ ��\<6˕�!�ʦvŷ�cS�/�J���w�SmhJamQ��(V7��k�C�O��L���u��DS���.�Ea��n�*̭:3[0[?0��q,���[ Z��/�W�?�Ƅ ����hGx��Z�W��K���Y��4@���
@'����s�&�h#����������Xn�6��ZG�F�쬽�-�0v�D\[���Q�˒��u��>O:{'Kڌ��e6�>���.��K}
[�ǚf1D;�$�G�]vq�����C��˅<�[R��-�@��= �1S#� �����@ـfh�1���U%�T��1���G]�z�m�rvk��,P��L|��C�L���4���Wu]�k�TTF�������Y�htz)�Hu:pcT���yj
������y�h��oM �8�2�y�C�IW�#OV3�⭐M1m����I���X9JK��uReW:N6�gP;~̡�@E�ٍ���u^N�D3��O���RP�;ΰݾ89��w�ڤ4�Ǻ@���:,�,�������-/&�ɿ%7�-��[�
�\CȽ؃��jC��Z�Nq����@9�rZ)2�e�v9����ɰI��._�;�I������B�gF\�^1ۢ��A5��̝9Qd��c�{D�h&���Dޥ����cS�)w��g������*�B�n���0@C��2�Z��bS���HM��R�;Z0O;^#+���b
����D|�[�d��3z
�Y�1o�Щ�; ݿ9V�v臍�������\�����-ޥ�������w�ܗ��Ĕ5F�����u�g��DBςݡ|���Iw��)�e�5�v�i�,�ߔϽ�� �����gS��dx<�nL��J �Ļ=��2qk�����d��p1�c�-g��}�#|�&z<��?�J>@�B�Ϣ��heƽJ{�r�e�Fc��}�e�)�v_�Œ��d�Nͺ)}��v)XX�b����Z0����b��<c`�
3�Q{SR8�,��
[��xژ���\)p	��v� :`x����;���Un{F/�B�/�|q���j�n���n����O�Z|��}��)q�S�z\y)+�]��Gߵ���φ�7��H�����BS�
ʵ�0��S�jOB���|QV%r�j�T>;��:/��w���P-����9�s>��1T��C���!�Ye�]	uf660��>»��ߙ�R�UC�Bm)���Χ������P`4c�ga��fI�i���i����I��
��	���ss� �Iά��64&�S��i������L�6z�����ڥ��aJ|�;�q��dk��=-�߷d�S.�z��rA��t}�M,�@mH��I�μ�m�^W�Ν�����W"�g�	������7������Aw|e�̼�+�X%a��r��5f�/���KI�|�&���F���6_���-�i|�!�������9An�*��E�y�-sPn'��4Bc�Lr
��ɤ��cl�_@�$�xf��f��o��фTO�oqig��4XS�����׭�P`��р,��T��9o���%�G*�r�7U�[k���l�d�\���P�Dѩ���m��u�]�Ae��E�iڏ�edI4������׀F�&������[��9�ggDL�i���f�ԖFz�g��)8	�4*������4��܀�m���⎰?�It�G]���Jo~���I�啜U9��!�(!3�3Nqv	9�Ƞ̋Ѹ9S/D+�,}wl����|ù��Ge�tw?3�&��n{"����?]��r�_�Ӊ��* �D�v��$��q�fO�r1�eL����s=��+���a��WWΐCvY�k���.	��d�|�lr���t,onr�5�:�(��C,�wO���8̐z���c��V~�6fp�׻f�R+u�\ZS-��y�V���zb�C�eL��i�*����Ⱦ��'v'�!�cmcedF)C$hxN����f�����$u��U y��r+\�!DQ�J� ��s�e$�qt0Wޒ�bPT�I����[*�E.��$���$�S��#ж�6�j�>�~\K�%����$��l�wD�t��������6�\]��dPyu薧����?nџ�P2�W2%�����~
}�qc�g�xu�qxW"Q$�w�!b\x�+Q�E��M��!�� ���?[�T�>q3��q? `��L9���w�uJ�s�Qu#���������?Dᜒ+�j�@�ܭ������/��6�\��	)m�ӔY3��ʊ-c)���Z5�
b7�ro.Ձ"��K��䞲�*����
D�_Т(��� �F��x�xr	'���l��Hf�B�Z��@��I�mH������V`��I����$��AJ�d���t�߅vl/��0�o*��YoQ�i2;*fdjUL�"�P4����Z�<���1�G�o�pO�����4垰N�G8��ȵ�P��bǸ�}�3�Ue�rg���E|c�����#��O�S��cFn9^( ���F�yG1�,N).vD>N�Dr��+�f1���L����I�'/ֿ��XY�w�Y��]6�ɢ�M�V���3e=�#�<�k�-��%�Z�i�ڍ:�R�^<�
V��'�W�	 �l�S����]�����q�\����6��r�>�麵6L�*�Y,p-���y��7�b����ףd1�,f4_�%������F�|<�AZ9y�>�P�H���v�d�{���:!Z���d��|�16ƕK����j�Z���]B�4`�v@�
���ʊ��p�� ��m�+�V[(�Vj'$�qgB� ZsM���ui�����,<�C#먶�0������k�85X]�<��,�;�'�Mī2S�'+�p�!@ƿ��S��Cj |*[�9��sQ<:<r���K�q������Lؓ-��yZ#�)z��-��{j�q��~���U��(1`L���_ �aNbbŀ����~ˑ3���^	��h|4R�-�^P���G�.���q�{�<��	2;;Շ�F������I����Ѕ������˻h���b��LY�ȣ}�A��C,z�N�OJ�/N�-s��wO�J�zplo�򦃛
ı�zxo�_�.�N)i��*7�J*X���:��p�=] Ο��b9�]�=�8�)h�1�:O��,nN-���FQR�}��@�ZP�Kjՠ�?�!d�:�Tju��%�Xs������O_�ᡟv.��)�٪s�*�&3\}�(n��R\TX~sH
�1���K=�T�X8�H1���qޙ��l%���z �4�˦a�{��]���dfhH�B�!�����?l�=C9�����miŖd��1r�K_ODLZ?���7���-�v �Y�����M�x�%{,����'�"?�6K�t3Fʁ<Y�`�y	�	3��o��~~��kt��)4�(39��$/���彽͡e��@���+�Y�f��Ҿ!��kwԄ"�?d{0�9�W�p�{<������^�@����p�/�F�Fw�+!�\9��?ZP�?�%%��Z������k��
e�w�%�P��m���/�a��`�w@m��2t�=���x���#���v�oѸ��d�;}K  ��0����Ӽ�"Zvb=��{m�Ľ���+ ���)e���/�΂������$��_] �JQ�3����y�w�����P�<������D�e����M��NX�3X�\� 擻{@����~]��t�2	��4�m��w�n1��}�#i @�8��=��w�CWj�l�Csm%�.�w��%t����r�J�(n/'q�7X|�o���[hp,l�H���.�>	��
�W`��3�Y��M���j����`M�;1�^���2�ǹ�?��i��e�c3l���@��h�A��eF�~�Al��c��|3�w��������^A�>cZ�hWE���L�;�Ӣ��'.)<j�Es�b��|<Tl �)�3�Y�!���%u�N��r`@+��o6F�����9۟���I��2c]{QY;V���h3��}M	��c8��u�Ұn�gP�+�J5�T{d�����&��eh�[��eWZvZ�û����iINN_�QI(CIm�aw���G���a1�o���#�����`Gt�����sv����!�R� A&b���?�X����ZE,��F��]�Wk��ѫ?(�!���,�	�Ė�̾�'b���z1F�vg��C_;f/R����j�3wu������́�"o�ԛ�rӉ���+C�i�E�&z$�#�E��f�70��mpL�Su]���q��d����Ǳ�e.Ը��襛��ݩ$Z�_�wrϬ?K�����}\�ui����F��0���;�������ϜW��0�Q�i�ԉ!l���9�n��
;4�:���[�9��'n~w)�?<��D��KUcd=Iu�h��hVi	�	��^2��N���l+^����w?�s����[Ջ݂�߾��^��fO����%�o�܄~��8'zn#|z�4�c��U�Nw�&�g�BWR���Rm��ff�ٮ��u����?�����jc׶L,�i0�/i!E}S���.|�:h��/~�ĖH�}���+�ڇ��ߞ8h�1���{���ʔ)C��p�3E3���#L���ZE�� SLrL;L�YE� ȃߝ��*a��"�`�}�ճ8_��~tN��n)׵_Ml�x	"%5>c��Y@=+4;���[k4��������m�ĬM����t؊8�Q�T�1>���v*�`����o�0w�>.��4����.}�<>�7���N�O��P�l��na��{��x�,��h�oG�^E�iծ/��y�'l� )���-w�_��i�v�,�Q)/�wr/t�;�TW�7G��.m��m6��(B��F�d�~��ʎ-�]��ʕ��m?`Rxb�)E>��g���kmS��]+;ӎ��Ͼ栛Tze���S���S���Ϫ_�����Kh�4bG �O�,��	*I?8h�*���3�Ja�\}�W֡K�{'��|��lM�lr����O��G�V�D\���c*�?�B�O>�ُ���W��R܁�����<��$��t�Jޠ���t��ML���{�4�����ꊇ��c��E���1y��6�g{��,�*?p3B�y�m��I�`A�K�,��ɐ"l��z`��w
1�ΫP���5�+�$ ���x�1�m']�+��T"�5E��"�[������~�龂�t��0��M� KDuX#9nmp�g�"�5@����QS߱��
9 �)���� M��i����ę+,��O����`�H(�H�Q�ݒʯ�c�im0�5� q����~�D�Nl����G�'̭n;t�k�̸�1X�|q]a��eћ�C�C7-3�t)� _�ʗ 9�"=B�D����7���5�g{{jt+*g�:����G<�)�j��Ww�%�S��`Y�� $ϣ�S@w���L�h�J���9�Wr���Ď�e��%��z������^#��:�Rl'��@�� �W����τ���i��	�}�^�{���?5���*���w�$�*���Ӷ�"p��L��p˷
̇"M�`�<�?�dtjμ)���ݑ�(gݷR���P�DV*$�h�+�q������Tq���&t�'���/�"���x�/�� ϲPt��a�%b�s��;�/�ɔ�������TJ����,����.<�fߣ0 4:�FI���g�]�\
O���0�3rkIHa���\��$��a�<��M�	ɷV,j��a�.P˽G��Ӣ�ad�L 5��G<rYK��f�R>�~��>T�,�G5��y[��ð� ��m���ǻG���wv6)��10���O���P�X��dZ����d#ߧkA���>����y
���l�^����M��qH����Y�p���4��F!>�J�%x���h'�PWx'=�F���3վ ��t<�'��������a��Ϸ,#fm�.�^��_?�Q��F�-��d���������wB+=�GJP˛h�(���Xdӑ����n���Ƃ(��(W�k�a��c�����$�����0N+7M(���o�4�2"/�������r�̧�82��������S�u� ��w^t�X@:��w��g�ے5U WBe�	x"Hv�u����ڡ��"J�z��1'�:���Od�
�C���Ñz��: �o���6��c?�J"j.e\� �����2Ϥ�z�)ڱI���VJ� �(d���^���/��a���Ś��A�#��"�� :#*Ou>����F��x/��F̋N� |�3]�@!`.0B�9�"l���CV$��(՚�����30�V����3KN},�4n�#��vsCa�C<��me��g,���ԕ�>�vg�g|a���U����]�19�#j��ҧ��%��/����.W�Z���R������J��6Iܻ?P�悾��.ؤڼ�#�w(���}����'���bj [9~M�Q�iY��`��ﱻZ�\	~o�R������D-�Y������tԋ><�bW4�W9͑��:�x-��Y�L�zz�;�Tgw��%�w;�GTs�Hq%�ӻ^��	iZx3�A�5��~���� ���ʢ�6ul��ۻzk,�gJ�(�ÑL��\h�	4M�\�C�Bsi���+ �>s���y�E�fxٿ�~����< �����0���d�.�Teml �_SfA�݉��Od�hb��?sh��47
8a��b;���ُ�Z��<�G�Ip::�2+�(���nݥ!���'n砒z�����y�]��du���;��j#G�[�%`(u�4YP��*�6El"��4����	���e���n��@�(�0q)#�D���̿�E���4��Fγ�V���020x	���c�U-g�H,��~>-��e,��岵�H������O0�~�Fr�eZ*1����̏��(˳�>�,�e�i�h���s����/L���H�@�;����)�jk;,$��}�X��2�Pn�1�˭�,��oM/�Y�g�Y٧I�X�y�G�hq`.�I��<�_,���tP��� T�d;{�r����	�O��[�&�����V�q�]�������f��E|�r��}n�W�i��geF�4�(����}�M%���>|04�biUJ��|�t��`�}�9}B���L4L1!^���)�tNy 8Fw���Z19���͜ ��4�{_TKL�Q���W<��l�C;����R���U�F���T����`�
?7$��2�_`��o&��i8PщSƊ�M��o\��J��V�����]G��+�����Ewb�k��� 3P�' J�z0(���g��8�w/#�m�K���d:�0�,g�o8s�1�����M���=��J�t���(�6{��QbK�XYS���d�75���ug���DH�~ҍ�k�?9d|�_?����u�iM��%#�ˊ�j���!Pd����-����$w6c<0��X�@���B�����-2��&�i����B��� �Y��w�!!�h���Q�E�#;꠾"���P��1'y���02%�.��!����(
�h����C��џ�kp9
&�h�e�{3|�u	X#�C4���
I5����|�f���QgWE��9��)zfR� �A�:׉�#�Xմ�e����%L�R�-���� rۨ�>��y��P&��Oae |�L����W�u߆�1J�p�cΠ�m����V��n�٫��p��~��R�O�>��V�3St-�(�������ꏹE���Dr��B�3��������ґ�\��z���N��D[�5jn��I\�uy�AZ��Ys��7매5���;�`�-�xS*����uGm�I�AJo��d�$���<��d��#جOv_'2��9?Ӗ�H�.���xA�w"1�5 �Mt�$=:�ʆN�*���8���o.�7��y��zv������������l�\uOD�q:z�8<�嬼�k%x�9'0�'������@��&��N�du4��	ɜ0��[ �Ӓ�淤J �q��t8i��ULSl��?{�4�
g=5�֝k���I�@06n��=�D����E�#Q}��;���=��6��l�D�	8��� Q���z�1�k�e���1���7�A�P7³@QoI�녢:��C]VSP��6d���,Gb����=�M��Q~����/NQ2fU�(u�מ���@Ӿ��~4]�5� ��rv�M-����� �}�f�`�1H�
�j��v㑒`'�P;B���~m�W�b�A����B�äx��Ŵ�\��t��8������bYn˂�:JM�Y�֮���)�cj;J?�����D*u&�O�9�G����*���� ���R�Z�ޕB�sM��'��H�%F"�]��N���R���m�z��Dg��x�����*k�U��7G�q`�L:�Վ��',�h	�G��&=;������S�,6��蛠�S[�$�6��f�dW��)C�*�)��g�k�Ƌ��GJ:Ct��ڙ���~p�{.�^�> �s��j���Y>h&9E�?��������`���,�
֯ڴ㊼!u+k�2�6aj%�T�`�zOO�\����?�������3�%)�_��mO�]OvK�3�6�ƃgǥ�kø4ϱ���>�T#nz��>߫�k~��r`�t-ޡ�g�W�8�~�=��rHH>���L��O%鴦n��Ԣ��r0�dmz�Iό~t��ީ�$�Ϟ�5H�T<2���re1��������ϳ�Y �q��b�Z�5�B�]�/�4LЖt�+�%�������Trb0���=��^m,K��3نƆi�,��_~�	�K<�>�b\>�0�3�41��OF��u�Nyg�6����T�}��t�)��w��R�6���c=��>4���"F#�4�U�i�
�d@��.2~�N���KQ�?�ЯB��$��KƁ!��-�����j���'��e��K�W1�"�Wa�K-�k�!�R��*āw��;M�u�i*���]��4?|ߦh���x�a!���xx.��p��7�t1�RL!�ߪ~gW�B�]oS���0�
����G�u�8�ym#@�Q���,wQ����!-'%M�ֆ���ݛ�ta�5���F�H��ȅ�����Ǘ3��ʗ�~)O"E�,)rRa�K��'9������@{˖����W�IT�O���5��<f���W,�6�M�2K�|�7\Wf'���齻�Mf;�3'%�6N�rZ;t�t��W3�J�-y�1�կ�e�.����?�8����+������qm{�VhTύ�Y_> �5l�8�R�F;(e�3�4����Ƽ�v�ߣ�e�"0P��؞��r�
�M�-�� ���#�f�샴/�&Zf�-^�$d�҆�-��'69�|%a(!����L�s10E}�*�;>�����j���� %�q�к"��#WL�ؤ�ǯn���!Ȥ��jW���J�������J�N����Н�ճB�[./�F��̯������ЋZa��|ֶw�R6=M"IT�Ũ�z���c@!�|۽]�;t�n�U������6`Ǫ�㬤���O��(?_Y;��uo9�SҸ!� |��8�?���o�i�!�&+|�x?S�PZ�͍`�ؒ�No�8��P.g �(�2�m���0D,�U��I�CϪ�e/L�2
��l�E3e"v�\�<L>?�rA��?��~;�W�;�A�;#=�.����t�<{|���K((��Dð|S�;ޗ{�=�%�'���w�D�N��%�$�&�]'q��l��@����o�$}��$�|簕���U��@M��������O��[L���P-L��Rn"���v^���Ʃh;3�׾<?���׈F<E*:8�؟D�=rS�~�6���Ap��+Q�Y�\�ܶ���#�;�+�/��db#�Ng�֍�AcoX��M$MJ+�C��|�wW�!�1��p$�r̺u!G�*��ݸ�l�̣Xt;ȍlZZY�P�����u'oз7��z�5˂q��F#fYz�L5��t9s\��zE��-�G�I�@���t�]� ��� ���tu��g�H���4G��ނ�����1�$ǻp�IO�׌�k�w��3�4|�-nY(����%0���b�|�s�{	b�k��7�l�n�kkNͮ5�U�8Kt_g:xMy�p��;Tj��f�.�~|�էt>~�Hܶ{��IN9�;�'�7�@aB��\8��Z�L�5�n:��p�?�x˾�2��k�͹�������)26;�G Kc�C��+*����4��$ӵ�m���%�*��V��/�L��ɍ?���,��/�m��n�/ʵm�3"�Oq�?$m�m7=�KO�#��؇�����GvQ�wӑǝi��*�8~��_�åǎ����Ψ	,�Tm�z��%I�6E���}1������֭*�N�O��R�Y�Y[T\T^^�H��D�JA+Q����[4<xqU�c=�T=������}�9$�(YE�q:5{��I�+���n}��	*��5�!:��` �!f{j�ډ>�9��+���S��]])p����������tƙR���,���j��8,P�f�pk��|W�2 eyO�4����6N�T��V���;w�륊�LɎ�y@)�y�!1�%�e�H������zu9+�M��
�ԋ��/����;� ��
T�m�{��s)u�پ��\;�D)Ͼ��N���B��^N�$�����.�Z�hI�ބ�9Q:7��ȝ<�~کT( �FSB_�aB(3�H�a��[(Sn{�P\5XZ����� *]pYw�0]�G>�ƞG�^�c����Q�aZ	
,7��J���\���Zg9Ņb@�U��	:X����XE���
��h&�-{nX�9��8��K��CAJJ���5Y���A^z�mx}ga���SN- �홐`�1Y���2j�9&��Z^�����Fjq4
6{��/>�ފ[�«OQw4ܣ��W�z�v����9+'������%B�+�릭�ՙ��Z"���Ӌ�=	��rC�}�t
�����Q�ay'^v��N_���3�%g�q���b��E5���MgC�b�eRs��A-��}3��$���O` ��UE��x��}K����	o�k	�3���q,��i�*��p�����?<��;z߲*��\P�G���4�>��4]�$u���hg����<P�n�aSF��V|�dZ�����������w�Y��QP�/�D!;Dd:f�0��&�a.P�b +��v��B�7�	bc����%C�*ʻ/�N��·��Tc�(H"�?�h��6�����z��˹��� �>��%����q�����0 ��.�}	SD��R������p����o�W�wL
�t�-bˊ�������`vX��^�-�
����΀��㪓��\�"7����.����[�u�s՚6�95˪���?l�����2=eYU�#�3��`E��h� ��pf	r�ä�}`F��g���
>� I�<N��*/�5�Eg'��0�'�8���k�Ѻ\6�~ෂ�!���j�a��9 d�Y�|㶽���}���#(]���/'ʶ������U8�~��AsW�D����
_u{�u�\>g�'��iOd��i̪A<H�,��H$��Nܐ��ͦϷ4��N-�R��5�����d�(#�����R�`;�j�[\��{�J�'w���Ta�=-��Gcj-*2 G��3e��tp�L��U�h �
�FPp�.�:W��͐۶-X�kᬔ�m髎��zT�=��RB�H�L�n�|�asl�ؓ�*B�N͔$�ef�cD�s|G���BK�C�p�9�O���&;7����I�8n�
?�=r�v�^O��WR���Oz8��^c\<�'
j �*eꈵ)�:�}������Q+-Y�K.� Å�)��)�լ��Jb:�~G*��q9-��ZR��Q�υr�_&��(-��f1y���v=	SPԲ{&�裢QM�tr q�zs�_�] {Uc��*�|��An�c֭=(��RI*]-@��`��q�ݬ�>�W���&�v�S�r
e�%��} s���|q.��h;�sGpw����~v]f�a�|��5VF���1�)h���\�����i ��s�����#�\��驞�3�8*k�R�-qX�B���4X�����T�Q�O��B36���	�%�tor���tQ�sè,���4^��%�&����gOK��k�dn( �A�X�/�ܟH�k��wf%8�8��b4Wz.:V
�]��~F�b�~����xS����&g"�Vi�����Cg�τ�7{Qu��_r�n��^*t	�,�v��s7컲p��f1u	d|��;�!�]�8M(1%q���`j���x�-a]x�#?	��`n:�~�'to*�d���)��.�}����tA)�8�Bq��2�s�p8�ٌ1ߴK�D�iV���SW��z�1����Ԫ���8#<��i�gѧL`�;g�q��f�����M �!��$h��0�Ҿ�W)�g)'g�/� ��&.0��!v�v��R����� �R��	��%�����%�5����N��r�]�|�אzb\�؛�m̨�NL����\|B�ȑ�\��/�˺�3�jvꭎ~� ��o����=b���C���Tn�=n�$>Qj����ĩ��8!ҍ7�4D~8�CJX%S��\T��쒺��K6���|�08�Ǻ�]�·)�+����^��T8,�?���`�ØK'B���Y�yІ)8m�D�Z)_�����_4��X����\2矒 ϓ��+��k������J���A���[6���4��z��<I.Gv��0i��<c$Ll�N�-z�Ρ�޿�#<*Ǐ��5�W�x~;�����B3iN'�H�fg��V��1%"K�:h��`5��,K�Hk8^�c���`�2F�9��x,�'��K��$�V[�@3��}�4��!\���ejG/����51���85���-� ��_�����`�+��>��"��4yP���\6zt��O9O�(p֡l�P�n՝z@m���`����Uk�6���h���B3��1����+�aJT����t���@�S����rL��6�lmS��g��$��Dy!+�-]�]��<����lS �T�&�"9� �b}g�(Z'�E@�ce�O���1����N�{�{�Y�vƁ�U�P_q�t���+ӑa�;cp�xO���������#�c���}�˄���NGF]˼�1�*k������ )Y���J�����b��� �>4��F�a^�g�i�dɨ/�f�����P?���e��[@�`�����:��o���:��.+f��,H��,�g案w>�� �����B��͖������9�TB]�Eɶ�?��k���0��:���+�*y��S�	��8���-�.~�h���)e�i�Uǳ���uǁ�Ֆ��@BOx�F�$so����4�S%���Ay؉282��E���V~S�J��t�ftĠa��{ѹh�E�g7P��SP}Q���k�3T���|�U\�U��,MI A���ceY�c�Gd#9��u�S��0n��-Ce`<���Jo��z�yc�N�Ggjٌ6[�Z�Ϟǅ��l��<��O*n����q���Z�g��jٺ�P�����6
,�"PA�N����Ahᐏ�ڑ��3�V݋��PI�t4𿪠�{�hiֹ�Xݑ�ւ��`�gar�]�d��ꇐ=V@�0��I���v?��J��\�l���5�nwZ�Wó
I��W/�d$��e���5�:�)�m����n��,G�+�0iJ	`P�Ĺ��E��đ��I���ò��t��ހ�*��	������4�y��l���N�;\�c�.7�ol^GI�DtXho�������l��?�*��a.��R?+�i��q��VDϞ����58���
��j���@��xa�c#���R���$:׌���*��A-�A[��Ym�A�_�6�.
&N�s"[�4����c�����%-I�{x�������ܳ�0���N{{XbpF��"���7��$�t��3e��@�m:ZK=w�u�E2��J�f�z_<IB^	dC_�?�.����Y�\�v?����d��3�=�#D&�Ҭ�Y/( O�s�k��$�a��[폏$?��9�����Yȝ���!����}*:`S�誙X��r�X����;�`�-���D��������g��*PXz��b�D6�vb������"ை�\l.^�A�﮺�Y���1��4��)��ӸȺf.�[��E�i�c��/I�9/�	>�,5�b}P�.��Eg_1kkeaU��p߫7=69U�d�b���t�(̏d|��T����δ93G��YB�T�[����t�Yza�I�%|����_��D���S��v�ّ�>�|��ޜ�%R�HeE��.�簻�e��&R!:���*��j� Ba����
��!�!EK��l'bvl��S��������`���4�q��2n�Q����Q7dp�?��j�T�/E��+�`�犷�����t�0J�]��X"zD��M��1L9�E8tP���"ҲB+l�O����Lc�Y�k���0��|�h��5�Tz���et��:_��0x���n���A��)ՉI�^�S24.�[�"���E��e�:���.���I���G�	o	�S�ů$�=m��*O����WQ��~/���iL7�8�Bp>���y1%��I��RC�K�fq����J�������u<wۥo����j3ƅ������Ve�h��I9J��p�U�k�w�L7���p�$��j�EȻj8���?,9����`e����7��9���<�]�6��ݶ�!0�8g+
�YSF�Ix[q�t�����e�	�T�O=S�i��� �=���x�HG�v�yTDcGA��Q�Ώ7)���,p$mw�Yf�	(9��x^wߊ�9U�"1GF�H��Uu�#�ċ�g��ΘL�L������=b��{�����/!'��dk��6#O��ᗒeS�����q���6-;c�`R�L����d�b��(F�@��E8x���yG�Ye��떂�%�OpC�y�=r����Q�`���%��g��	<D�eLDh��'o,d�8	�fx�٧�M��V�na�R�J���� _��[�(h�r	++V_�[w�3��ZhN��݁�9�/����в���y�����K��1�H���apP�pw�N���Q���!�,�k4��c@}P�Y��7T�S�8P�}��@"VD�����U������Bf6�
}���~ċ$u�ȴ�O�tް���Ҁ�s�Y�!�)+��e�,��e�7`���o}�DFǭ�0�!۾2:)@�8����E���+�Y��d2������!��c��b�,�<�2��&����1��(Wfw�![`�BZPm�Q�#�:9{��]���V,�xb�?W��C�d��/�7e��E#�h3�2d!����a&����M�z���;`
M����`�+�`ˑ���I�%=�΢��sF���O��p�R\D���!�/��/�l#h'�A�0��t3���V$й�B����a 2��%��I"��p���o<-p[8h�\�X[���4b�>y���S�q+�-.v,wi�-����e��^��c$��9h��l�B�H}�}���j�zvg�6{*6Xl;���/�@��/z���N��j\PE��	F��|��W�k��W�Bb�O4ؽ�;쭌qV`�o��[��*����V�-��,�j����r+��D=�4�e]�/T�l�wi‐RMМT�����KN�E
�����8���c+��$ن��=�Q�l����fAß�!�y=�gr�x'��a��\˚�aQϕ�8M��F@.�"�2".:� ��� h&�S���`4�_�$�h�ⷨ��T����w����b��|ID�n�U3��?!�$f5ph��4.?Nꓕȴ�@A�yah|�#��N)��ӿny*U6/�P4�h^Y���B�`�w��?�h,AYi`zh1h��CR.�	��DBw<� 6��R���O�ģr��|��hf^�ң�Ϝ�K2�j2���
���(p�G3�㍈,���*-cӋ3Q*��[��j�묲L@�fκs!����f7�	��1�2�0����:6���G1qkF�f���.GJ���8�~Pa�c����.v-·.TTG��CIDӖ��]鄆tǓz5φ8�r�����l��',Hf=4	�{a�T�Vz��iI=w�֌�b��mw���*:�,)(O����r���Ň�?��qn�������@6����!T����;�A��J�^0�dSB�{��T-��y�Ю���!.�D񸼔Ӄ�'F��&�?�ͥQ��	Y�xU� �
��ћ"���A��rV��jk�%��p�����)��kh	`1VL�)\%.{�"��ݹ�N �>߼��FM��D.=�Jʻ�f�;d��Q���/%ưU�� ����.ݑߪ�"�:8٭�1B�!�ࢺ�I�g��\?WJ�����V-���8:r��37͑�k2�������\,��>CF��ЉZ@4���aE�#�6���N�4M	*��@G�kF��x=��]�Qɨi��>���@��oB��R�Dxs�Urʉ`���5�#.�HJ� ���/�8Ȼ������B�t���t�����7+R�5�Y[Ŝ%&V�5�"�0.3�}���
r���g\�R�� �_��oU�s2G"���%�m�6��G���ku�q<��*�>׃�:e����~@�o����C��=��z�(S�)ܻo� �(#�������BBg�Ɔ�ċ^ã���������[x�����B��� %F�@gBA���"��
y��=�᱈{��߿I�����-���Q�hKW�θ���t�wy��#��DX:�D:���K{�c�'���a���9�G���r�x�2A��mu�w����!�)/u�ca�덳�{H�R��n-���t���G%C+����c.��<�Դ42���n$����&�
k`'DO�/��V�|���y�&<L���ê�\��>T��e<���eg��h�ݕ=�`�Ps(��rD9��3|���T2��m���S���$��us$ki����Qb�ytM����w83}˾�;j�N���2�֢�?��՗~�Nq��k�7�y-�O'ɬZOb)�i���f߈��V�xb�똚Y�0��>�-.C�fO�r^\�"?6����V�W��:U����D���Ї)d���0&�TUU�ON�;<!m�K��:���~�7<��	Ji��Ou�H��p�qbݜG5$�1��]A@ĵt�4{G.O�}�A�:�C�#c�o�MQo)3����y�r��>B�<�%ڒZJq���l3X#� I�Vմp6~G��h�@4Ėd&�ڬ�JX�2�>\ W���������NAю��)���b�����)����Iw�ғ"��s�OC�Ew̨	�@�F�O,l{���s�:&ŧ�2V�(�v�a�:ڿd(
��蜋�� E&Zyt��B�C yL������-e�L~R+����w���Qȥ׍����+
�dP8 �4hG%��ʱ����iv��	ih��C��U9<�(���"�Țџ�*����u�Ku�v<W8c��>����/i;���c���s�OAQ�% �nAC���W��,xCzmibV�\�A�ֱ�tA�h��E�N�,Uwz.
�ŧ]�"���\���0L�&/{QM?S��p&�1���z_�h��)�!n���3�3�~��Lƛ4澕�o��`CĠ�F�g���cC�T_6�k����
Hp��:�`c�Ű>��֪d�l��i4� H?�z�3�`@�������Vp��5�C#C镝v���{䮀�u����e//Hyx��c��ONs���,6)gV	������zX�$�l��X;Q��Ή6��I�"�	�OT��S��y�qK�R�ۓ��>�د>5�jό�!^%s�@�ّG�G鹏�I�X	Z���+��Cfw���oc aB��C%� �J�t�9+\(+�Ӹ�c���>�M��F�Xrr#��%)|r��h��´����:�_�Ե�
�}L�Y��1����>�2��@eD?�5E�9�4���$O���/�x5&��F��蔭:'&~Y�k21��C�;~�����̛>I��ld�h�Q��nQ�Vs��࿨�מX�Y��`���q�J +y ر�����n�w��dh)e=.��������6���e�_q��i9�o�	g��'���q�>�7�ޗ������,�}��
�s͎۫�2$L��i�S�"�I�����q����:sV(.Ԁ䵾��U�f1a]�u<�=�a�54
��w`���W��1�C������wI�G�U�C�:L�}����: ��H�9EG�.������Ђ��z���z���ON��P!�?�U�����GcN�a����Oc�c宕����	ך��9�U��^�K�ȝ�ʤ�1��@��PT��#H.Ą��\DZ�`~�_b��"��[��M��N��aw�8�gr�.#@���]�����.tp�Nu����t�呝�D��O�X��w��0K�%��n�Aр�|&���A4��&y�鋉F����Ŧ�[��l�E�,�̾�w�e�z8�q`�\҄d	�f�����d�@��=pVϯ@&��¬Qb=�!FFus��HI�וj&�I��E~�A%/�]O�e�����!�F�;�8QChq�](z�M�H�)��^b:B`IY�W�J.[�	�h���A��v��X��lB-*1�9u����/�F�ˏ���(ZE��J��������o�9�=�!��t���5T�f�����Ϫ��_����\v�,��}[6�$�_㩱��>���g�X<,��|bi/���,N��®�ɡuy�- 0ځ�WR��.��H�+	R+g�VS�<:�+'��7n)���@3m"چ��&�b�A��kz&�5���;�}�5�h��R�e	�uyNص)��3�1�C�~���u�J�֯�v4N�D��)Co0�f����C��j�XCUq�_�s��e,�=41��(C�Q#� ԙ/܃ ����	���� 'Í�ﳬY)J�}�
�x��Y�j��bwX�U�UAy�t� ��@e������y�=A�	|��_WP�e��=�]U�	"5Y����UZ$ys�{.���H���o�E����[��Pᇒ��>��G�+C�j��8�N�6�BD;Fk?��bmy����,�x/��7 ��]"�7�~b�d�"n����6],6M��.C�΁*`�$Y���n_��0~O�0(L-��4Z�y�� �3",ut�Kv�tAY���~o� 'A�vU�n �\��p#nׯ]���S�*�ŒQ~c���~*�O����瑆��^%�c���:{H�}��V����Y����m��m��I�����[8	�����1$$1b	���,� �Þ���I�:"�O>�($&�t�.�CzZ1�=e#�P�k��l�%3���ZL�����7Dg���$u3Oa�
9��*��2֖,�+�f��_yF�_�lQ肙`Yʃ��9�-f6���+��ц��g�Y��`�p��jf�C������P`H̋H��b�↨�ͽ��w2XF�P�"���Ia�I���+t�A�s���*j������2�%>��y󪰗j�	]r��0�#E30dH�����]q���[��M��W��T����r�W#��ݓm��@��{~$.<���bU�0�X�d��d
��P_����opLU[���t�Mс��')�n*�Gk�N�m��$ǃ�8�M���[5�����e���O��l-=���a�b���
��%R�9�/8[o�Kb9]JXƱ�X�ْ	�#�J�t?Ѝ�t���
�|Y��u�[O
D@L�;|L��pX������J߹)-��+�#��%C]�T��b2ԀS��R��d"�&�E����vyxAX�T/W@n���\��[�nn\Y@�P�����Eok�0H�|{Z������<R����:�"�>��
�^��Eߗ�;c*����0/D���r,ItI������Ӓ)��Z�����:@�)j�Q���$.Sy8!@Pq+=��;;�gi&Gk'��\h�~��#=k�oL�g�A�H&V5CױT�WA�%,̿�0I6��q�:��/�5�pY�T����<j��ycJf~�x�ro�g%ջ�N�`�6Y]<0P���ŐU����&�]h{�֏*)PL�ATԢ�h� *J��B�N���I��vƆ.�w����L��E�=�f����9�o����d'\+N�5Wm`Ax�+����s&�tch��P+*:#0h[�X�3����ԝ��ȸu6�ED;��Pn"�h<��Y(Е��ǆ�W�0�F�2�Ͱ'�]�j7�L���1̩���i����p3�=p�����jD����䪳�P�tK��(�@���_.�:/���H��=L.���[�����zO����>
j
�6��;&��I3�g�$5W�p�^�bس�n>�)��la��*�)�먥����`�
;�����1��6?ή�����U �i��ș��%�2*2	k�,��Z���#j�U��ߞ�?��sQ��7 r�kC~���̓U��W�=��h��4N�5l��t�DX5���(4�2�����KH#���!B�bE��#W<dFAmǚ�.w�4wZQY��E@0��>b�d;�$�/O�{Ź2��݃����T�p��aV,ƌHEO�y(�c��l�+��b�p��1��g����Ѹi�";{Q�F��9��{�q/�������?"o�2g<�w�8઩���ݵ��XS���g��3�G�*/t��/K��^_��	�����y>�ɺC�3�]�E� sޢv�`u��r(ͪ�<�C�@�Ϋ�~�v�.M+�c��r�~�}pѤ�q�v�]��Y���S�s�R<�;1��{8 �У��t'pA#=x*�yIX(5�_y�"�V�qy�p��8�ʐt rk���`W���dwn�5i�I8�4����WvL�0�"y"6��K���:-d�ے3�]�&��l�ֱ�l�6��Y�O��,\����#�]_@|�F/"�׈A���.8��pax������ߴ�P#�2��]����b��tD��|�52��B�n�/��w�Y4zF� #d�p��g�ֳ�O�J����ZU���Q��H4��iK�
�ρ�q�e�?���G4kIh������t3BSA$�t�)wXz�̘�@���ܠ��v�^�p�E?�G6���kɺ�?��η�B�H�@3[�4=_H*�8��[Mf��Se�T����*[.Y%����ei��<�2���Û[���ɀ����DË��؄pz���hȷ����!�>�kq�����y4o���J�6�``�!�����To���U5^7ɩ��?A.bҏ#\cɱ x��'Q?V��N������XҠ��\1�b-����c�>E��o�*5�����QhF5P@��X���C�[��"gY�cH]�-�-���bG�֛��hJ8��е��'�
�fM]%#�X�)8`��
����N���.�v͎�\!6=��][���n<݋�`�����dA��೚T
F1��q"���{���H��.O�P��]���p���U�I��$��J*��M��h;$����:8
������I��~0ᩝA�2������-	�0�O�P��VJ��x�%2*]=܍�]i^th�2��ϗ���"�n�c�N4i�]V�0JM�nd|]Ό$@���eF�^=��L.?�Y}&k[]��c�/����0G���BY��,�c�6܃~�!�f/��W��I*?)U������&b��u�i���)L�V�Rl㉡� ���ဓ�.�ԏ���d	
�X�>�]�\��v�����1������×���62#i�<R�_l��v�n���T�(��jX�H�X!<�
�t-���J���+��b�c'��=P<��(�L
��^b�����K���8>`��t�D��z4��؆���Kiy��C ��w��W�	н�_��oR�Z��t�iC�3'��G{���C��IzY��{Q
?���[�[{&��L��i�)=u�:mx�&�ռ�v���C�I��"H���K��i��wAv�
���z�A&C�%u��fT,�K�}3��䔢`�7M"EyS��'��B?�)�T���!K%ɏ�)�o��>3?R�,�o0�������n�_-qq��e+���yH9$~�Xs��)��X� T>l_k���{�S�-G��磐�����C����e��	Ĳ#ϓ��m^�2p�GO�A�Va�":��q���R�"��i8���L+�?^�"������W��qa���� i'��/Lƶ-�$ezѲ��;��*��f֕Lmza�
r�4�=y����6+��,�W����7����'V�ۺ���+�XY,��&TN2�
]@0�����{�U�'�j�8�����"(}������oL�����v���ҕV�	��a�X&3wB�{*8w�ֽ�a6�BPVC�ɥ��C"�l#����}��r9�t���R�d�]}w���(2���Ѯ�����:�n��z�H���5�f5Us����˗X��2�U�w�U��	���`
�5;5�O|�ߛ,> \�}��G��3[�](���?��܌T������5��|����� 2�x�R]:Tn����M����xa[�^I���j�_�x`L���]�ղ�g�J�h�9�l��Rxg��������Kh"Cf��0�:��sW{�(�HQPJbZG�?����cgF֟�t��fȓ�eᇹ!�n����F%��9�g0��*f6H}���v������>$�^D���$;L�|~�D�*�f��t�K���+~c,~ �C�������j��ή�TF�m̌�:L����\/<���$9���8:�RL�o������j
�������y�>|�*��f�΃b�eQݬԚ�w+. *70���Tw�_�rѧ)�^�FR9@�쀨Čl�M@z��8�EG�;I2G�(�E8�}��!�Ҕ�yP1�|l��?1��I�A;Qru�5��,�%!W���xp]�B�8�(�e����2�)��/oo����k}&D�w���?x�� !~����aUb��z���k_2Oڧ�iA�BJF{"��2ۿ�%�{�Qڒ��q&�LBFg�s$�Z����{���@O�*�1Ĭ�f��:I���;ٚ:�*	�𡄄 ��CI�P���5�9߄�XE�M�T��_�3`��<h����K0֥�>S� ���F�G��g���q�T'~`���uCp���st0b���/N;%�kv,I�����ʎS�F�񣤄�Q���n�?���h��'�	-;5�ÿ
!��e
�)ܖs���_VB�Y���">�u�C�B���o�8p���:&iM;=&�lmNb~cih����0B��C��i����.Ac�M����>���O���ƃ�mꕯ����*)��^�!��i^��9�I�f8re�KMn>8:����#�A���J@=� �%`%�0���WB���1�ͽ�V�^�ν.�W�Aޭ�O,x��N�$��������Rh�H�y���}y��ǣg����LGn�̐Z%i��Ʋku��F7�	t�^�u�b��`@%��bBz8�W[t���x��c_�r��s1 �s�h��^MǙr�����`��SC��Ǩ	�N��!��P�YZE1d����a|�=�$�V�qk��#�o� j���=I���K�gv��_)�M"��c��A���ɕHu���1-�۶OϾ��v�t��c��g_�8��YW���}����9c���S��!x/|i��4��� ���~%�&��2v`tc`�ن�0�*���xq�'6!�3�g|���<�����HUc�m����}�? y���
�����M "��=�jD:by�AG&�1���6��Q�56 ��v�O�c��C{�r�ؓy���[@p�N��L��g�-�6EO��i��(���A������g�F��S(o{����(Nm�v������d��V�k���y���Nu�5|LO���������@\D�
:ܧ�^p���Vi�O�*�p4��|�� �um=�x���a���'A=��h�b��V�DO�""��ߛ����ہlF���vj?Ω�ʨɾ� 賎�u8g�uf���������������J}�D-�"�M?�#J��GQ���º�b'-�U�2�
Q`��jR����5D���fʼ����v�4�>�����1�����[�'Um<���c�uާ���À4��c��}s��T�}�J��u$a�[�]EK��]TJK�FӰh�B�>���b��o��4H$ت���&�%;��A}�
�:�u�y��N��ggL{���	�oj�ϔ�׺"9@y9����/��{�KF�az��>�1��@`�uTm`�0ǿ�3-����U�A�مG}�m	��F�9Q��j@���.7��힋����E�._�~)$�tR��2��&�n�B����������D��\���7_���8J]�������_E!�lX-/�9`!cRx�;�\W�����#@~��Lӑ  BqD�ge]a��wv�h�\f�G�S��G�A�[ �G����m���%a�^3Z@CS�;ǝ'�Le��M����"R��їJ����sԤP�`/]���/��f]C��tL��K)1K,܉��u(�8sXm3����a�둑���!�r�
��K�ܦ�+ʀ���X�oR����!���^$��2�]% ��5�j����)�D~�%�m��&��
�ۥ "�{I��S7��;x�!�vf�R��+6�_X�!�<O�>�uQ�ۖ[��`��B�|�MgBx�w���*>�i�G�f�C[^�*	��
����|����NYd��j4;��ԽF�C�yM�~Q\�c|f����0�,�҈�\h��],7�[�h�\�u�v��6�S.�A�r�[�:e퉙E�~��1�g/����v��*���7�~��h�e�'뻽23{Lo��i�!Z����	�"�Y�������Ot�B�u?(�<B����m�TOuA��+L"�!֚�"XO�q}�H��4?�<�&�|_o&}��A�Z��zfm�8{()�ى X��L��r�l��}i�"��x���`}����N�w6*�){�� =y)��?�xY���4�����0�h�xGU�؄F�	�7���j�4�C�a���:G�,>ޗ%�\�\�B.6�K>�Z��:w��U���*W�4ܡF���z�οB�PUOC��kf�$$�1]&K��S\���Y���?2��e^����d����@��y,��5����lsp�ҙ�v�39�Up��@�������FKK\�z�ȡ��a-eD"G��)��7A�O��ZUc��̞��
�q�d�Ƨ�}<�=US��L��f���y��jCؾ���F^�'���Im�Ʃ�p��H�4yyS�ʚ�E|
��R��[h���t��C�<l��G�����,�{vF�>b7�9�m\5JIѕ������C��|��h��ڕ�����^��:|������Y�}�I�G<��/3��W9͛�(?��qu��Չ����:,��(=��q��P�����?=�M��EE�[�c�pD~Uq�{UO2�bB�$��*(�i��#�q���(wh��N�r��&邿�VM�����y�!.�"%�_߸���>�M�����{�_B�#Z�R$ /��W��9l���Sـ�* ?)�⯁������3Nq�� �Q�g�%DtM�M2��+9�MY �������eU�;���{��dyַ�<�B+~� ��T����/�g7�]ҹ���e�0Y��?���\EH���T�����tǚ�I/�!r�"i�����S�"6G�W�����8����_��o"�H�2���}dI�Hvjq�F��⠯/���|�f��0�n�ی.0R��g��}k�Zm@�M �x��YL�X��|~��)�&�Q��/�3��E�օ
��0n  �6�:t�y����E�>�;d�_*��T��A��P�����;xD��}9l��4�=5qg� ��;з���, ɂ	֚g����F�ACf�@`���D^e��mv��	�ؕ����X�ߤg`��~/�Z��ˠ-x̩��J �tC��b�tʉ�՞9r�3��3�E�*�K���L�-
����2Rڏϔp��݆��A�O^�Ag��-����8]=����A�D���r.���}C�S{g��4�eᱻ����?E�ڞ �;�և��S�d�^�m悌�{o�=NR��hQ���`�LtW��n��qXP�v��cO�}�8�����7���[/�r'�	�'U���
T��S���m�hM���������*)=����j��=�5NPB�U[@SF,��*�	](��f���B�(���p,�T��h{ ��6�_3���%C�J�%Ț{}+y����T7|��"L�@��f��j�/��`ܤ�$S��r7(�H�n��htP���
ɐrEw�}
o��v7�LaC Kcޥ�2���wOe�do��p�W���bý�ƕ@]���c��+U�6��'DrO��cn_,{�����>殾�!Z���cb�t��������PI�!����tB$~#NK�Z��u�C`�G^����Z�n1�������/d�%wX�6-����N82�"���y��:��OL읥�xĊ�{Xi�� ���k�c�T?U����O��^28��t]�x��eNjg��Τb��(Mx{�'��%te2�R�?��|D(�"�S0�a�cQ���IL��byZ�8�fJ�X;���Kp4 /b:s�ǒD�2c�͕�Q&�9�t�X�������Rz���Ja���t·��5E�$��A"-�_�i?�o8$��O�U)_�d�U��/�%���U�c�D����p��XЊ���S�e�O�~ٽxU� �Sþ��s���x�GC2�����y�	i>qo��;'���_�O�ᴾPS� ����3��Y�gq%��*�#�9,�m%Ah�2�q9�Y�� WhkT�d8�J��0z<`DB+��3.��ۊ��v=9��X��F����dc�`��=�OA���;�B��[�w�:����6cZ��M�+�������c��~�#BBq N�!!����G�1f�+:�M��2����=޳Тs�gsA/L��aϾ�j����'k�B�P�|���9J8�n�=��u][��,E���0,�mum'�Ŗ�K)6~C��V����%��q9���nt�LS>����}<����A9��n/��;����fT�AD�*E�2�񦂚���(oB�}�'O
QJ��w}�;�˦��,}����\�࿤L��Z���˴Z�	3*��EW
J�m�[0h
L�H܍�M� ܟ-uo��S���k������(uW���m�]�3�ZD�Nyge:MU0��~��q�X��c�/��i~��eBlo2yoK*22ić�cR���S���,��6^]'~PqwNE�m��\�NF����K	Ҥy�7�o0�� ���Ճ��̑��X�8s	79jf���N����fCW碮&y埲��+�8t@02��T�S�v�9���:��O����a��֐.�zY����H��)�^��{�렦;x��¦�u���#�#翔�*1�r��!�`f=�h{ &4C<�O;�Z�6q�u��_Ù*�j�����9�{������������,�$�TkI٧�0��咦S���g0���?:�wfϛ\��&����x���)ДLͩG�Ef���@ �~�����gO��T�e�qi��:�����~n�ѱ�.eA!��R;e&
K/��hEp�]r�6��ח4.$�|���,a�E��zeI��oW摺�{/!�@���a}��`RR�䏅�u��%�ƜӼ����R݂4�qm��m��.P��Q��t�E��۰�l�*������\Q��2H�r�+h��!oK�a�^X�J��d�v9뤀"Ƙ�M/�(a�ږ ����$)Z��S^�A��ϱ�����L��9��\���cަi���d?6�xK-?0z:D,�8;�y��bLA��N^;�_0ώ��({X6��}�$2%����Ϲ��T��X�7t����I��c)<����3��,�5R�-�?��0K�M��_�����5.���1���� ^h��: ��]wR��d��k�E�!4�SN+ҭ�������������\�茿PfA�}��=G��ѡ�p;a�5�Gw�Mr'�1&���m��I��hk���u���i��F]Eˉ�)�ź��SO0.���R�;��PT�]AM�Rzn��l��ي���2¥Б8�fr3�̪��v��Ʌ�(f��X� }Jq��M}A�	� meL��7����/]�U��	Xq�\[z�T��Om�6�����7�lь��MԢ1��S��cUF@&�%f&0��{��^�vk
3���v,RɴC��P�0�=ƫ�a��B;�$�,�c{>3��Z�9۵;���6	�j�����Z^�Z��������A�_f�{K�[H}�X9����k�H>%��$����YĮ|z���ӇĬ��`��ᯢ�L.3ك�����$���œ%tOڭ  �A�^2Έ��QO+�c(}@H���Z{̮���9:�{��{�N݈�Э����s6�F��s��L^�i�sڊ1�%�tٖ�D�L��.4LE,�������0Y{���)�r���_���kk`�iP8�[q�Ǚw�����6r3"��D!{���pE�q:�IJ���=:Qҝ�)����F	��\\���i���&͆Ǘ����uم��[�/�	ah}5[�]�e��ג8�Ã���]�p�md����%�n�����=������H֘p+�8��U�"���;�pn����T����C��
>3%hm��d�f�V�g�����|�׬O`eD�4�f�o�Yw�1Mw+7 ��wI���
|=�+��c8�!�G�� �ȐL�xG��`1�~**9uo���N�Z#��C}��ӄu�����7aL$��]U�X`҇����&t�b$��/�u �됀��8��Q��/�v����.�/>���bW���&�ֺ��y�^������M���T��=C��\����-�7B!�5�ˣKb����Z�@�t�BG�����4���/�z�y#4uٍ�A��	��ބ��<޲�+|(�c���E<��Q3���-�����<�<|՛���P��3�Z6����e� �یsF�)��+7����ůxVHCs �#޷�@�^�՘Z�?ª����Yh[}�������H ȯ��6�)^b�7I�W|"o�N�/Ğ�^�6�s��S��|w?��5{�mj8�,�>� ���rm�9��g�al����v�;��ᄚ���,X+iB��B0SY���(6�PD���2���UfX�!Z��ܞ��F(XwDAB�>�%]����:k~��$�#=k�/^~�wIzP�R:s�ȭ4��_B�'\�+6Q��Q�Q�*�/��Ӄ�������[���}R9��Kn�����B��31RI�/
�;�]1�=K�:fgƄ*f`�]�F�$N���u�"j�Z�ǘL���^n�|�f�h-��ÆJ���\@�(��Q�e��֨ڸ��z��[cP��C�8.�+����ﶤ���k��j�8o@*�pNM��Փ*JK�Px��`\e����!&�
6��F)�$݌�Z�T��~U5�YbAS��<�����[eh�烺+�&=��N݇�rש��j���9Z�����ͦ]�Z�6�W���[�g���S�8x�)��V�q�!��[L/�u&����a�(ǖ�!����> _
��C��ƻ#.�D`�<8��9=\����.t��e[)+������h�.��~L���P����{<�c�c�>���ሟ����٬fK�'�/�;��_+��N������U:Δ��gP�Ў4��A���rI����P�@H:"�!���w�C	x�E��ݩ~�� *��F�JG���-�<�Z�&I���D�u\2�8)�)�ҿ��1HD����-7?�v|wxVi��/�KҲ_�#�i՗g����Q��w���O��X}]�s��1�F� >�գ^��gV6��Ҟ5��揤�vV�c<� `���Dޠ��7ϣwli�D��瘵dM� ��6BH��p�gܶ�I?!�"�b�,�<���iF@nR��CbF��B�쯍�v`��&�1S���#-|5�y$:���H���T<Iz\|T<���-��t+H��k���ҥ��^K�����`�<�28�P=o��ˡkbS<v�F��G��Ks���kRG:���Y����YJ�h6b X�v�,�E!!{��'���%�G1�V3U�e��A^X��CUEۦp��N!F~SԄ�sqDq*Ƈ�z㔫�e���eC��H�c\�+�I�Z�N[צq�".-���T����\�.�?�)��%�N�$t���wO�M��Q.���1�'h�&���
����|* jc~�	�<�<$�_b&�8�\����(�R�q�a�ފE���m�a�j�[_���2��F��Gm �:���,GotABr���@�i.m�./|]��w�,o掆޳S{M���Y�4j�F5�UhX/6/=t�U*���̹G��$sI���!Ȩ�μR�`X�N�D��P='���"4�cU��K�kC���A��?HT�2e�F׾>�%_2�ԈƩ��g��w���~�ן,�2+�8Y���c����B�������|X|��tD��D��*���vT�{��ū�!����q6��w���:k%����&s�=
sqA��v<��(��,�*�nʧyD/�D��!xY׌�f�H;I���(z%A��Uf/f%��h��md0���~���A�;���7��Q�Ò�P
Xg�c|o~#��S������3 �����!�r~q���Z�F|� �hJS|��I�#���r$
3�<%;��{(]H��/�������g�E��#3J�XY���l����n�,u�Z��O��˭�*ž������B��ڢ����I�A,F�[�D��q`�-���� bn��WH:H�?�c��׺)�ȥ���9oϒ+��CyL�2FT'�2���,D.��_��	�Q��#�34�4)�7�p6�ʐ4�X&\E]>�r��H#'_�p{��<Yn/�:$����Q�)<�Ť�v�H��%V�� &R�r[~`��E��R[q-l�)�"��S&v�f�F��_g� �6�!fgA���!`"�||zl�&����G�rѸ�"�m���1ʆ/+��~!,����L���f1&����F�2l���*�ȳ��x	R(�O��yb�tNqE�׮G*w"��V �u`W!�,Tݧ"���E��61�;�=�['���a���70n��E��	���H�w�_�L^\�=1��w��(V�_ce�"�&���<C(:���.J��G�v�KO���Gu��U�=�`��|Uo�ZS	�!/&I˲���.�\�ycf�@����{&η�J=W�է,�4�퇀�&)���z�+���N�8E%kA33q=$��4�(��L����LL?�|��1A��c���kˀ���,:}6L`���m�R>�DP�j6�~�#:	����p�%O���2�%g�M�d+��(���a��E�������ӄn#ܐB�4�i���!X"�e��^(%IwGO��wJ�]V�"���
�!2� G݂h�)�D@Ya[l�:z��]�B�;t�2�sA�w�T�й��n-A�j(��KL���͕�����o��g�'�R,2_k$76YK[δf������3�T�hCg�v��r?EA�J;
gTe��4�ǳ��[�3�ƽ����7L��d�N�+�T��P�.�����Fs	(,�F���lB�.9��Ԟh@V�ɨ.@)��ql�bJ�uZ|�_�jތ��B��H�u�q[��G��'@��d��H]IڰK�b��="Ε�9�s��,է�y�EF9�#� �E:�S{��dL��S�����^&�'-�R���)
SS�?�Uw���u)%zOOOE{|�a���Х9��J��k�f�<��_{m��|�O�����:�>��׹Y��E��T��>�j�k���wr܆׫F�poa�����ߨX�o��=!��%A��`5�m�;8��` 	��M����<s:~�^-�����a�s��σ]>?_�]]>�"G��H� ��Gث.�-�}����wc��H3�+�����!�/RC���K{9��Q�º�"!@��̍3b�1���f�
�G�x��w���.��U�P1��\�G��;T9S�wֶD����/����,#�.(�{���}T���@(8��W�X��Cn� !}U���b��K�d�<ѐ<#w@' 0���݉e��'O�w�(;&�T�aY܃,���wQ�!��'���;5�
�����@H�+U_߁;?���󳪨//�Á�3�?͓��!��ON�'F9cR��"�q��ԃf�P��~����*��fi�l8�+t�s�|�DHm=�����g�)��$ҳ���/g�@��9�|���v�oV�v͹.Q�Z(3E &�V7�ur1�|���q�:U}c��=wQY1��X��E�FH�+���]��o��ɡ�P���ו�,�b}{'��D�Lz��zN��������Pi����ð�cH��IDl��|��m�7. ���8��?�$�J=����6��I�;<���9���'�Eo �����o���y��5���X2Hb�~�5��Hs�A����R+� 7���̯h��u��%�'��g5db\B��"b����$ն"(ǒ�dP�	�ZG"�)ӎ�Ȩ=����k�����d�Oz���&�kP�*�..�5kDZ��գy�~�E8Z�[�Bs>�{�ؽ��|%�X@d�(ķ8K�|pwN䭂;li�:%�Q�a�e����lP���뉕,�ө*�j3��V �\Q�[�ϣk Q2�0�W��m~�����О6
������.�∬l��g����#���^���m�ƶ��Eq�':f�w��a*�o�L�(���yq$��*dm��%a�W�c1��\���D*xu���+��#Es�[���L�\�4�l��@M�gj�������g����V��+=�Pn����2Pි;�O5��������Ј p��q&��������&PI�T���c�V�EJM�X�v�
|���Ԕ�VH�f��u�+��mY.�v�wm-�*��?��!��tN�����{J�eh9~gFYe�~UA!bNR�Ĵ�r�
k"���s��(��J�6����U�#[�}B������P���z�_5=�?I�d�	��Y��t�Up�䆑�:��&`��;;�������C���WĦT��Î���[��3�D���^s3���W��{�o��[���_$Y4^#	��a�t� O@���3�I�Q^����v*۶R���p=Y��������tC�jo�d�1�Nk0�����͉�'m��(v����|di��h����+����3�JJ��%h��i(�������_d=v�A*��-o�Vf*1�pY��H�ץ]>z�W�]+gH	Nk�4.���������)8ػ҉_ށh����!�d��8�U�z��DPvEs��Oa#����W�[������x�I:��� 2g���iO|8ʇ�w��2K��Z�a���y�&B9�ы�)u���S��;{��RdnI����P=�X��Ԍ(;/ٰ4f&;t�p��Z�"K����Fal���йX���ͨA�耔*��٤���"ܕ�a����YQ�O�P���9�*�k�F��2���t��X�s�Yn�kL�QO�o2 �M
�>���9���Fg�d��:�y�o�'��HX��|�fOHս���j��O��o�s����`Ģ�p[�4_��o�L�5xc9���P_ZB8��G50Xq%�z#�F���#�F��5�E�4R<-y���^�q�C��J�`C�u���
����-�S��s�ǹ� ����2G�������^k�E���P75�Tf�T�P 35Z@W
?|���o�+� Ft�O�֖��2�b�/�T܍�/�S�
��L_F�T��4Jb��+��~BQ��b*n@�섢0����f�{�qg��q�z\jwW�Er��z����3g��CC_�MJ$v���Z�s{�{��D �et�Ҕ�Ԗ���f՛��k�/�xVo�j�$����g��zJ"�s�6���i���S���'�b��y^���`T�mx�@U;Li�F8ʬ�-�ϣp4��4�����~l���h�"A����N�D1G!0�K=DUWN%-=��RC�k�#���]Ġ� zI����QVO�++��X���U��֦K�2d!~��mD�͡�8�+�Vm��G���[]{�j ,Z�jS$��U}l�)�f%�ܴM��zSؗ(4!�=��Q�O2֊��l�n�x2HN�ͽ,�!��#"���6T��zX	��|��_}�(�I���%|�Eq����s����)Q��u�S 1U��L�K<E��D�i=؟vW��Tk�+em�`�\�2���$G܁�Ű��r���2�|uՂ�E���D��y��d��B�H�|���~���{!�\W/�B�c�ii�'n6�ћB0���[��H���D䳫/��	PIt�b���^*&��G2) @u�?����r(��|7�Ҷ]�V@��O��'�.�&`�6́!U���0*2�J�N
��Zw�v������h:?���16_���0�1h������ő�t=�����g�-5���l1�,���()r6�������"�S��u�R���+dA�W�43�^~�Z��>PSS���B ���$Ecv����T��`�
@��1�� �u;��v�ZO]PA�c6*q�O k1�ޮ��`9x?1����:�#�F:Q���}xO������;f��wK�.'A\��x��tȰ	N�����h�G��L4���Ať���0]��e1�o�?,Hc5��p ��*�m�Ps7�rދ��8�I��Ӡ;i%��O�q3�K�B<��a�{�r�+��� ��}����G�τN�Ae��>���?d���
���/K�j���ox�l�c\2bB�c���=n�j�˴7�DbA��#Py"�<,�h�q._�n��svv���*��(3��eZ���bxB�!���R���bNh�S�v�7E\������N>�(�"{����p
�Y�:��LcE�1�Ԓ�ȅ����ަ�6>�è�����Yٳ��gb���9QyC|���ל�z3#�H"7��Z�&��Etޠ{S="ɟ�m[�oˇ�%G_C�B�O@�`�w�W_�S�/�}��U{���V���.��篚Dy��	���g�EZ8&�p�r� %�@K8�."��!Y}����%�k!�3�]V ���H�w���Uh��@d?��V
�*��y������"��>�8��e+[G���~ChUT:/��[�L�T̋7Vg6҄��#�0�M�ݏ2E6)�U�~�]����>[Cb�p%�˵M(s�
|t/�rqCC]n��=��;oƺ/���J�z4;*�L"V8��v:7(��)Ѿ���R=��&$��T4.�f�����IΚ:o�	�4�O�@��w����(����1j:�]n���.l�f�ط�p���CDYl�!L������.��N��$�\��:t]���0F��g3�#��d$ᐢ3��m��r�����i�;'�?�����t�ڥm�׵k)�b�,ɂ�;M����|J�����U=|�,B����l�q�!8����З��C4��~<�?�m8!_n�O�G����KoKq��4m��*JK��f�7>���f٪�r���M̫�﫷���X?���C �"bN)�r�&�g/?�}�%G-����[��9)�O{�,�-#l�^�!DQ��B��6\ׄ�k%��29^�c:��^�s���o�R����k�-���@w-��@�3CTW�A7*-UФ�<l�y1��E�D?� �.��v�!ȋ�ؔ�����s���y��$A�Ok��ͯ�TzTJr���O��B(<��ypJBAY	�ط?���Hq�ӻ`�~e��������4S�s$�NkMv�{�i�P�%�`B0%"��L�D�=�,{P�����b���p&/h�`r	�ta�I��$N;����<�o����,����o*�cN�8OG��$	�W�]�#��9t	*Џ��+�+��:tKű�3���ts�� �w�n��5�c�w�D�:���*W䟯34 w��b�
�'k1��� Q\s�rAL�
����aíW����|Y��$n<��/} ��T]$�- ��fh���6�W�ha�Å�1ܼ^H��x�wiK�_��ߕ�R�!�v�:�L�����o��P%Jd,%�����P8�� �E�fV��Q'CAi]
ÈV䁘��"��:uK�o���6ʝ?}�!z�.sc��� �z��'���/��>��E�d��d�w�p0`2ϔ,�ݚ|�/&fA�����6�;c��J*�瓍�Ä]����>�?��!�uu�����?�Ȟ��c�p�[�>7���
,�~�����	��o���/&�w.��x!�/��d$kq9���x�87�o��ి6�N �"�'��A��� ^���̠M�J�r>�9)���I�9ݪ�C:yf>Φѥ	��:pDK��w����gƔ(u�\��^�) �Rt͒����m_�H�Ɖ��� j�����]�����,��s���xq4걳'2^/d��f1m�,�b���!�[��ct�f� �� ���"�[����ó߸N������1�*g�]����R�s���ľ���ӞMֻϑcgN��U���<���Q�]�{��ڏ��5ul��ܽ�E��Sne>a+>`��S�ՇX���~�`G*�ͧ�
.ɞ�M��G��v����l����k�5Q[�I5���i�Y4	��H�8q\c���e�Fۚ<�KՆ5���W��k�k5r5x~1��ΐ:D�v��'�яa9W��D���S����v�6��~=��b�p<D�j6;�zb��/��X��O�������p �-��f�!�݋ wU�$:#١m/��Θ��&�xE 'i/Y
�M�w��j�1�2���D�߷NG�~��k��P����ȱR.e-sAL�7w�$d�����ii+Ahb�̃W�u!�+��N滻���y
 ]qJO��E}1P�jj���,�)8զ}�!���Ƈ�B����$�Y##f�V~�3�Ӻ�o�#�����,z\�J���D������mǻ豀1Li6�C���8�WT[j듴�"�?���Нc*��*�V��QwF˅F���XB�����l�z�2���N�Ώ�ո�� �s�:�M�b�����&H6�)�d��7�ۡ#�|�r�LГ4��� Gh��r�!m3aiɥ^�"� "�ω��n2���,�G۰�BU¡
����k	 Ox��5����,ĥO�7u(1*��Z�C6�I���M]��\��f3~#Uq$�5��x5�.��lTo��/��o�kHׄx�Z�~�7�r�)D�2EC(�a�g�.9����
��n������ge$b�m�>^H�˾ק��HOF�P�Kv;�U ��*m𚼎k�!����@V^5bv���E�N�瘇��RNa�.��Iz�'��iJ[�\�j)��#�������R�d>ɶ~+i5
[���U����o�w֢�)H�P�F�~1k/7�nO��H�>[��BLt����E��몤Mx?����0[��O��;���1��^�vH���gKܠ��{�&�w}�t�Px�.������UgFh9c�LS�B��X���m��L���ʄt���l��$a�Ŷ�ӎ1�W'��i!�x�Ќ҄��w�s��)>�T�O3�R����>��=4y��g���d��������ɾ>'�&��i�k�2�PS��{���3�V����( ��{��G���N��Ȇ�9?�@yrU�>`�M�	r������A�@�V|�S�՞ '���_��xZ��jL��O�h��`^<0�B�F�d�5��n~׏�i��t&S����-�Im�3�l`�<-iD�+1T��ov����эN���H�Tk��X��i��P�!�Y��<�I%0��o�_��(9�4Mv5�o68F	̕*�S2��a�攢i����rqݧx�zO��?�wR����i���������.j><��ÚG�@�8���_�"�7(�+�
;@�*���G�'���hv��Q��`�W6���_�Q-G��Y��D�Tmo{�S���Ń��+W�,�t�"|'�87�ɣ��_7Q�
�rˬ�y�u�$&��V�������2/� 1��'��kq�1D.��� $����h��"�Gϫd;IM���� ;��@�˲Sp$�?aPZ^+���V�uD���V�=ǚ_4�q�"Ym1:��0F1ނ��p8�g��!�h����=��"!�䣓oI������	d㾞y�e�D�H�0�YK����{��e���UBL]�\ju��� ��W�������w�N,�D������ߓ��BG9��p^�r��(��^�X�kL�@��9��O4K�9��� �����r����(��@��A�1��9����y�_X�#�A�2(�1���pv�w*_�WU��Ϲ/Ȅ]p�K\��
�ZO�nL�M�c,���jH~�g�L�&��О4c5�2Y6���.�P@��&]e`>��t��;��.P�AA� �@z�D�R&@�=M��u��w`���Ed��P1]����W�=�4�����Ƽ�hW^���-ݍ3Xs������`���iy~�'���@Fw�WYܵ�CA�ĝ/��<O��r<uX�s<�����L#�ReT�D�����Z��E�suf{�&g�\F�����wr+�Ё�C�)T���1A]��w�EBTI4�(�bi;�/�ꃃ9{�繕9n!d�]���p*��{m�X�^,�
t�Bs�^Y�!/�����_{Z���h�������C�S�M���*��2��YTP��1�E!1�ܥ/O&�>H53�tmcI���G�X��m�� ̒�'-��؉3����d��`U�`F�Fa�.a-����+%��$FڏHK0lД٪�,X��ғ�I�'�l+%6�|p^��=�1� 6�V������[*�b��]H���cJ�7L[�U���=Wʓ�髆*�'��o�˾$W ��+K��ڪ�\ۡYf mmq�ںUX/�)����w,�+�70�J��H�h�[z��{�S�iR�-�ICsH\��nz�|�|}���c�ߨ)�V�� y�O��s}J��iy����`č/��rH�?z��?���G=1��� yR�Ե^nG�a,�ت}�I���B�LƲ����ǫ5\9�|��W�1f�5�ݨcY�_Z� ����D'�D<y���hv�l�=W/?�>r�i:J�t�9`�$.�u�H��������*z�=��� Sr�n�OW ��d�!�~lo	�ޙ��z+�%��eO�����l#5�<!�u�҅|��S�!Y�}��d�o�?X�I�MN;��'N��!��r�ԧ0��SG��5�k���s���:=�b��|m���s���VW۝�zW��l�\���T���?�x,,d;L����'��/�O���>>��p�]PE5:��w*	r��b����'���Im"�9v��7p�&�b��g��j�����R\w�C�������a�1$�DD��bF�2��{ɡ@Zu�!�he��a(�8h��z\>��͡��\Ђ�16ł1��Ē�g�"8E�x����C-˄�js������',�4�ӧ��p&jI:�<���5j���AOY�����=���U��Y���.[-��Y�hw���k�]������B�'�{�+R�$4;51�(k�� ���;�x��Z�Uv�⽠�^�	V�u�H#�5��7EЎ+:*�p�k�$�����s�V��!%�ȩ�L{}�N�IdI�Q��bC��z��[��q껸F�G�E2��;�C�w�'��<68 ���v�xW��<��6:nS��k~�%s�.�b/$�2�U�Tyq��-[�a�^�N��ӏ]����>tw�4pd[����9d�َҭ;"�J%�0o��ײ�.U[p�U��t�g�P���b�r�����B��Svկ���K"�P��Btuu�'��(&c(�z��,����¥n�ܴ���{���>K��m����>����c��D+s�NAy
]�!�h2/<-N��j�A���t����r.�>�QΠ3�2�R��xI��oQ���O��
hi����(*��W�r��\�f\�Qs�wWW�(|� l�n`�a�r<��X�*�����Fߗ�s�+{�c���㤇���zj�M��_��m&�Xv4Qx��ސ�HC�*��O�0�0'+�d�\c8	'q	]���{�~���F)��e�F�� �<��v��W^�p��Iޫ%�����h��B�IWM��h���B��\4��������,�E�0e��c{�n�F�*�;�N̈�t��%�jXA�O�`_�H&U���[�[�O����o[Q�tռ��J&&�q�Jc�+r�oo�M������H!@���/�r��-_��>�Ӿ6�c������k�Z�I��6u����Q����w�������er2����
M���+w��H�,/���:�������w�%��*z�P�[ك�h
j����Ԏq �����чT�ɿ�B4�q�y����0b��k�k9Mˬ���Nv�z#˪C���<�En�����
SV��t��Z؅_لRN��jf3���9���;�3�ZL���۱*r{jӹAq������#��l�3��Հ�}Db}gRK��N�w�ǝ�A�}r�����:�Noֶv��12��5�r������(�u���ih���ƨ"�z�GJ����2���^%"P�U0�<��e)���%$-]q~���4���$E�ì� 7r�(6�\*V���T|��{;=�!K�ms��aT�uw[�=�D�ez-�0i�����V����#��-�y�gw�[s��&PQ)��.��6?�:Z�2?�����_�L�~ݱ���9�"$�r��H�}@L�rHYm���~�c��A�1
V��0��Y��=���h6ˆ ��t���o�F�*�g�mϙyM܇�N�@������	�Nя4B�}�V��L�6"Y��:8�>�"�qYȒ��5"0�K��.�Lu�s� w�y;]qK&�9�1���y�(Җ98W��2V��))����a�fY�XM�Ws.��I�%��R+OT�[o7�I�F_��XC���pʒ�a���7�tv;�AV���L9b'���	��t�t��C��l�a��!$��Dc� �M��6�d�w�4��3���[���<�m�*�&6���uh�h�L�c�!Ȍ�ɺ���9hn�T�Ra���A���7I�� "��k�a�`W(Ư��n .YpD��<�o��u9S���E�-��H�N�Ί����[0�@{�}	���c�5���w���ԓ�.aN���jT|�7�}���[#�*���(��8���x���3�n������=O т+�����k(����Vjl��t8IF~��͡��l�J�n�D��E�4�Y��Q$:	����}�"Aq�F�f����k|I/�])�k/>���������_Hٵ���*s�bt��� �2^aU�'��x!�ٌ���⭞���By�1�Ik?qzcf���v�)�y� ��&��8x�yeP̿�()��Zk:�\�s�]�'��	������.�^��d!���^�!q�;�Qo��Ge��L���&�]�6�֧^�^��{��� ����L^%P��y7� ��kɁ��"��)���&��.%V�d{#��֌��d.�.�L�L`;�.U�Nr4or��C�k��#elJ(y`�pVJ��3�L*��\u/aG�|2����Bd�a�N�4ꇛ2�ч�t��`�w2$��Z+^�d_lg�yD@��G���ɐ� �>չY+;@s���:�	e>�v��z]8��`�"��ziz�{�;n11S�ص���(Z4#�:9��TQ冟�6B�������Dm�o��O!�ۨ����	���@I��2�D�Ei<���I)#_9��Ϙ�|�JJ7�O��t�/���\��-�c��t�OF��0>�b�F97H	ǻ�`&źH�5�Z�=�0Cc�����C�8�,�c~��|����7~���@b������X\R��!ȇǐ�wGH��'�f�t��>J�(�}�B@3��Ve�x�O~����2%������لCj�$�Z�<�	�� VL�鱫����ڛ|I��������?���@�
S���]A'�И`����'Sc�Ŗ{q¦�;k�j�"zVi[M<�N�U�bt��Q9�+\0��V[6��+:y/6v�	'Q�<@�"�����q��S��G(�)0�/����@���JI��˸4�<Rqt����տ*zά��F������Ͻ��_��2�!-6��t<*U)^��u_5.Ip��Rt�(8�� ����;�`�IQ��i� �95�o 3�;��ak�Ep\VU�sڿ ���Nn;d���?�)���6Lp�Ok�v�T�q���]�u�JL��0��5Ny, ����WZ�\h�.v}L��ߡԶ��}�au��J���;
T��=I���p�[�ɧu��FQT�[)���t���c}4L<�x�ikpشW�l�l�
���4ΐ�uMa>Iz�>�I�B�l����ad�Ci;��a~�1ks��a�_�������'bҼYrB�yM������ez�xw㊩��z!���)@'"(�y�J���ʁZ��t5Yf�������8��&�Un��kd�$xx�挣�MsB����
8����W@8���F�/_�2,�r�%���5��hz� �-�$p��d۞ٺ�
��鵷{��?Iz#�xe���Y��;�{�/L�� �Ox��)�5y;�L�uP�O�t8&Z�z���b�����K,��dn�R<���I��jD	콝�K�e���6]v^����b�gn�c�r�҈�l���E���|��Fr����8���� ����]��q������N5Y���߉��*I���,W���/�5��(�W� ��B;m��q����qq7Ŕ�����5��IBo��M��梷sg�b^�Ky8�!�у$�=rԷ�Y�xRV_���<���@�9�!蘜-[�����Z���'wB��C����v��z��:�K����Dy�b�;������
�M)����9�#1{J�	t��W�Ep�;�桰��8"R�"Nu��o�HYZ,�X�
C�B��n������m���Q�9ޞ�v��cx[�{7����HI��uXk��¨!x�u"ꓽo|��H��G�i���/�:�}U�.5jy�G͠P��q��ҹg�~b�`Ne0��u'�I�������:O��7'�,:u��ɇ����:�f�|���E�����)�N�| �O8Q���oz���I��V1k8�Խ㓍;4$�`OrWf�b�W�HxOâ�Ԩ 8��S7�¨"h&���e�z��L��8U@���&�n�/}X����{������n�浙 �"� ��WTmn���|�l�Wq�k��� W6K����7�E���w�6-!���5��FsW������f2�������9,)diϐԲ+��o���IW@CC3�mcB�s����l�y*綥̡S=��W�9K,Dd���π��ɶ�?��pu�rL%�>��8/Q�حwl������l�)Հj�d�*��j�MH/5I*���A��5�0ov����t�$ʗ/�)]�d2�19W�CO���t
�yAcS����(;�[�7�r����:x��Q�Ǐ�
6蒡k�pɄ1�$�f��������k[Dk�䩛���
��r�`�.O�M��S$y���B �gnl�_�bbA0'�A!fDNsEe	˅���|�_K�g6!K�c'�M�1�S�������栎y${��H�+ig���*���6P6lь�q�)~LM(s�^�_��s�Xz���y}��)�z����R�VR�Ml{\(�8PX��m�<{i�8$����y��,�/hCҁ@>�9�`2�!��Z]��v.����!���İ4F_���F;���_��<t⎙����E�#�|�Ab����gp
�kJ/
׾�+r=:���+�I�f^��'�Υ(��d�Cz�3%�}ij�a4��漈��l�E�oמ�5ޝ?h����⫂$�?��Em�;��t;��PyyGK�:�밯0��4��D�u�KG����XW� 	���Ɓ7 �աA�N��ZZ�o`B�kϹm[V��Uঀ������0]tԣ!e�r��P����52���M=I$�P7Yb�itJ�9�x�?dO-^�vU�dD���p�a����n߃\,OY�I�����SE5�	QL�N���N��yO%܍�#���<��>�
%L<��߾@{�JL�Z���8O7���.���rV��b��@TS���jC3�cyuu����l��ڷ)/P��E�ԧ00[��W\������#��P�����0T�_��+�ha�E�>���x�a	]��p-wP�q�g4t���� س�H��ӱ�7�5S�h�':�]�Ml���)��"��}D ��s�@�	��;��W^0a� �u��f�j��M��A��O?����B�>�DU�Ԡ�IMƹ�me�ֲ���)�lD���mN��]�� i��27�	�R��'8ZB� ��T/��~3<ؼ�?n�:ԙ����?o�n�$ΩH\xo��b��Lڟ������|�D��|n��Ձ�[�#� �m��'?����T�ꯈ1}A�
`�P*�a���Aɺ��[,ۯ�j#��W����E�Yz�-m�<		��a��shⰊZ{��F� ��J2ךT�(�陪]���Y�Ϧ�5G�+e;�sX|����Z�����=؅���6yX�.�q���e~RV"�k�ӭ=�����Z���ak�f	�v-�kh��^<�|k\-D�b`�"�e�
bќq�I��r��z"�5�"@A���|i�ӻ����!¬�9܎X_� ���`��+1Ը�W#e�Gf��NJ�]��my�.2Yf�����%��{�@�U��{�J�6�1Pr2)t�����=�+��-�gh^Rc��a�lCj.Þ\*1�V�㙤����/F�C���Ɏ�� G�F�����U+��I%����X֙ޜ�=��ڵc�'
��\2�����
&/�r��Y��r�\U��"����mSY�}�\:�1݌Y<մ�MI�oP�Ga�ǅ�Rw�u�|h�i�q�.m�A����P�;�a�_"�
���
��3Os��,У��dd���w��=�m���WE	�%���	u�K�a-E�4[�������b���`w�jQ���]��!�����jtV�L�n�3ƥ,��R�K���l��'�E�	�I�9M/��q0�ʂ���Z�_*w6�S�=N!�yDH�ژ~��$��>��'��ҕ<����Z^,g0cF�������dC�
�jr'���5
�a�����jȒ�������x�꼣+V��,�낓Q�
c6��s2$d���g��5ְ� ����x_���c�C8=������A���7?�E�
��M���jҩ���\�t����� ܈Ės��`�s���֒�m_��]���E:�u������2�)�� DB���t�H�p�ql��N�U�&a���W�9�2���_�l%quԝp-�&��0�@_�o���19"���Í�6$<�����\�I�>[n9��r&� `_���IB�����d&��%,�ܷx�uװb�aO��;;���]O4��h��(�ɈL�s�j���n�D�e~�c�� g�K�#�����J��5�g��0@�:���r%X*��\�i���,�8�+Zu��;�+�� ��=�`����G��Yur<O��Osx��s.��
Twܦ~� ��[���؝�MqE��0��r�5R~^�V��ޜ�!/�:o�T����@q�h��oV�=��@@D񏣞��w���H�Zn�M4���BY�9l��$�+9I�0�S+�[����}U��H�]���,lHq�b�����Փ.�N)n�Ŕ�v�z����@�]zc�(�bA%�9�gt73
zr�nTwt��9*��u�����,V5�/5�G�n"�Y�\��k�*evh�NPB��KSJNC�������8Z�y�$6F��i���q�!���FcF�KfzU��(�N�l�E����t���c���e�J[�f�^&�L�r,.�I�ܬvM���u�)������wھD��sݾ�zϺA�{��i s��K�ދ��-�@X�����'b��	3���P�F�kr:��,*, ��b�3��<�P��p�8ui�[?Om7+��7U�ޔ��s��������́_*q���D��?t�6��Oޡ��h�6	G����Г�=/�����G�*81#�>u/���9)]��:y����6*)CIqJ;݌3t��]����]8rha����.����yZ�e���yuo�7JI�r" ��avog	\&�b{kr/��h�fj"aܶwZ$tCD真���š��G3Ʀ�1R5�ӔG\ȹg�&@�`��9�c���\[�%r�������ʵ�� (��W��4NL�Eb�w���{�HX+_��s����b���<g~,����E�d���,�@G�ͥ�;Ɏf\�ڬ^@��9��H��fd9��a`4w��~��R�r�$$�r�?&ŮD����_9X�-�󢸗D-�s�z���-���;BV��^paǜ�m��[�+�ioK)͋/5C�#%j��.Fh��Ws�KbK:q���J��aZ>uY�������T�S55$9"���*NC�F��s�׬ - ��{t Y�X�+�Տ��q|�r	׵���Y�75N�j������܉���%�7��#��8��nJ��m�5�K��X�t}>��3��p.�n�#Ej̏����βY��&�;}6O	�R(�1��.8�f�nunByE�S༧��/[+�2�W���`�5�'�MH��@�~�ۓ8b`+x�M��H�t��FԴ�L�lj�4�������|d|ia-�pT5p�#�ĭ���l���1V���F��U#=�L?�5n�]8:(p�;�Rj#�0��<�s~��u:���� ��c�-�Ǽk�M�%͉FYF�]EJ�y~�H��p�|٭b���Xד[�Ԟt�"��}N�Dȋ�mC�`?��yČ-���/@J�yg���f�G���#��P��7��˻�+mdN$�T!|�[���*��� ���"Q��0�Q=J�%a�qIU����d���;�1y�����t��{�#;4"�%Z��*J�x�h����	K�[���A�e����!N�X��Fw��}�j�o��y�*�y^�{�1��|��Ez��``���U:d��.�|eI�g׵*�̥���X�B�*2�M�+���"뮿�`%�5u`Y�?f:kw]�~]��Ḵi3Z䬃�x-$|��-�+���rpLIB��	n����������Bb���/��L�M�fP���d������y(�{AG�g$�R� ��!.л �xYy8���ڏ*�7�c���098��B~ո��7m�^5�:)814j4&r�9�!Y����`�Q��H��ŝ�Ҧ�O�Y����RIW�Mŭ�����Rc�궻��ht܏!h����+]RxW[5}H���?��F�z�T��-�����P���.��B�/^I>�n#9�l��C]�-K������rﻰZ�	JO��:&��"=a-��es0�k;�u�s.?&�O0�!�Sn�E��Vd��q��תB���h4�u~�[ϽD1m
I�b��b7v��$�:=�w�����Ƶma�ή)���<���A+
� ��1��)A���Mq�C>��]Q>��,k�a�G�+&Y�� \�9��:��%�݀I��i�~4"e����W�F���ǂ�~��j��^��-`z�a%�yS+�NO-�;no}�Κ�D���g�˨��i��,�����Rp ��j�V��lt>�w�[I�#�$� <�����	�ڀ�Q����]M�[��
bC��`s@��(�̃��7W(9�7EI�q&�u8���vto���7�#IQDOS(P�1������S)W�4�n�;|+Ͽ�&�f������K�ܶ�M[Y7K��UOn�h.�����%I\^ g�W�L�ވ�+��1�5�����+��Z
�)r�KS�����9ʲ�W�d�V��`���dG��,�8I�5�nUqy�`����f��^(�|C�G������o^��6�gĈ����<F ���H,c]�c|Z��f��S����ĳ	h���=/7]/��(!y�_;�h6�$�@|%�j�����~/7����yb���f�� s�9^�W6��tT>3Re��'�(&ОYS��	��Z�I��\�&�^�/��<�(��OR��BՆ��"��/!}�U�
(ћ^*RL� X�[p@#��aFn̔�Nu �_si���W���z��6��M��1� �y��8�J�.�(�Ǘ/~?SE���7	��	�n<Y'����W��if̶��&86Ț��A�`:�Tvo��~2H/����9��ؙX���I�O��=4k�Iw��#��'2x/��c�1�h֙�����g�m��1+|@im��\Y����b7��K��	��0#!&�|eG��ᑊ5������j9��X#��|�_$9*�c��e� *��O��.�->Z9�+q(����%,d��O�g]\��&�F��I����<��E#4,ɽ��\�u��o>�qC�����;���,��ߺ�G/�H�Y�O�����&�G���mh(0�=�Do@R$�1"E�X���}5:��ίoF�W���S���
�����|�%�dd�Q�b�����8^��g�$��o���[�9��yG��Q�w�Z���d��<��\H)=莥68�:�9F�67���e"�����o,e�Z�lq���e9l�>vV�������>C��.)����!d��;K�e�c���٪�iX���	�ՙ���z=19)O8����D,%H��/ܛ��Ձ���3���x)�Z(��V2A>���yy_G��<�D�%'Q@B�C!��	�5��0��	E�#Z��6��#�~�W�/F����f$�y!��<����9�m���ך�y�؃����X�P�<^|�ѹ��S3�A:�${��T��w��0r��&�ŽY�T0�O0��R�T��r��=$�a�k?,��)��j�����J�<b�,[KhD*@D+�eqt��a�7�ȝ���� �5�}�]��6�=�T�5�O s�,�D1�7��]��3�i�mi�8���{����J���p�uL�����A�����c�r�W�tA���f�l�!Y���3��ª�]*���
g��A��㪩^�\��܏걸���t
������]��-I'Pr������(�m"��D�]��	�B� �V�vԾ��bb��mg��ʬ�Ft���Q�x=�����c�����fSV�Ϳ��$9j'�/��H��}le��5���"%!t%i$5�6��D��-iK��vOD�1�/�k�d���l�A����3`�t��k�(0�Ԫ)W�5݊��9s�WԿ�|��h[����	|DZ��O�L���N	��F��w��������,�d^����زR�(-9G��h�5���\�O*��J܆V���<,eEM��3��:�%A���=C}��g�]?0�$4^�gj�Ny>p1�֣�9���Ix�/��un���4;HY�i�=IZ)�:��C����R�0��"]8�X �)~Q���q��\�P�;9�����O���;/�{�JW(?��7؉��O��ns��c���;�r~�>����+�Y��e��6?���&�:r��3׭��y��*���\N��B�$v�#��7'6�L��n���9b<�L%��F�n�F1�qnJ����	��c�WR�Ȏx�
�;��K�3����_�W5H���	��G�yz�ӕ��.b��p��`�Q�U&�_b�r�Ӿ�((���I&�0p�`5M;�sJm�,7�Hd��h��J���;�q���� 9��Z�U�n~#o	�3�8���mK%�fC�Z�[t2T�x�k����`_�%���o���A5�зG"�����S�VaVf���*3�=ay!��@gk2t �>������m��+�⏽690B�B:x��7��~޲�zeM9��r�2�@��'��qc��P�-|g�Y�|HVq�(KA��ՠ
�ٛC�喩B���3��������m�b�,pL	�vނ��!���C�wR:���ٙwrn2\�2(�M���4�$���S$�Xa� >]L iK�=ɶ���d/z/]�չ�淵�R3��s|�����|���A���n�?M�;Jo�0rJ�x�d�&��[	��9����h�U�C���H8�mU�-����H)��t���_��I�Xx�WIϒ�;�l��9d`b��+�	c�T��A�KK�SAO��{+Y��"��ޜ���/�=��s!衭�u$�bo�Va뽙>�-�h%	��O~�jG	*{��V�!ԋV:��2s^�\�����'/`��P�����*�	���0�U�Fx�YX���E�"IC��*Ʃ�v�-CF���K�{G�V���0^hỷP)D���"i1�1�'�p�=`������t���\s����_�HM&a�c�=@��76|���-}2z߶:�IA<<�bk�w`ڣY��\v�!��@��<�i0-��2�i��[q�%U_7 8f�� �2`�0_g��^�_�5�Co�d2&�Π���%s2��z�Lu������;�D`/�`�<ܔ�hn_&�ce S]A ��k����^$��0�Y+�ӆ��'X��G����#���j8��Z,e��+Y��Ƞ�#N��U;V �sP��,QO��n	��F�H�#AJ����6�o\���z�*�u�P�����
��9>֋FYS�>�y�8ݳ�|����+T'pA���`���<aPɰmF!_ҨMh�}�\����ܶ(�������2�$���DȾB��z�	�����ăƃ��:����g*�J��c�?Bn��_�R%l�;����X��/�Xр������^�?$��k�Vg�IXԿ��(�Q�$OmۮQ��%�F�C�V��]�}-˵�0��MyF8��- u�?�tu87${�:7��r|��#.V�7�l\h�o�ZC_���+�Y�����+d���
J7	O�+�����k�C�p"��pJ��:�2Fp���\bH�NZiv��<�Ľ{�5�vt:��Q5�VL��E�C=`=���q#�z4�W�R�k�l�|?�����%qhX?v��1�z��
L����]��8O��-�?y��J�%ϯ�d�с7�-C�]�+  ��Y�^>�!
����2�9S�����u!$�$(�wM�q��������ݦ4I�$���~�x��	�N�jF�&�zm��W'j`rϢ��r`/�T`�1;�\�<�zcg� �m���X=r*_]�:h^M,"�M�ȇ��B>�C�S�*�}�Y��"v3,[����mjIQ�ػ�:�>zkܳ�g�J9yFķ��6�[��7��]TݢOOq|7�-D��B���.���D���S���Ƨ�f��Y����N�%��yP2��c�"���~,�F��k�rUZ�o��{;?�{�,��槨p^��Y�2*5�
�g�9#��DQ�%��n5�
��̚�49L��N#����)�-^7�]��W�����UG�5�Ьʦ���c�yD0�]/�N��dȀ�|���o�M���ޙ)�K@�:�������05��["V��`yN�dd䔻S��uޱd�"%C&���ڐ
�2O?���Ѣh6��)����[4�ֶS�b�'=F��-�u�;ճz������M�~xEf��k�9�����|�>Y�<��s�)t'���	)	�v%��}�K˝D��P��ԅ��A>�q�(���\�0v@�����%O0[݉�nǫ<R��S����w1R9Vu�I��=Q�N[��տr�QzJ�������͠�̽���Hm<6i��vm�o�(��ةX�p���^T�.����E-�HK`⛻���a�	v��ԃ���yD�qG/z6S����1�3���y�:�;�+��!�F߾�"O֥���x�UP�-���	�u5��]?"�F���D��#zB����}+yjloFh\#�͚�k{�@G��/,�������,F��\��$��nn@rz��Ʋ.��7i�.-��9d ��hI�
��G{.l_��#��0bC��8]�
��HgWl�:�"�y�{�=H�P�|-V��` pn�y��5�XōT�ڽ��Qr����_u��#�Y����*�6�)�W�AJ�V��՝8��*.̸s�? 7��~_}�O������	I���Xv��>2���-B*�&=�*���iS���ldsc�lV�y��<3Yw�c,����5$yc���$SK����&�NN��G��[�G������'��|��^T.CG\��,��T[5:�}@w P�#뷖T7�yյ�E�:ш��q� �2i^������	��p EqP��Uy:M�>�.�����c'B۷wVQ���e˺�/|�3�H�R^s�L���`Z�RfW�׳
�����W[D�f����
�0\r%�y?��jX��hwp�?n�`�S$��iiT�3&��
ඝuHx`An���������x������#�u��o3
nq"���h��)K�?��6�vy�d\dF3!��M���A\j���F������P�_R#�����zGg���5-M>�-%خr�@l�-���3����8�l�̃9�k����2�lf�@��'�u;�r�qv{p�	����AN�E��P��s๼8XV�3ʥ���4�'qp���K,0�H4�fQ`):|���i�p�2%3���`?q�*�����fx�w�Wq�7�'~BD� ��B���O��b=�fP�'s�����9�݄K|T8�N݄jJT~-��m�#ƏX3���n=��[qi��qxo�<Z����M��O�*5,\w �'u��L�U��^DFGa^p�9��0�'9��N9�'_V�E�N���S� ��h����ͭ�����ʠ7Cѿ�#�P-)H]�2�у�n'�t��R���W�F��N՞���Q�[�/��m���=�U8AZ�I���B�1*VU��;̲�{%�{��%-�b�?��
���Hn[yU�X��L��2L�L����O8X͂ƛ,,,�����ҁ�����1��p��2�������O�+Y��~$4��r'�\O���87r���p��zu�Z�k'\ҟ���5 ���3�����'���24i�6Vk��f�1Z����t��j��o h.��x�-O6M��v�.������~������A�����[������V�R܀`�tا8�@�0��{�Oya(+%�����NRg���6Bf0��� 8s£����N4n���Ll�z�Qt/�S��F�fvD�,�D`�D�z�_93u�⛥�y2x�seG��6\��K�1a�L���^��N���cR���������<oPS�b�����L�\�yYn$�E�
U�c%��0����2�����w�L5��\�"��@�`c���?)�̬�X$F9�3�p�u����b�i�K��#^������5_���q�邜��S ;�k��;�g��Fvi�- �� V�A���Yh��Fܶ�/���:'&mǊ}�PD��.��n�Fh����̓1 �5�ԇ�6���,^�0CZX���3o�a���ұ��D��ZwE��2J�\lv��� p�sF8���|kQ��Ǣ����_:�F�O��2��`g����&5�i��iᶻ)�m�-�Rl-��}3/^�Pt	��ֆ��1�GJ�����X~������ȰH�cx��U��#�%c� `��KM����7�yԋ�uY
C�V� ���&ݛG���+O�
�F�ֽ*���u1�2{�wʥJA~�6���b�:@T-����b��O��7�����R����v$��s99BWĪ�gaM*uɻ��k����@Z&�ުB��ޝ������c�A��7�t�����Qߛf���K�艨 �㇌͒^᥂^���I���g����x�g�^ �a�Lѧu�:�P��P�E��q�Ycvf ��ϻ�I��GF���W�ڏ5gEv�󂡽��NI��R2 ?p�O'�d }����4f�3m�	F� C���oO࠰�g���F��[��hAg������O�j���w����r���ۆ�4��5�qi�����_Yp���9,���m�!�	��i�$bg�E}.������/�נ�Rg"n�DwľddbХ B����ئ'��g�@Z�Bi�]�bw��h"N��V$+w/5=�T�[��m���^�LHC
U��j `����/m�<7q0�8Dݑj�4ȵ"}�_��]��fd�8��m��3Xk�{ҁ8c�������Ǚ�9r��Ӂ��A�j���5�0T	W�p2:�
����vb����j_��\qOc�r,�VK�Z*�Bd璷LR2�ڮ�6Jo��+��|(&�e�x?��n\�R��M�|J�7���uy륓w��j��(����9\�D���ّ�#z|��s��$q���j �6�\%}��� :Vd�V�z�[�ֶ��pA�%��s�_q��S��M�\� |����<����.̺����5��r!_'T��k�F��`��B�B�&�=~%{递�j��v䦯{i�塖~�mp��车�6c9�\/����V���\��;��.�-� ł���:.܏&n>�0-~ka��]M\9���	,q����nǝS�J�."L����E#�7�6�#�
}�>��2����ecݏ�I�o5�Gx���x\P���g�R�4�h���^Au��#%�v ���l@���s��U����}yg�F�HQ�&p�d��ݧ���Lj�!�˙�g&.���k��МE���Z�\|��j> �<�'�|�[oh�X����+�� )�Oڮ����YM���:))/uJ��l��CM�w*1�l�r�P^*˯UJOJH:#�=E9;�e�
�G{.3�#.%OI�Fl�G��%��[��7�ϥĘ��6_bՎ��\���Z�vǟ.���@X�~���_��.&���[֛�U�\�>�ݵO������l��8Ç.�h��m�+�Yy���n�5�Tx_�DNZ�C�\%e��^��ALa�� �I4C?Vm2���O1�<S��(/zy:���J�uׁ�>���>�äI��QXg2��W��,��
���C��z����9/��c ٥��2��2�@�<��?:}P�!�@u��(���$���&�� �����ֻl9��EO�pcH��(y�0��Fʼ�r�L&�-_!�]N�K��uO�|IZM�:���b�a�k}Ŵ�&���	y1�?�[E����lz��#���m���1�4 �����K��ik�M_q�|�]ەJ�h��o�\��[������TR�>Ȩ3�H��f�yAn$�c����7U2EZ1���� ��s;3?�0B��*m;|^��k��n������@���R~�W^Lm��Y4��a�
�H�n�+���]���3JxD��<f:v1�LJyܕ'+-~ֈw���N4�p�@بף�R�r2�F����+�*u�;�dU��I=&>������.��
R/~|���OAY��]��P�GJ��k��:���cڌm����xk�C�� �c�^q���?g?����� ���y��މ�U�2��V��{ʐ�ڄ���oI�'i��4K�X
�	�����M����XGk�7k���*� g�1��	j����n�p0</.��)��}/�9��5e����Ŗ/,��*��7�P=)�3���\Ȧ�琢A�1���D#��{��ξ� ��Q�S�7{3�%h~ʠז�/]R� �.�p ʖ��s9oL�Db+���q�c9;8�p wE��0#���3�S��Z욉��4n*��&Aa<��j=Ns-I^�[g(ݚ�5(.�$m���GSg"blzY����SAc�O��vI2����=ÅJV��E:%4|��w:d�NX!�&eM'3}�|m{{p}R�,H��E�D͎Bs���Q�H�N%�[��f6e=�_�ncT�܏gv�Q-AG3�����)ؽƚt����ol-s]Px�!�V{\w�.�2S��� u���c���gDasE�5o�o��e,]�پX�
����@�#�*h��H�ìa��q�Iٰ������s��>��A �I�ھb)z��E�T�6�k U(�@R@��5u>���$�~����|�?����P'��[�O"|��hê��&��m��\�h��r�؃�C�vͬr(�Ktih�r;�j��%[�|X�FɄ�U";�!�yJ5�������~��m �׌�����8�4~�L�`� �k9�`��:NY����o�M�������."�R�e�$*��Jk�|[mň;�؍�;���&�0N��lQԭ�zטf����[{:��/�"r��d�`��@R�"���d}+w����D�ﶷs,F����Х#�g������1�h�6"�Z��2 HJ/��3ߕ��)�7>�+_5��r��܄pb:� �5����Y+c�֥����R���֜�Uso� h�=��=�#z��d$�T�Z���L�2ɒl~J'�7�.l��j��f~_l��}���DlfL6�±݅����h�v��0̆��9��{�ں-�H�"SmSfw)3N���Lz}�ev���2��!J�"���e����sc3"�麱�bEb��|;�$7�=o����̺7wʶ��nh�W6.Ly�N�I:������5Op�\�*9݂<£���bڿ�]�.2!S*�A��]XXC�:��3��K�� ���@�˨t�/�H�a2)�#���j~�b"�j+Q�� Ƶp��>���F*�<y$��<F8@.w���{�@�ٻ��b�E���?V�W�py��4���P�����	W���0~d.e[*��JZ�7>����tooK���Nk�Et>S�c/�L�L�����C�331[u �ر��sc�f�j#����s�׃�뫀��î��]c�Rw������!<���ֳ>R7#���c�q���Q�_hE�R1�>�����ʣ` A�%�޹?-��JX���$h��9>��GhE߾.���*7 Q<$D��2M������6�&gJ�ƎG�P��'�+�JߣR����p4l3��e �-Ct܋�5��R�H����G}ܩ��'U��	V,e��	;L�S�>���OD(�x�`QL��{���	���K��<�A�aa��v�o�UC���3�؝�.� �ħq�n��������g�҂��XbxŭngC_�l��Tk��+��+�<]�����J�2�`N���t&���lLR��gP1&���b�R�l���>����/�� �}�F�Q��Z��1�%N���pY�N"��w�	g�������-��繿�^���|W�uO�7[W�䣇a߫�s��y��.ShL�8a[�ϻ+rm�tT%3;j�ׁ��q���RM+�
-@��B�` ��;~��0S���M��%��nIן(Q]�Px�T���0Х���I���x%��t|�6���m�J�f��7eя\�u1���!�ïb�h�	L��3\ ~�D�~N!:����}����׺���G�Jw|5�i�mG8����Bz�]1Ǻ����20<tC���_|�+�Htw�^pH�����prV�&�Y?9�/gBa��(���`'|���0Y �p5|� ҟ�YP��|Z}T�|�[��5�o�h2�	���a�a�e$��Z�b/q����%�[�x��|6�)9�-2�`[
Y��Ό�T�Ĭ(�ޢ���Q�KEM�麼�[��A@�F���Tl��o7�	cIu�����o	Y�T3̭/�'k�RBU"5��������Gɪl�E���
'�
�l��"�Ab�q����0�� ?�}�T�#
��&��h����C*�g^��qE)���3*����x�ܐ0�ϥ{D���q�p��n�;	J���� �
��P=Ɛ^g'0X��	���m�\�>ԅjFJ)���LMp��Dz��Di����y<�ק3Ww|��i�vP�<$�۳Nr��wH"�A�?���t�w~�v���|A���e��k�B�e�+K>z���e+��a�=V���7�*�5[���PL-5��l��d|c����*�g��TA_(!��I1_IBG�8̅�f;'��_��$$[|����6hzD<9�"��5�ꍇ��e#E�G@�F}����$��A콰�M����9z82ZU�!��[Y(��
��=^�$�ݑ�����J�Z�(Se:U��^��O���(ʞ��/%񯅍 Yʕ-��	����k�&#�#3\��Wy�+6�^�F�R/�r�_��A��������3�*G�Uk���HV���ID����̶��c�O�X@�-4��=���|O����Ϫz��֬����y�&�cl1�/lD8VZ�ZcG�THr4���S�M}_�0���|��%�>H���	I��4�w�$| �����"jJƴ\�y��M�����7EF��+�Ugk�X�R*�u0u�8�ؖ0L7�)��n�I�^����&=*�i�����)tj }�}�{8$SP.��r#�'*�������PX���ఙ(�M�Q@IH����9����� �J�Mc�nN0�f��.��_��R�����w�a�k ���r��4�8x�&%i?s?�V(ٝ��)/?�$يh2�հ��,��끷�a,J�eD�%����Vw�?������ֆM����ƙ�V2=�a�\�ȩ�8���?�F���i(t^Wꊒ����O~�6'W��"���fAp+���^�t��M�*\B��S�ѓF76z�UP���c%[*i��^��I���-�g2�Mv���s��e,Ar�!ղAyD[�Z2��WW�$l�H���7Z²$-��}Z��cg���Zϳ�
�����k2Z�$q�@׽�^E�y��U*�U��~�r�"$2�j�b�1����7��$�vc�
  � )��W��k�[������5�����f���5����̭�I���Q�]w>�M�-?�$�9/=F��N�脰��8�WfFx^O�*�ɫ%V�"1��@p�Y��X�:{���S;�/��i��o
6�}Gc�p`E�HX4�1L�����;��~���}Qo��cҹb�����!����~v�%A3A���~0V������ ʺ�D	�ʃ�������ԨtIC˝ܿ�o�.7@y����c{� Q��̲�Td�W���{�>cN0a�dn������ll�<�Z}KI���:㑆�G�4ʩ  8�p?������Js�)�F�J�(����=po�ף,*��c��]��� EK��ԑC'UQ7"|x2��}�`��&1�I���oJ*(�x�)���>Z��R�Ug}�H�A�%�'�M1i��$�-�J0[��OZ�o�6p*�] z��s��FP������ڌ����E�|s$�%�ג{YJ5`��9j�.B�2�*���� a��PRI5'ÂL���U�7���āO>)]_s�]wS���!h�)p ��АK�:�B��V��C���Y�ŗ�DT=X�$S�a~��TsY"��Ǚڝº�(}�睩��E�;�
���æ�� 膳�䁁WE�ɷ�ګn�9��� a�ɗB\�y[�6�x� �n�$��]�9��ӣ�l��\+��C�aY�� 5K�|����V�{4���� �:O6�v��ESb����a��Y����o�plD���ԟd�&�C�m��K;�`�B3$� ��'���q,��I�}���W��q�W�#�".	��ES�J��	��<��O�ZaM��g^�O��7-�O(]5�����,��.���#��*��y��?�r��`���_��z��ץ0ō���M9����k2�v�,��B ���y�PGc��li�Fb�9H/��� �!R$�+�d�
7��&S��8\);���E���W�WV�]R������ndt�6��5�g������o��{�CZ�7& 7� -��oj�|*	(��>Ï���
%��V
C��b�Ż#Y6�`������@G�XP�q�1��4�iؾl�@4�Zz}�����?Z��3�\cj��Y�z����X�} �/E;�\i|���-I�/�g��m�{���bI�)�d���5��?^�L*RY��~�&��CQG���Z�^.�r4(;�*��eQ�1�N�C��������8r��a������Z����!�d�ۜџJM�s5^�t7�[h�w��-� lx��S�q��MQ��a�4=���1Y�,����*����iǢ|<<��Y4����� S���S����A��S�I��\�칁+p\'�0�&�������\u�8�#+�?��I�����\@��t2ho�����ؗ�>���*c���W�5���'5��Y i�m�2�={��AWؓ���_`F(0�(O	0�Jm�$��"iA�T+��qQ�t�]>�n8��3����Fzp�T%�LΔU-��T3���<D𛪫�����P��+v{�B�o���t����}'L���z���� �
?��c�F|�9��/mi05�G#���/�\��^K��롬�9�!֎�$���;�n��U8�+�F��t톴�j$<U�TꙌ�͜X��tڒ'+�,3d
>-��+s+����c(ʢ�Q)#I��� �N�`�!&���T����tx�� $�����<��L��o�A��l��;��z.��ƺ�T�2�W�E\��G����q�� ��k���m��C92$��ѫ��-�!ѿ׌)���� �p���Ix ����Oo�X���M�8��ۘ����*�ǧ�i?�$f9�ѝ��=F�㲀6rA0!H��=b����0+�my/x�~�n�b凯4��V�[�g/��јvH��v�wt)b��:FsGq܅U�0f�DW�*���0ޛ�(�2)�@{�cG���/��������-�?_�A���CW���$���O��}����(E4.�13)������Uy��~iҁ̕(4B'�W�S=^����ɲm dG��|�]�A[�b4�Ǒ���K� ��1�&k�E��E��Ԍ�I6�̀��y��A��7�k�w�S�����"C����}T~l�i�+��^�P[G(�<���I���l-��XL�+v==�c]���̓��V̵3�|���y>��6-�̼Fv��'�t��h�e��:��$Gy;J��� ���&v5W7��=i�_�%Qw$��V� A������~g���}�r��1�+�`1���7СaN�[h�z���#7�B�����!�� ��,N�u4�dR3,+mX5���^^�D� c|Q9}ffw�PՆ���xf�����u@�QO�@�_S�~�����#z�j"
�	�/#�Ǚ�T�V���
�Ú���T|_�S�}����:P�J2H����p֛[$9��kHU%\���J����~���6�Uj�v ��L"���-͖��������6e�l���-���=��y���#Y}Þ�����[,֐�!��e����]\L��N�TK.k�Ȍ�2�wiZ���{��̾�O��Ս�WS������Fy�i�~��@�G�;ͲM���x/Q���m&�،�S��z�kY�k�.���%��hR��3�Ν������IX,� 7�U[��Mx޻����f&��������� �_�hUą����!P#}��
�J����ĥ�Y+��k�w?�̨����.ϺL��?ku��S�a������N�[���������'�o�w$V�?���.dmz��=>.sp�8�N�GD���p���4��<1�</N3��Zi;wJ�iCb��de��Wjy-y���Y���fj�cof.]���v6�=������x�[1�2(=i���/E�4�����T6�G���M�瘃����Y��z���mJ�ݕfq~�M���pIA��g���?lN��i�TS��ב���Z�>�CpZ&����Z�h#�Wݮ����&Ǘi;��`jo��՞�)�ܼՌ�0���k�������E�bT� ;��*:��k�T�v���w^���(�)�ŘI���1�,#fSh<����z�ou% ƀ�$���.��5�r8���A��mc���ur���W?���b���HPF����K�NT�ګ,a"��j�?
�9v��'-_5J�_�K������ e��^���ǥX�O+��5"�I$�l`�Fb��$�*�_|�_(KEY�,�ƭ���o�~��Z����ԥ�0�X�T�{�q��Z�P��m���_a�t��vmފHp�%��I���8 h���Bn�z�[�v�}08N��P^�?�z�����M�:V	�?ͨ�;-��;U�$P���,e�oH�8�M��,��{�?i��)C5C�843d�)1�����x�����7��8n4:�� ��'}�cQ@B�e�����8;�_�������Y�plA��Ј�/ '5�n���%{�c��
�(�V�(E�ә=�	;�ښ
���X1�n+�+q���_Ze�'g��eݗ���8��B������b��>�:C�]��'CB�q���f���'k��:���P��
�{���ǯ����	�"��0��Gm�
��)��]&�H#]5�����\�"��&��B0����tߤy�\QN~_�[rp�W�< ]��%xiϞ���.̟[�Ҿ��Ѱ?�%�o��Z�{�<�k�o���'ͮ�<����a�6����f|����d�p��^��1JUh+k�8p�Ŧ)�8�Q�}���v/����&i����![����hl�Nr�I�c��{�6.�*h�]��	��O���秢p�V�v����J�l�Cm�2{����|Ǝy�~Nv��Tj�pry��)x��yw��VSex��
�i�(A���4�ȣ*[���,�s
��a�:���v
ޔ��%�S�u�ܟ�����%'��|Wvo�k�$����m�'/�
��%=r�Bydl-D� ��w�v^��sc�_޲��E;t�����٫C t��~#��}�h7zJQ���9kz΂=�i�(�j���7ߊ��35V,����*���No|� �����%y ���
�.�.���E�x�1�][�Z����K�٨3��W��7��J,	ߢa/d�iE�n-~D)~k�t�d
�#�%N��*�ؘI����P�G��-��٩Z��ޗ�G0x���TKG[��*��|v� �P�I�0�t�]��s�e�=���୉Ŝ�%��J�����c���� ƅO$ھ��](jE�Ӌ���V�&�臾鬨�*p�;�o�vdcp%�IťpO�!�c)�U]�A�Ƥq��ݮ��H�G��U1�)�c�=��U�W��#�=��I��}��VL���|w��x������+S�JR�CuP� S�gP���g�I�N�I�&�_�7� "�0�2��O�p�D�����5���[�A
��<�7�z�F���1�).��OMM?n������ے?|У�L�1����s��QjZ���^�k~��g��b���,Ay�o�M⢵��>6;xR�i�X�����_s:��]pǝ��ZyX�P	�
�^��X�z��l.�2Z��юI�&���U���	v2տ	D��Rq'8�kp��t��i��T��� [C�D�/�@��4`�*�W1�˶��4ّL*��Y��ӱ��М�=���9�
S0\_ݹ�ڻ�m^�)�Ƌ;Fn��!ed����ѩt�\u#�N�7�|ۀF����p��9p����)I��M�0U����󩋝�ȷO�D��D�������!Vpwf�Z3��4��+y�^�����[�̌�O����G��i�A��]c �q4��3��0�}��!Q�S3�K/s�Q�L�Au^�tc���I��2��T�Ge�F���&�.e���j�+%����ɪ��T]ऀr5 �	��c�y��ιi-���Kb�Ѓ��Y�N�%�x�9����@)GC2�ڈ���*sr"u�w�ϟ����:����l���Q\L�V�[�^�c�Q�ꂲ�M�K�p�_�����G��a���?!�Zߠ�IP�t@����/�}+B�1om0HIF�k�7�E�a�yif�=Y�惤r��� ,�`Ƥ�=<��̂��À[Ki���=�	��`��(Ȋ�ׇP'�o��B��#�έzg���$\uv6�:��&�Tl�R��-�Y"L�����$E��	�"fZ���J,���&����{Ć���!����aD�4��6��ō�������.�i��}�>��{�V'����DFl�)�� MPo��b%Q���M��o��r�k��0I.h���ɫR�����dr�VH�P���9L!KiZ|&��5��m�a	9�}SCMI���K����XÁ��ɓ�1���/V�d�~|B����u)�^��9~���Pl!��r�ל3�"���2öߥ�����g9y�UJV޲����[OY&��ΆĐa3@�=Q-_�ڵx �T�.w!J	�N�d��J�D�4�诣$胠��2F6�Wˈ؁�����R����u�����St��鏶0$��5����h����Z\�4���55�l�tE8J�w�p7��g�[#-����F���<+���Y��~ۚ�Κ���