��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P��v�"<ߞ��&'��k%P碶�R�ӣ�sĞ������FY&v*9�ho�R�Cr��?�LL��Ԝ�t'�P�����}9�*�H@V�h��rŀ��Q(K �������vcn��}l�a�.����ݴ���4��_n]�N�s�øbJ/d1]����潯� �v�����V.����(]h�+ޞ�"�,ܹ�ɱ��S0�&E��E����Z{��P|�_-=u�t�9�Hy`�q�I8��gP��������i�����m
jї;���پQ[����Jb�:��!�)�M��H�쒭�TK$��ߟ�r�-I��0�u�Al�>�����&{��o�%(|�r�V�"��ܽ�[��jb����>ҭҒ��Yic�o)����O����̛�!Ԭ{�X�u��;��`~�
�%<���/r!���ҜE��.�Ԋ��^Y���LUB#$��|d@���RӇ��A>�����w����_�X��Bt�u[���p�M?�U��?P�̝���y��(�wA����<!f��w��.��_��3n%���u;�@��m�J�1�2J�8�A��%���.Ƕ�|p���tR��śh]�R*���\�$.0�I*���~�ݿ�<��f�H�Z��u�\l̋Wc�`Wz�:^�K0B1FO����	
Ү+��W���zO��}d�Qa��� C����TT/B�V�MJ,��W	=iT����ʑ=� =cǪ�Sx���8�N����e�LMZ�������=��Í>Y���%7"k���4&ap.��*�E�y�C���������`PM4�yӻ#�?���/1�	3��:}{��r��, '^-s�Vض�D��G��Y)a.Tb�p���.Q�Y�.�:Χ&���^�ğ�;(���$]���' �5� ¯�TZhJ.yv4NG�q�,���'#��))Z��u�}Úh�l���6���+\�ɯ�<W�G@�M�)�e�l��-����Q��˵$���ń����W0"T��M��i;��`�UG@d���Lkx�K����H�n�</�%���[9�^T�uҥ��\�ۉ��
ӌԛ'	��x� ����t��'ϲ�}�O|�=w\p�mI*u�Y��[�/����� ��U�a[���h�SvR�EIwDz%
{?�rP]jO cmXd�b��C"-�SU*~��i���5m ���C3?�)
�ȳ	S@����S��-L��&��S��T��g�D�@&�*�we�^R��<2�VP�H�6�K��J����A��f���J��{~��L
�t<�>{�&�)�%v��� ��7G�?�5�2�$�Q9nX��~yL�W˯!��ړ�H��W�Ņ�ڗ��WХVW��\Ɩ(/�m���ѯf�b ���F�CH�u�?�j2�Z�����A��n���)Q�U:*[DG�-�d��*��	��&�O4�%�u����{Y;ɢ�Y�V���S~��o��Pc��R/��fLL*]�EnRV�� ��3���`z��`���ɖ!&z0�� �Ay^Me�V��9�fF��.١&�ǧl.6:6�U�-Itsy��וR5��n�@� ᓏ0���CoaM�Y�4���9 P_�n-lַ��bY�5�)\T�K#|댥�h�3I��6��Y�H��J�FQU������6�͍4l��b�wfQ��C1/-kW�XMބ[#�
��:���Wz44�����"�0����r��#�i(I���y���JI�1r������;qA	�'9x"����M���G��3�A<�����8{��,
� #�s�K�T� �LңS*�?) z���r&b^��� e���h����+q����g;v��"�;���-4����gMKG��ǥn6;+:̯o@x��H�9����>1�����;�M��Q1��8xqe�XO ���	�P>+%�꒝NΉw�G��*S�X�t��Q������(�&pW�8���/=B�jl�ؚ�K�<\Y�(��׆g����[(_�ܣ_�d�I}���%��=DD~��Q�&���{���	"����Mt��R���C�UU�a�Y�Z�1D3�mR~/�U,y�l^��sl{��C����T��_v����O�'�u�5?�����Tk��Uvy��C���啔!�T� s�U7}����!@r<�����~�6�0e�,+	0wHDؑ�c���:X� �h4 ���q�1�����0&F�x������յ(?#��1�� /�S�W��R`�(��".�he0L�[W��Ne�6�t���4�3�s~M`ݻ$�7��$��7* ɑ�M��S,ߩ�y�me)y�Y]"'NE�-� }B�Fj�2��wўʡ�2zbR)��6��16� ��4q���)7�YY"��#Y���!��?������z���&i%d4����K/������(8�A5[_��Cw� �Wal��$qTC��=�#��p�K|ۚ���>�=1)�ύ�
R'�N� ?Iw�n�ޖ~� K��]K�8:�mw�ٹY��1BzJ�t�/��V���E��.��r�6yKw1:ܴBN�5�֧��e���˲ d��~ �@#��} T�˟�;�I�%�#�C���T�k��͌���f�4��ғkv���m��uV�:X.di�m��"FI��_O/SmJ�Ɓ�#�y>
F��^� �i�wI�~�d<�:pj>���	��^���I^���>���1C&r��h��v�6��۝V�r�(��"��9@/jN�l!KU���K����������>���{�$�c�R6F��H�K�֫�4�k��g�,��冱nl̝d	:N�Z�#�����k�����@����]�ȥN4U�%�%;%Xq���A�zq ��Qq�!�|�CU^[j�KT*[v�%,��֡c�&��ʢ�x�;
�}�d���_U';����jW� j��}%�>Pj|�1�w*�`<�rr�`jq{0}y��Ϳ}m�����p'�]�����v�5n�'����N�̸E$5���BC�"7���NFM�/W���j�Jg��V��J�+&��	*��jD�1K�Ȯ�����,z�PC4�jѲ�B��Iw>�q�9Y`dq�$��BҹFNl�<=m�rw}%ɟE��[��Z5Q׀��n���=�UXb�SG �<�}�yt`tu8��B�iy���i�����O��M�bL����`6�q2u���&��x��%&ls+�/$���w��(d��3]�W/`H9y�b��a�y)S��6���j��@	+��E�coᛃη#H�6y��`�ᶘ�+��t��r�7�x3}�<�.���0�z��;��f��T����z��8Pc:���_�.ۆk�=f`)t����g��O2����r�q��S�:V���n>�MWi1����~'���3�&�n���N����F�<���/�<�eՏq1�u-�.ܲ�x�9����[��W�:�҂1���2_�9QVޓ��<q�;@�K��:�5n�s����}E.8/ ��e�C�ƴ�[&=s�T��k�8~�w�	�N�r���NE7�9[�*�Fq=��h{8�J�X��R�5��������}��L�ī�X<�l��jm&T�u+�[Z#{��?�]Obzu������G���WX�|Y` ۭM��[S�>6��Cs飳��]��tO9�pK���(�֒���'t��|�}��ɘ�h��La]u_�0��[��
آ:0O��X���l�b���2�w��j��4���ܹ�����/s!���p���%1;�cZ�����խ�Q�������%�Dș%ˤm����?�gV^���|�I��~^e)'\�����gVۍn�(�
H�yԛp|��J��a�H��!�.��*4���&Z	�y`W���;��;@�u�V��s��f�Bv�V�T��k�А�!��	�pr��kB'V;Tm�?z<{�W}
�*��gmP��&�򺕀��L0�*㇓��I�x������m��W�dKJ���H����S�Q�k�Zn͉I$;�	v��Δ�b���A�u@W����F�4d�C��y�z�#�&A}��#ҡ1�S�������ODG�IŨdR_bKM��NuS�|�4�WCm#��p�e�k?d��%�n�\�OW��0�ɿ<��3�o�ʟ�Eu/��NtTg��ԍ�ۮ�SJ�ըH��K��u���H�[�388���$�q�@���A?^G����Q�0�����+�;�NHO  ]y[vD�?��zO�����B����pX\P��;^�Қ����!�+��s��@�2����fg�8