��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P��v�"<ߞ��&'��k%P碶�R�ӣ�sĞ������FY&S�b�Q������j�-v��U0�ĎP�F�_*��8��(�GMq�~(K�PH�A���։|5�X1�I �9)�9Z�OM`���c$<Y�8%��$�U	� #���h�:p6S�����A�G�1�K]疣ڶi<���?V�ʈ�4�,j9|KU��i�K6��C<�����9����^Ed8�[j �)KB/[/-�}��<�C�ڸ�y�9b���wE��%w|}Ùf��m�s����Fuv���L,�jM����37f��S'T& �5�3~"ha�S���
����c�+�t��m�q;*U�(��N
'2/;]#�4I֒'9����CIW�2���g��f�f���ʝ'+��%����w�;��iX��^>K�Uɚ�n��(��4�#����F�#���-$�Rs��7�1C$eʯ��EXn�����'�x�yX�'@����_9I�q�P�������p.���\��wV�3>�
=bd௴*�	��f6mD����p�D�	�{���uˌLiH& B�-�/�b��0#��0s'جV+�t��v200KT6w��I}�r<K�	"0O��Pg$�r�&�g����Fs"��j��(���(�SO�կ�r��v���O�"� ����&y�s6^bהJyM����z�n��O��c���#�,�7) ����^���T1����PěG�4�@L+.>f�|���H�No�o*b�<]\��jN���5�Zg3�Ǵ!���\K�Ҩ{�e3�bVJ Ȣ�P��wY��fUJ/P��O��M!��~��Y�>�D��#��"�>��d���ѳ�u^��df��^�d:��9s��0��,��	�;������?uxƱL�eƬ|�Y��Ic�����^��G]&iCVZ�X�"H���¿I�vD�k
``���_�S�:^��,^ݍ������s�ᇞ7JY��5�dXtz�V+v�5ΕCH�KPZ����w5��^�HE8	�9d�n��SU���`3��#!��/W�bxTǾ?O-T��'7D�J�A>�Ȁ�(������v��5V��tZ� �/�}c�_�?*��J�k�]�F�=F7��(3�&��_��ߓL�B]��� 2ek�<Q�2#�fn�9f�Iҳ���s""�;�^�����U��I�~�|f�Þk�'���c�vśpX��5�L|���(��ט��K��{��߀N�_�%>^��Y�CSy�����\���Ɛ������<7x�uI[��9�ʻ���\��/�nq��W)�� /���{t`�_�ɯ9m������v�K8����D���{�{�0�;��d��Z�jណH�b	���/��WVM/��`��.�5Q��3!� �Z���,7���u�����
4�bz4 J��"�S���a�Y ��wevU1�,Wj��/|�V��ވ#*����h�[:�T����h:p.0��z���L{���k�����:*������cӊ�X�KB�����3J��,��Owʵ
�@����A�ɽ�5�������Lu�x�m�%�\C�^���OHߟ�I�Fs