��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P��v�"<ߞ��&'��k%P碶�R�ӣ�sĞ������FY&Qw	��PpD���h�D����^Ry��
Д�$Ws(���;������!�W�V����������v-Trݴ_,�^��R��j���q�����M����T��+FlT|����lj�oLh7�J�uD}z�@Z<�;.MK7|�`�/z��@�z����q�D���f�N��u3��u䀝��#]D�̱�l@��]�i?��4�N�����e�2���Z*�����D��v90.#�/�'7�J��9�h����ثY�Ӭ{����@�\���R�jd�&��w�qI���L?�����;E���;��㍆φ�Qv��8����˨͍��(��������)K���UӽZ���Jw���w6D�·�=ӡ�xq��X�ᾁ���$����'��Tu�d9�撀&|�]�0�~Hɋk���������&#��^������p� �9��Ss�s�O~"�o�׳��MX�N15���B'��~F�{]���[[�6cm�+���m���������G�aω�l�
=������3p(o8���?�N�������J�:�єQ`�v�O��y�����*چ�"�\�Sz� �Lj�ncm��Z* �>�V��rK8�#&�01��]������u�3`�/�BX��e��$#q�8�*�4/����V�����6VfF+Y�F��(�^꓄�r r9�w�5����9�d���fN��Q��}2N�Ļhx)���`	����#
�F%���幏tj�7ǰ*�G�v$Ë�<e��Y,�Z��1b�~N���#Bܶ��"1TF��Il�FC��r����2�0҃���#ad}s�<@r ��A}�����"g�������=c>��`���}�А���X��%�����gnJ�r�9�x<�v�IԖ��v��K]_;S�d4���߰j���g��1��U��q�V�'i�T=r�IfJk��!��r�l@/*���~�z�h]�����BWB���EJ�Ty�g(�D�-�м9;���A�x�
G+m�oD �{��������;�~���>��d�r�-i~��e�YX�(:ь���nE.�����^Kn!X�[��br��jO��k��q,�s�t��vz���^h �b�ڶ ��~�u+���9�����dy2~-�bV��:���m�)h�eL�hlT��!��xG��_]OR5w3sK��ha��n������0ӹ4_rK�y��XOl��t���%���B�ad�[���fGU-v�℁Qc�{��,W��[}����dlB�os?�ƥJ�y`m�R�����+��������ȵ݊���}�~BJe����8�Pi���n!�X$���̞���y�nd*��m��p�^'�� �g'����ͮc�*❝��/�ɂ9�#��~��:|�߆�è�n�VؔG�¸��͹s2)��D�VW�u->��l�F|�t���NEU�[p�	�w���[�����q���9_�K��2��"�u�{���V�%�m&�x�O�H5�O{$?��̽�h�`@�^�w��S����o��HEE�.J�鏜D�Fp�)���.�9�ͽ6o�s񚂪Y9!�SJ=�[�+�w&$���Vw�@�.v���{�ǧ,)|e��ǋC\&�@C��-�!�
H��S�[�,q�)��������*�ur4$V���ݎ6Q�n�����B�X;ޣl�4���}qA��&ޓ�pC�_��mQy��Z�YUQ���!+q�s1��f�*|�~�D������->!�O��S��I[j\��F��A�rS\a�ļuh�Y��襜פv"Eh�(?ELv��_5f��j`���Z��6��7^��{]�bH,B��.:�����gd��!@7��m�]����c��q��^㩠���l��%c36���cƏ��������@��Y+rH�{q�=���Ёq8�������k�::�K�	��ERf�o��(���~m<x���kf�=\���D׌�rI�_��o�˃1��Տ�X^��F�3��5����od��{����y'f�X_2����W�����=C�L���8ъ��U���O6��vh���G �]�N3�1=��u�("��~�:� c�o5Q��7jf��#��mk����zw7����#E6k�J9 n8�ndeuyk݊2#�놰�e�5�!0��9>�B��:�i�xi�.Hd~�T�|-��42k�b��~��l���"`���/+�������A��+��-�bY�*ReAA<���l������k��&<������cs����	��܈w�Xj�Vm9�>8����%��dJa��������+g����
t��~�9�wg,�#c�Z)��	f����v]�~���G'o�#�# ydh�7�O%y�����_L([Ɖu�۫\��5&�������Fc�Xʾ*�S�0$�&�!�C�����!ޏJ�}$��ŉ��<��g-~�'�E�㠪��51s=�=(���O����rNj��;�/2F�]Bx��P�fep��i_�#��n��{.5n\S$Ff�s���!�o�ߖ��۟�U����l E~?�N��ޯ	e�h>�`/�$��j�mt%D*�n�/_A>F,��oZ`�o��` �yl�uNټ�9��~�zx�6�=�Qc@��I?�b_`�0�)�]�9���r�YX<ME��ŷ*P��Me�k�0͕�#��m��Ȕ��E2^�%�V�ՠ[l}e^��jWz�k3H��/fS���o2���+ŷ�$�)�C�
't� ".K��L��ΤF���3YR�g��o�1���)o�"B�*�蛹D����h�#�ލ�l��P�7Y��#�����bG��i�tZM���y���%_������95=P_��42�?��Vn<��������m*���&(�����&^�B�+�ʄg�Xyra��*s�k�:櫝Y��?\{WT�l���
<�F�ze�<����@�-ډ����M�P����(H�7�{�Oa��}|Ga��?��EX�ׅt�����Մ�q��s��|yvc'ӱ�(��Q+qm>�Ś��ꔯg�A�%��5�H�;�w���W�&��و��g٫�P�>�����E��p߆A$�/�+���?��E��{"J+*���Z~�n�%�р�k����S1��ah�ҕ���
9�v���;Ymi>�s���3�Ѽ��*d��w��K����yp'��l��/�>����N%A�+8ǌ��h�W�Ycj4��qt����`��B�w��o�\a�SN
vO��b��0���/��wUϫ�+��&(2�L��3xnf���ԓ�5������_ �=k��j�~۟ ��(Gc�+�v�*�RM{�я�f�0��o�~& '�T.m����U�m�_��Ρy6P����pcb��H"f��s��X�&�I��F
�{�0���OM2]��eKZ�����/M���p�1n��`?s�Y��3��o,; (g���Mdq�~�yJE��T����ş�-+Ǵ	D:�X��|�]��-��.&�%"����E{ws�0�	3���H�Fs5����x�j�p�Tk���Ƒ�X�9���e�*ט��r��b�q�,4��롭kqy��X�\���<#�Wk�O��\����H��f���x��s��ݔ.���x�ꎃ�m�Z�i1�170�,�+lΏ��x��{�5}��UT%������Қ˯JxLk�� �J�O8�_�x闔$�򩠢EN@0�$>9IK�`�Ps���HZ��Nw�fhr;M�ݤ�ZtAyt\[u�j`E5���np�zb��>��kɩ�nh-3u�ѭ���
�]�Ъ+�FJ��-���3�Px��K�O'9��R1����Rz��y����{[,�t��~��s��:(�=A�*PgI����Y�e�����7O�Ϙܝnq
PY�4�P��6!hAQǔ��1י`��t�1����O�oz7��\���p:�bwB־�-��z`��LC���m�Ig3�Q6
A�ڱ���b��E�џ�7I�Ozʬ���G���=%b��vwt���iqXS����1h������Wp���?G�q���X���*ƆLPr�����nR�cX(
7!�.���at9�����hj-yr
R���j���@kp���~6�zR���+�z���u^���&X4]g��R�bXP����5X�]*s�c�]���o���������=Lb��3*�~�\�u���t<�;w��[!�/D�7�-,_Q{	�[�ŭ��9�)Ö2�y� T��\�j�����ʅԃ�"Rw3n�TH������u_���b>d��E=Vg��_{��&m�L�qJ�0pQ+��#��P�A���9�	%z�G�� *���vW/��vs�d���/��;�θ@M :o�K,��O]��E�o������sЂ舶���2(��SMx�q��Ļ�6�pm��fz�~�b��C@��b�s�`��v;�9-7���e�s�V��ѬW�{�&�MȺ|�fp�kj�e!3�Xd�^\y���ů�������^Ll��C���}a`�)ǲ�v��x+�V�0:�k�^���B*H�9^�Θ���.��`)$���`��D~��P�by���������O
"� �ιqH�_`�9`���iԁF/H�>�!~%u���������xFFo����,�xB<�2�����oY� W�j(��:dVe���.=��O[]���}8>y_�#�����Z��C��: k�R���R�b ���UH��S���z���c��V���w����i��Y�Hp[�ٮ�뫌`�kB��Fr{,�*@5�*��w�7A)�WNliY�:��Τ"g�N�#R����:\����| e��$
,���~J���)����.�e�޾/�^Wژ�Gue:i�pX4��H�>%�����Qs�ڦd��+�]���-=�-����y��?o6i��%�#����p�F"ㅚ\�K~L�G�\4��	{�1��@��'U�ͻ(�DHQio6����(8��n���Y�&�����t�R���e�ZS(7;�PE؜��AT�)��N���U��A�E���7�8�~��d���݋�߸�6}{�g��3�|_&dKP�������V{E�zTq�#�x��,�e`˳R�%��\�v����ѢF�CG�?Ƽ���
Жݐy�]�Q��n�d��:"X^�g�4�
n�?�I�����`Z���j��e�m� \v�x�C-�d~5���KON��Y�.�.0B��g��yr��k*%��W/6Y�3K�Vpxŧ8b��+�i�`�Ƀ=�����4'��*����?q��B�HΒ��Q`��<��Oݬ$H݅�!䳃�ibD=�ڹ�!�DDVY/�Dȯ?w���l��/Xge�Vfm����(�F���O޴��:58j��ڮބJ�=Xx[�I�@vIll�l:���Bր��Ȁ���q����'�%
8c�Oy�}���L}+?��=F�
g�U�mک��9~�iB�:�(oh1hV
��=���4�uRG�۾n@>�P�06i��pT������\��ݯ��ЇE���?�G�1*� F�p���ۢ�j��_��8ie�m��Y���*���)sw@~��x�p"�,�v/'8v�ܣ��#h�ʏ���6m\����?���\���+#�]�4�/k��F��s΅�jߤ�[^<��jh�r�q�Z�w��;!0�߾�H�nw��N� s�>#�Ef���wk$�c�8*����|69�5q��f���,&߰;/�(�|�vݟ��y��+ޔ����.�v��pW�Ķv뚡K�%y�P?_;��he����*|�?gX�6��	r@)���@-�ÞP,jH{E�����#���B%Ն�P �(�겛kr#���"Ir�l�LK=$���T�CU�?��~SG�_D�5Y�|�31�|�<�1����B��a���`ѽ�l�����sK��N�ʽ��e���/^3iҧ��F:��`L�
�Xit��uur�����'�������C�;>��QQٳ���C�L��{�Ok@x��lP��Q���B���Z(X��K�g*�HN��L% U���WF��� T�mòG8j���Q�.7��>�o��m}"H|𨰏zD�+}�R�ٺy�&'���!7���ٮ�˛��'� ��v\���ł���#߁��c^�Q|�@�&{��e��@���,49՛��ؾ���v6t�"����*��S�Z�XK�k��\��[�2�q�7���r\:UV��P^� ��L���6Z���4%Z߈M�n�R����L.^��7�m���6�O>�#(PZ)�w�ߥ+	|�
E*��a�D��j��?n��߭�Acw����)������u7�m_�X�����e@����u�,�e��->��7�7�Eo�f�Ȑ	�Fn�~��2n�i*<�,�F��fZ�G>�Kd�v��+x�ɂ ���%AYtZUN��nB������S�ua��q�Z��~q�h}/�55�P�!�c�v���ѫ�1����@�"lp o?�(�X2� o܄��]u|~�r�醀U�ZHSlZ���Ru�5qRث����O����_���%r�I |GL�5����q����{��;�P[���'C3~'Y�s�).5��`'!�P���Nzn�H�1��'�D0�ǜ�t��fP2�ސ�����Y�:rD3*�p�s�5Y=���&~��?��c%�X��r� Q跼y�s�84l�[�%O��3�/�/���ЛW�[s��/�b�tU_�1l��������O�UPf%��D�4!u3`Q���e�]�z�,�К���lT	�P'�g��'�ע����X�,�Wˤ�+�$wA��SpȻ�1���@��%���i-ɬ C�������mv��
-�����6K�x���0�Ӏu�|�f!�M�nQ,�?�}*��~�F��� �xH����c��<Ź�P0�_� !�&�B����;$
n拸H� IƯى��/i���S�4�dȲ>�@
��[���݃� ��:�؅����؎�FDD�o�6�ٽ���n����N]��d�,�H��wV$3+���p*�0\ו�`ZV�t[�dɂ/-=�;��u�Lߗ���z0y���'��c�b��������_���iC��-�`����h�w4�nK��d`B���u� 	���PIx��/�SbNW@w��%�x���+�.H�p�Þ�G�q4_�������u�\*12�5ؚT��)M�L��ɷ�^���\��bl�!���6�	���ֵ�7[���\��P@Mø�sD3�JʜP��D���B7��2[aB�$V	7� `]�l�T#"m�����{� �(c����V��j#Oq���$��#8�ѲO$O��oa�9�Al�0q�0��^������R1��)�cd�5*��7f�@c�6�ʞ	��o)׶�62`]�{�0��γ�6y�����9B$K2�i��^b�G�{2a6-�@�'ͺ�V��/�b���æ$v�لǨB�N~���<�sr'��*�<��)\]�{�}E�x��`�%��M��V�B3�nT�����v��"�	�-�A����a�A���r��_&9��bp�J�ߚg�Ke[�|��S�ZA�`$���P��\^�h������Vٌ�����,"��N��Q��K�ۙ���^F���>W���<(��˭�ܶ%��Wl�Y�R�k���-��������t
z����tƖZ����9��G��/�-�V��Iʌ�;�D�E������A�Qƻ+:�ިʇ�k��6����ao0�j�G��B3p����ڛ�����,;L��D��gY\�D5#�'%����|��'b j�p�@9��'[�'.Y�)��}^#'���T_[i�ĦX�ߟ7��$C7��6�e���˨�Ku�[&�o�P2��qT��^A� �x�Fo~�cF���V,⪡g�?О_��9/�k�ꎁ�.]z0�GL�z��w���q��05{�y%J^�d��ۀ�1j#��1�A>�y釫���$+����)��H�&fJc�W֠	(�U��D$T9����`9��R�o��Mθ;��7��,�7�	���;�T��"�Dھ�:��%Ҝ������m�M���&���	�IvI��h���c����*U �N<*�{�A2zW)��#��LŞ-�.� ��B}�@|f'�8r0�7��ko�7 �R(󣔤�~�	�CJ���a��Yl�)8�RD��� �Y.��x�lK������B8r��:l�\���u�����U��K���YRĢ�
�55�F�VVP:G:8�Ms7��"V*ۯ�˖Xh�G�I'�GBm�^$Q{��3�7@��py���n����X5˖_����~愉����6?�eL�Ջ�a'G�[0���oh1������G%��(d��F�}��RrB�O����[�s����@��f[2�*������f�Y��CU�x;;w5�vvW���T������zi�꩹
ϛ�OI�5��y�se8n:ɜ>8X|C�Y�ќ�l�	��oF�1@��R9�0���V}v� $0�&q1ъa"�蝧�>�	����ќ��6W�����Y�C_��sp�;,� �.����e�x���V�$�����y�t*�4���Y��c�ј�Q u��E��U��k�#󼐉4�4re�*���lV357��ĖUy���Yw�4�u�mG��1����SpM�Cn�!�8�H5y��0��?��"���,9��!%B&���b35
�J%��9M�_�:���敷�Og��`g@*�������>EF�'���q���0$�y17�tN����<��ECbs�G��dJHe�
�VA�&Q�J�|g;o�����U��M��,���sq�+���%�ĵW���
 Ebz�VyP����f�+�acQ�8v+�i��@��g�>�\?{��^4
�Q�&fg��n��C$&�^s��ܸ��v�-�nt*4}����h������\i4
v�;��/�p9ʩ�W)�gEn�z�v��>E��v���a<�z�@}�S?�d�h��ٍ����Α#��;>�Z�\�,:@W�=䑚9���!�����B��B��U_�7�0��{P?��oR��	fI�[S�Þ0�P���C��i���$22%�H��`g�� �7�|���� ��I�VQ�uڎM��v����� �Dy�*,��/X!�9�g�3�	&�J��l���W�Gl�]%۲7�내��n�!֊b�X/j���c^�|��~��t��N��WA_=z�ۭ%��v"C��s��qE��ܹā�N���L��
B�p�jɰ:29/�z�,PT�d��S��g=����,�Z�7����;8gQ�](ֆ�%�U ��k�ƥ�ӂ@��$)	H��܎��h�b�3���ӛ���]�19ʰ"�����E�n��X��[����mȌ�O�:c�I��r��Mj�������ꉨ�ʻ��z{B�L�)7Nj�󖨨��c���[�x��[�?
�Գ8�N�eX�����(&�2U�Z}#��S�5@�Q뛪�o�owP=�A�6��j��}�T�&�"�i(ڧ.J(����Pٍ	�i��K@��Ān�	^����?j\q:�b�Rs���s�˘'v�$��*�樑W�A�N�`V�Bi¦N`� 7�U-�)�������%A����J�ʎh��ò�Op����s�X`�"^�<�?� ��Kn�z�[��[�R�V��|%�1�Iڛ�S�c2�1��ʒ&�f�`�������-и�٫�a(�q��U���}	 Ɛ�i� (�-y��x@@��j�G|h�4��!��ɱ�}c���d�T��ABS�Tۡ+[fܽ�̐c�C�����uRҼʂ�y�c�Y��k�����RUX^;Wl?3�����b���T�&�zȽ�)����`)R�����H�����P9g���S'[�7��5G�����?�=ku9Y5^�@ؠ����M9l��5{
P� ����:���gVh���~uCA�	x��F�@����J!�Lnb����lu	%����������b�N��L-t`%� ��[(�]�}+�v6C(r2)4�|D?�+������d�Ex��&S�U����T��lg~E��G��5YN�!7J�@�M-���+v����z�_/$�Ja�B/�5`���;���n��z[M�@�"��m�ONP3VeHm�Yk���9%����p/rf7���"��dxb�u�k^��u\^�N?���������x�s��-m���Ng�Wױ�q��<g z( ZvU�`�6E��xH��d��3=�^�F-X�CP+����W�eg�m��툚�����[9�n7�a8��a������ӫN&Nf��[��.�