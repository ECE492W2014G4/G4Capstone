��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,��.��̡�+P�FuX��d-��N��$%�I߽7>wN����u�]��j��ܹ�Ucל�|�=í[~��k�5�P�ؐ��T�5�����#�p"&�l�z�Fr&b6��,���Fԟx�ɅT2n�x��p����Xh	H���9�Ҿ�z�1�� dT�h6��[I�����B�?Oq�_2�9Ӑ@�p���G:26�[�6T%,&'�#JeR�+񸊎2�Դ��E�Jc�������5N�{�����Jz����+�:��G˦�<�_�	�'��k�Ov-��5l��|~+��,�Z��r(?�! WD_����J���K���םcE4��%2���qb�B^���p�G�A�tx��,��66KEك#")����,�y�I�2�$r<f�a�\)��?<��r� m
_�
|�P��i�����	������9��4��uRˁ���1�{~Kr�	eM�.O��+�e����Pņ�мfƶ'H(Y'�;���V��j%W�i��}��b������D�g ���(�����4d��"zf����[��B����^�ގ�L ���R�}����W8N��˟Q�v����R�w^UO�à7ZW����2�j*{m)������ ��Y!��+>q�*kf6�C`[w�IB,[���U/��W�%��h����J���|����U�z���Kc0*,�Z;��WM�2�+�v�]3��h�r��ף��gk�����-m),���2v݄�i#8
�_B�w|M�A�{���I.TF,�NR\z9׼�[�����t�@�Q���~n�^6��qfV�y�q�ǓO���F��dM?x՝&㒎�q7n��s 9�d�i��+a��*5�z��a�]>�6`�w��}�D��U2,CB��3��]M?�D�D	X�7^����dǞevԟ.D��mɅw�K�K ������G�}3 �c��L������W�6�i C�:�߇��ȖMҸu����@]�r��b]�<�W�p=i�R�H���v�$�lmy^�h�$��]�S�ݕ#C9��[+?`u�RVTc��n��;�٠�"�~�%O�lк�E��S:΅��v<��:t�a�����ﶏ��I��6�M���-��Ç�ysu�!l�����N6�=ҵzx4*��}�7k{P��n"��qw-�(��l4a�p��H���em�30C�v���m������mD���f�i��GQ1s@rt��k�n���:��-&B�D�=���#~�;ۈ���4��hi����B�/˗�w�iЙ$:R�V�g*r�~�����UNf*��2;��P9�`\�E���!�a�b��X8h���{]�6��F�%}�H*_AbS�p8)Ԑ��ۉ;j�yx˧0�6�@b�PTL��ZW�l驐Ώ��v����_���n���5vp�A������K����򼉾�`xdP��!�	iWֶ�::$�ڑ����"�T�0�8�8e�ߍٿ��޶���^�T���A��3>9�V����|��B�@��:�H��y�R��V��[��N6sg?�k[2\�)�7��DD+�ڍz:$���ͧ+ΎLl��_�_ݎ~�W{�g�iv풞�M����%O��8I]n<�Wk�ju���M1�� FJ��\h���$͟�bMNɣ��}�v ���@�k��6f���޻�E�
p%�-i펮��`���^�Q%�
"�Iɰ$.PpoCI<^��*��s�W&���`!��K�Tt����Q�Tw���u��r9�@'ᢃ��v��y`��[ 1s�媜�b߸(�����2���u=��֊SK92[]{iH�uN�����g^������<���X*��(�����3͝��������o��VȤ,��������8oQ<�PC�ql�/:�4�D��S�X2|�c|����W���f�ryù͟�Pw�hv��b	I��(M���2xEp���8��\V����1�4�7']e^�?���?����(~�
�hH<�欛�m$p�b�@O�i����+1͐Q(�:�	����=�s��W��{IVL���������J�5�f�Bۙ�|1�_<�z�,�-[l���S�Y6�e6����Q�����
�=l����R#U9Y8mHHFp|��+2�De�NN!ذ�[,x� �-�7WZQ����
)���*Y4OA3ݭ�-e/p��=����Zɼ��!Ux֙_���O�('<hU�R��eDd�z�-5�뭟�Ag�V�<��oZy���1۬�H���я������ �FU�Q��4x�����|�ѸəX�~�h�ua�J��d~�N�^~�TQ9�F�3� 
Ĕ#��e�B@Bֆ�CQ��(���I��N,�)��v�
��ǧ�:�1�����F2ѻM����/eZ��/��H�C��Sʁ�Hӟ��1�_�9�,�)v�F�/G�Ua�������!�߸h{����
vp�:y�a�zD�_XV?5�L)�