��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P��v�"<ߞ��&'��k%P碶�R�ӣ�sĞ������FY&�zH���۔��RaǴ�{�˵�j�u�6��� ��',d�	T3�˔�a�S^4Jn�����F3~�7��4l6�mq�A:G��^�axD�i�R;��$�y�rǽ�%�1���ssu�*Aŉ�;�O��P�s����ѿ.�M^�mO��%ϐ���8��_Q�����E��1X;$���J��%-�����
��$Q��l
�F@U�k�7ˣf�da��n0]F��d��9�x̘Z��G�N�}Bb�����aw8�*�ҭ�L��-�.}�I�� A����GOmNш3EQ��;�q"ب�`��[��CN���
1�p���׽g���B�B��i�W<������JS�b�u���vr��|K���Ӣ�DRbl}��.L�s:�w,T]N}�[���0bu,�t$QM�T2;���o�g����!$�"�YJh$v�%I|��]���7�O��I�gds���ٯ�_5��>���rF���0sr�b�5`qw�|��&#�ؽ���.q�,��h���&0@xqB�W�w��b�$���_E���c��r{�����u�'�x�V�w��T4\K�{w�F|�8�U�������C�[I�e��}����D/A]���!���l@`-����2e�5��c<[S��	ɪ��w&X }�����9ӠsϼY�����R���A�aj_�?�핟��N!�ZZ��Kh�.��̨o����_��i/���f��z�&�T&� ��S
��c3�pY��N�L�D7�-�jk�(A�8Eg|B��?eu9�ZDg,R%6���d߆�YJ��N���)�3�� ����|ʫ��y����m�?�i/~+�?��)nS���J'����R-M�9d�qaSgE��FHf��5�>���/�pk���4=N)��[}�'9e/�^�6��Eܭ]�C�Fѿ���ĴH�-��j��=G�s���-dk����'�PQ�"�U�&dۺ0����HF�KC��.\ì��bk�(����Au���U9:x��wM�W��ҿIK�ozIWZP7g�@�*��C� ���i�r�f�ُ�_sہă�e)Z]��԰�Ÿ~$�>�0�ʩ,�u���˟���NS��͠����7p��e{�u�R�c�Y?.Ҿ)�{�Bc�b�˶b�:ߟ?��l���,�]�qRͪ���A�	ID��i.�֞�L�p�я���<z��ʙڄ��\Zt8A���N��.)�=M��rބʈ���a��m���w��}���v���]�,0�-��/�	�W�C/ò���� !��T��2H���Gj�&؀͇T�ݖ#�����,D���:sH|�)FT4�hg���ɼPS>��x��O�?+�d�&] �ɺ�H�QuX6����`���J�W�&��z���g�m�i
;�SUFul��
��ia�S��XjX��;:m卝 	�^�|֩�O�
TQ\��_��e�js����+��_<�]���30��Su��KC��@~O�f6YgXė�M4���w�����M. A�����N�t8g�����UmpW�����s~���HLG}v��S�6�NDQ�?*ϊ�u)z�]	vDA <(im���` >k*�����,e��緼ņb���"��[�W0LY'[�>Gg�#O�v��ܽ�����MU�fd�MZ6�f&M_c*Q^L6f�P�$�Y�¡�l�SJ��K�"n�`wE8����VL�z������p�G�J�v�Թfg���>�����mu͔�����ϻ��ӏ(�/��F�<�(E`9���@ic���B��8��{�yCoP��`hU{>�-L9\�	��Փ)s]L���l�?��Aw���:��4�U\�����5Q�lԥR͠�@m3�Mm�7�4O�������h��+c)��8�#�K貏/�~��D��"�be��V�5ԁn� \�ܼq�,���S�
�zN�\Ͱ��(z��=�G�"��U;�a!����}�8��g�m��t�#
�ڋd�|JЃJ���p|��eL����yL�����&@1,<��X��F�D��Ï�����w`|u�s��ǒ2j¶�m��;"����s��&���֛����.���9m|V��xz~�+���N�LS�]I>i��L���O�9N�l�|��S�u�Ǿ��HOjiނ������Y�?����I��74��-�N�o��r�A�?��_!�K}k=�*jll=/H�xӵ|�wtՁ^D3�)���e X׆̺����J[*��?����o<�}6�N�����Aԁ�ӬK{B���x�v��X$�*��$N0|��^L:l��X*�%���V[�֎��I��n�J�4�b�?�u�i�h� �W7+���nKȘ������%�P���:�-�&8 "���e��d���Z)9����+�xU��/���Z�3[�����`�AD9V�7-y����v��k�F0hՎ����1�I�yY��6�i��}s��SoԐ�\/L���	��0m>�[�����o�z�M���`v�5�B�!@k�#�ZqӤ
F��A������ʬY�_���8��_���8snV���e �l|�
x��(-�pW��e�5��������X�	U��WE������p$E�%<jTp|�;�7 �T��K�Jdy�g�H��#�@%��<ڏ�+�@Ҋ<��8U���5��*�$�i
�����OS[�i����D��c1g�M6sy�[2�Ştm�A
+�B���bM����Q������Lí�����0�^\f��-^���lڸ6�T��c'V�%&���p4dH�i[L�V�rlt��ѧW�I3�`��޿���7�K
���q��6������V69���$EPw��;���DÏz�U��dqz�;� �����rX�m�W�Q�~�4�%$p)&�(+-�7/K�gI1��V}>���K�j�L��V�87�Ը6�����SǣT�0����(p����Ŋ�L��?E�& *�3�}d�>hU{ST; 9���^��Q2����Q3E?�v�,��P�;����Z���HV�<#{��?D�����qw��)�W,��	��q�?�,W�$}��T�E��E�2ϖ!���q+�c���e�}���T��ax��&�f�DϏR�k��[��ɔ-N@9��f���+�Rb�����F��O��?�k��]_���Ā0��r�Kr�]� 1���B�tY"���] i�ɏܜ�+a�g�&&�T��#��#��n�g�;�\^	n�ej�����i� �+�(f����)JٻF��!d��~?��N��Dǖ>]��"}A��Hj�]�7�9I
N��,֎`�y9��=&���X�Lu%����ŀ�
�S���P*ip�Ms�&I<ܒR>j��Zǃ�ݴ���ģ�@�a��Z_�_j���.
Tji��:U��,�w�\�vJT�R"�`�[�� �-� QQn� �U��x\)�/Q�Z�҉׬i	aF}�U£������J���
7v���+'A��s���\f�cW�x�7eƍ�%F<9a,GS>'�i]�~[��Z�S+D(v>P_K�*cյ�๨f!�M��8[��T"Gq|�n�Ո /�C8Wq��Y�]��i��-i�2r^�'0�v���J�ߛ�7��Ŗ2�_��E"Ϳ����!Ǯ󧘰�}�\�.�K��Y�.�u��ƭ�<[=k�?BO�Faz�f=k[Ӥ`���C��$M[��/��XW�/Mfm�3���
*�c�&ǟ>`u4ͧ7& �=�ė-������7�`9N�TД����ߦ��{��0z>b���#u��S�����X�Lv?s����{aŕ�*А��Jt�qn)l��)+�v�r�V�9ݜ결���Ѩ�_A��99�o�<F��)e��`n��{�����Iʡ��;��~o	��ִ�?61�`2�jn�t�=�"����g�����@bQ�����`$�G>��� ��7�3{��]�S�z�^4�`��$o�:�����1,�;%�*E����-(XҶ�(U RC����
(�x01%�0�z�/"�K���5�d�C%�!�)|
�K丬���~"�y��3��Y�_ຉ������bv"�Um�7���5
���ۨ�'�)#F^��2Z���4��i���%�R��k�v�l�*����w}�"1WRD�^�&56*r7AQ�h;̞����e��;�m"Vl��"��~����{�'㧢�[�ʇº>�R���7��E�� �	�c�a��'�m�FE����t��{��.�W$�����6��Xh����Lq����h��8�1���yl�'-�Хv@�����T�I)�v4��d�sh��g.�n��M<�����$�gs����e�d�c�y���f/Z�G��1��?��}�D�'�������J�����v���va�����҂%�}+�F!���������&�QJY��Y����1[L�~4�_'�"?Φ�A(y��XcOQ9C�/Y��7�l�M���v�<�5X
pXjs�5�8�:U�����ir�P��@��E�I�)�8����.`8�����
L3셩��KR��F�CzY�G�/�����xK;�3�FĢ|6�z3d�U`b��A@IִG�BL�ݑ(����q��a�� ��K�P:��%U�iH�s�@\�=_�O��*��v���W����ז�gl��R����C鞙��3��ۓ�8@��^"94�>k�������a���R�p�X;S���^ע���q���D|����Q#*���Bd�z���;���b�׋��u�U��e���V��q��8�с�=H��\g�W����<�>p��ׅ�:�4����c����F��|J��6�;zW��������Av���6j�@���p��UU�����Ś�GN� y4G�z���?5�Jq����/L���U�Q�{@{>}���H��@O�N��_Yן8�.�<�������t ����7�Jn��y�}AU0��K�%:�ψ0��Z>99b8f%�������R��{�4�z��T��b�_Ϟ\lek�$����)���%�F�Y_�S@8�B�=�������1y~��P��f2���]�*&�;D�(v,�nbb�V�=�
�d�4���,�����!����rS���C��#���,����G[��ӿ��p0��J�X>�hx��{r�B0!a�7/ɹj�b`�	�5J��ep��b�U��)�3�*A�N^���Ⱥc��5���1�r�u/��C90�L�2GAiy�K�$�3�E����f���"�y%��)�@(5%�8�[����^�<��&H�V��Szr��<i8W��]���-�� ��Ō{M7̉�e��nm�C���l5���j�%�[>։�r3��?��u�Y�� C�=r�2�q4�%]:��T��Og�m�x������ZP�J���OK?GWM��?#��"�b��`�`9� �c�n�>D�1!�u��9�i����̮i��ݍ�`�f�����Y�4�_���n~7���^�ʑW��H7���\�Y�b����-�J`��7�Q[�~L�,�]iZ�����?�?Cb@��u���%�V�Qp�;���!򏟩�k�&�8S���P���:g���ߨA��M��!WA�|b�Qk�U娺U�6���^8E��j��.�4�u��2f�i_䓊�կ�
�Y�Wk��D�/�5��HI0�)�G4��M"�vD�,n���	C�&�%�	��D#���6A��,��0�9���m��*�v?ň�O�y�6�D2�"3��b��=�bvH�d�ܙY� 
� ��]r3k�1�P��]��p�[��*�'֊�y�?�Id�q^��)B��)�M��;���i���p/��`�{��ڶ9���RY�f��р%������,܁s`|`��&o������nK��Q�Ō����O�j{�0�j�������K�*I!	���G��_:���ߍu?ߨ���Q���/`���F\~WJ�+I����7,�Z� ���,��|��o�O���hQ�SwM�VZN�	#�{����	8�t���Y�R'u	����:Pφ�R�!�{� .�/�D��sda.��4VAk��\}y��]g��M��_ѵ�^��qb%���gu���\�N�%
� O�}u��C�ߴ�jWb��^,��{=u#��x ��҆�������@�hh�o�����!�[�,��f-r��[���V̋q�ڤ^�FsU��l� ��~����ߕ���]�*�+�"��oz�2xQA��Mm� HrVL���[���esİq �F4�<``����P�����^S�5B�3�?~�zpCn7��%�^Ls�Vp&�w{J8��l�e(�K�p�C�znM�
Rk���=I�[d�7���йC�3l�(�I�y)ׄ�[������&oH4(�rH)�M$.��4qe@�uZ�o����y5��&H�T�p����1���~��?��?,HΖa|�/D���=�7�gdK{�0����5]Ja*�?B4A)���.��2Sd��d0$�m��)�1x���|��?fO�@�ߎ+�~�X�-�m���"&z�J����k���T��/Q9�b+O�o��-*�0�����*�3�m���^@�; ���t��m��#ͿW�Tt��z�J�+:��Z�;#��+�A��
<���=�5��ec�3��#-L�.��93v�!��f��P��I(��S�:]���d�֗#���gʽ�م��Q��}�ap2㘼3������ӕ!�"!,gsrڞ�X�:�p%�_�u����+���E�늖�'����r�Y>�����3��s\ES���$�c�Fa��~,8dGG����qeL�&3������?>$�XL�H��/X-�m|��i~��CC�u.��,gOY�d���~��<X�iد]��d�^7�5��.`��"��b_�]\��ךU2fhT1�饉9m5J[D��p�J<��%]�b!��~CRӔ���

��t�*XC���W�oM�۾��fA����Ú��	�zK��*E4�b6^���B8��e��?C�>�~�c�Qu��A#�R�&��Nw���>��5���<���.��B��3�X@�1|���]d֍DH��N�3��ɼC<ǥnW���jnRC�J�A$�kY	��_]/��{fj��c%V(Eǽ���<��;䡧ʥ<q@�y����#�meIm��]�P�u=�/�s�(/~i�Q���y�P�!�i�b0S���"��>��<���D�ȫBEٚV��h��ل۳��Q5�au� �~��*f6��jS�_n�@�gd>�d�^c����=��y����U���%��H��:|DB�>N�
��C�U�tK� ��\���7��x���D�mR���8u����@hƄl���
� -��]�ǥ|���lyq�0h����_t'ʹ��-k�syA�u}���o��{,��i/��d���wM
Br�?9ّt��z�����d�41i��q4�P�msC��/�+�xM�x�2���S%�_����?9�_l�Y��@h���'��%���H��Ɣgq�b�9�#ʀ�y��t]��_����� �U[Ù��!�S���e�.x%x
f�D�^$����WQA�fJ������g�R5��y������~|��%�&�3^���}?����^X�ݪ5���' cg����P�!I�-�L��1W-3���{d���2#�&3wۇ�۶ �ר`2_p��<�PXXai�c"%R��	�oĊ���UWoĿ�Q�jF������,��vf�߅o4�`������8�x�(������z|�i�����So�i����}L���9�(��0���/f�����eW���Ոk+���9��g�����m'�*"��1E ��T�g>A�l�r���X�LڍeH �F�B���S��Z���^����"ufߪ!S�Ɯ�k�:b\NWa��p�����=�"����5�Y���
�F�B�WUA�����q���e`AE�υ�ؕu�^������4}E�UH'�y�1�u�mZzT=�Cu�������;��?G渜��<��0^��w��>ɟxx��]dO��3�#�K�m{�@��~�����.�2��������2R~i�W�`k�Z��u�з�	C*Ғ�}@�����%i|��F @cc����&��P��W"f\��
�R���G���R�GE��"�1�s�^��ޟcu��W(fyޕ�ˁ�&�����=�n�\�z@"ݿ�5�E_�D�6�>,؎&:�<7��9�]����3d �$p���8�M���vJ/F]���{E{x��� �fj��լ�o>�P'M.��-�E����s�-�F��F���=�A�u6a�<[k+.5������e�4p��#@; p��(��70t�tL�Y5�7��R�������G!GAM�$��r����C+�� >�T:����Ҕ��W��m$=8?�1�����c`s�V���aֹ {2T�=�l|��v�f 6��!m��X2��dq ��ԁ�C��t<�k�v.A*�ucs�ɊB��b�V^$�s2��F�-�� ԫO�ʇ]9���Y��+�w�Φ΅������mt��{!xYg�o��w�fu��jC��4m���]���ڵ���9D2�~�i��$��9�Ֆ�
&'�rt������n0�S��<�|�BcT]�XH��]�Q�Ϝ2;GR����Qv5 �G��)����O��;Pʰ�J���Rf�jW�Ӽ�]�awd�n�MC�¨��H�ӡ���eFo�
���`Z
ޭ�$
52bQZ��F�&=��^�� ��>���3�\�Ģ�_��)��Y�~\�s�e�f��P�Z�/����L�/x�yZ�<�T2ݸE� C���g�o�^��W8���:�|ω�i���\�Ԙ��)��1|�i����b�m��D�E�����d��ƀ��H�}�;�$�(ª[~��,30BU������"�d�H�r\7��C�4������^�ƚ�g�t���91$%-b|��I���N�v�R�
7�G'*<D;Tcc�,�F�a[�����F	�1r+���p\���[�c�fU@�a�� =������Bn(V�~���Jyjfc�����`W��W��y�'�C2� �3�)a���e{	5�x����X&�o����Y��O��#����t�h>��ҫ�T��$u9�	�q��{F�C(�N�;F��y`P��5��}_�R��KWC(�'�O�UȐ9v7��wV]�$!��g;̢Q#%�]�������tJ=~y��MQw<��~����(���l�����խ��C_�//���ּ�"�>���O�@\���������	�_{b��Vm�ݱE�`��ps�YO�njcV3��Ő�܆s��Z���]H����,Q�!�1/#	m)�� C�wSf��[J@U���$2�̽�:O��9�u�F��b����mĞO�fџ�5���g���Y"*8��	Kyw\��m�|g!��<��{�r������օ�o���a�:��F]��;%6U���X,�����������	��-Q:�g�����e�bK�W�Y@�ڤ�tvG �/�oZ�p���ڢ���j�'����L���e��[߬��۪9��\G�L9��]�/���������	��?T��b��@C�2 �W��n�Ε�>t8�Yo���ǃ��c�u1c�YĒXEi�5�#�H�A6�`r��B��	/�El�[�D㼖����f�0d�ꦯ����:���6�԰G<��Y�6ɜ�W'��O�T�mp�{��_��a�
�s�C���O�i?�ټ�����ր�g�9���GKo1y��x�tk��Yw�:2����:{J8?�]�2~P1�X����i��KbC���V�׀]�� ��گS�V�k�Ax�� 0���|Rإ꒧�e����q�
�?=�5�"\���`�������C�] ��L�@|`��O3��9�U'�*���I�D@��8/��s
M�"��3(�؄f��fe2�l#AC�$��߶[t�T���&�[���I��-�>�Vվc�.�4˭0�;��+3��T��\B<�sɕ��+��tc8�3����F	!�p� [K���ga0�� a�o':y��!���q�[tV��54tO��J�?�qp] f������ܒ�jㆬ_���8	f��YH?�5]@�QJ��L�Z��jD��U�R�S��&�.���f��� �&���4"��,;�I�o���q7�8��ht���fc�L��V�;�� Q�ߞH��������q��,ı��+��L��:�����{<�Ɓ���{���$U8�q\hǅ���2��z�=QI*	��5	��8�Ȉ��`�Y_�H:�fqct�ܥ�;d���O�%��@��pp��@Ս��w!���2�`������_m��F���E[�`��W0IY2�e������2[��;�_.�կ4�����m�|JH�H���v�3L5��A���`G`����y�)��N���|�c���qXA�9�W���ԔT�C|í:reL̈�ܥ���-��y�i�tϘ�zN���P��(c�t ���˰,4������ߟPo��n��~�|0*�T�#г}$��4�P�p�H�C�~i��o�Q���̎1�d@���ٮ�D'Nsj6��֮���8G=-�/lp����فB�~����+V��dZ[���s!2�Q&[5�/��(�oD@a��XY��:6��8���3�J$�&t���Z��i�n�=�ޔ�j�����<���ÿ��hA�ArSJh������{S� 0����C[�5�������wE��U_g��)0���|O�zSw����$�.z ���Y�N�Rw�����U��P��]�'ӽǯ��v�� \�M�/Լ��A�L�6�2�4A�&���:�`^�?��C�#�'�#	�[f���z>��+��00�ܒ���?�+������8�c�_a���p���aΥ~<L�҆�8?�Vss��k���!L�!�=_�Ms��u�Yxr,l+8?�|�h�Q'݌���B�m�{�	�����mE��Mw"J�� /(B�-}�7�re���AE�57q=9����K��W�\?U�^Ɣ�;��� +��Ņ=�R�?Jx���l\i�Lc�i���Ե-��hv<n�t|��~M�OL��>���Wo��μNu!�i���S�%�����K6������|r�����P��hCd�Wq�˽�g�LNT�|��hL{`�IR��}cLM�_������o���U�;��63V+8=�@���X٢*��l��tC`��O�
$x�9��f-�#�l�+��z7�iҌwm��ށf���(�(i�|jW���u��̼�Ǥ��S���d�yABԨO�U�F��Ǆ XT��` Z#^�2d��g/~��x��9�Q�8c�Yⓖ��I�D���E�ٙ�17�4I���ř� �N)HRR ���4+������K�$CT2J�o����)�3���
����K��R��Bt���3ʶ�0�B� �I��6Ev3��-�H����9�/Y��̿h�A=�H-��[��ܶ��V>&��S������!>�W'���OCm�i;�[8_C�:���w�7a�=�.����?�B(@�d�quNK|� �d"	gߋ^�Q��k�I|ڡ�=H�xY4�C;�:���U�^1ϊ[�>�le�Ĕ#���	˺"RЩh7�ju��hv@��gr��q��tg� ��%&WF�`\Yc�"�����k�F3���U���� ��GףԱ� ��&��h۔@��&:�]��0�U��0Ƀ+��ǿʑ4������o��2����7����v�,Z2�_��}��+"���)9��AeJ���"Ave��)�cƳcUO��K�;ߟ�B0N�LY�)�Bܙ�?� �CK��UR��S�ᆠoa
J$�f<��}�t�	��@�:�s��{���~I�j�3}�Q�zA�_A�ZՓe�X��O5]�ϔ�A/��O��#z[V����CPહ9���1�_-(ٜ�4�,��|�4X��c4 ��SC�DkR�Q+�gy�c��n���&K���@���Y�"a���DQ�gD�ښ�B��'Vz�[r�άlƔ�ڛ��	O����"~�HEk�5)����[�}���eذ+ͲM� c��H)l�Jk	�/�>Co��3�1���iP���qy҆(�X�=w.[9����dP����C(羋\�uE������mT�d��gػ��dmC8mt)��Ga�u�d�W�Ef��Qt�s��Fq)l7�ABYzg�G�����u��cEkp���n�oo��gm�1K��d�
�	��iU����d���t`���]��ؾ��%����O<��}xp��j�aP���%��짼�����#i;_���ˁӮ�����-M���j��\ꎥ)���&Q�	�t?v���w:?�fU�c��V�Ns�U��
�φ)WV��)�Q��w�ߵM2Tǌ�ɀkG�\����|"��D�N�����I��+��Fw���i�X�����2dx�Ixr�{�u�����X���(3<�m�v�},h���g�P^�S�4`\�%�Ļ���"��T��z些֥E��	+��2�@��<��l�[,���#�֨��.(>����ulI�lK'�.{#�N�"�WW�M�*Ͳt}�EZ��T�}����R����ܝ�޾��y��f�Io�������Ic����Fa�/~���a�g������~���f+#ڭ��r3�l����+�i/"�ve��*e����(?Ö�n�^ۡ��`�]�9��i��0�ç����X�4��b����z���h�rT����,⑆0�oߊe5���L?sr:u/������BE�+i�+Ddt��5������o*�>j��d5�'�&����U���
t��jN�1�e��	�p�'{�Г���ȇ��Wu���"�Ƙ���=�a!�'����-p��o"&8�iN�?�ntQ8{��@��N̕�Dv=�h��zyWL��;HGP6�O��l` ��4A����5={8���9�2R~l��c-���<�P�n-�]#��W+��tv���Gj��)�/��lx���g�O��~DO�k���T�j �i,��w�$^�����8��3-�JzL�߉ҁ�36�6��<4o��Tw��2��E#`���~>�!���`�Fc����0�>Q�rw�#���k�.۩i���DV}߭.��7߳}�t�c��>G�fr�ٰgq��y�B�.�Z��7 ����9�Zs+��W(س�+���ZhA�/��hyK�k��&���2m �"}�4�y ��o\������]M��i) ����z����Ŋ���SQ!J�k�P]�n��x���7	� ���_'8�6C]�1Y����0a��x��`��o)��9���f�v�f���!RF2�cL$���ro6?�aD�����Gj���k��}m���*������G+�<s/�,y�,�Q. �2�,��ߛŀ�[�Xf:稀��R��W��H1��/؏�2��2>�_�8!�0�\^�0
+��ĔIp@��,�Ҫ)�N�~A�N���&K�I�>	$���|u�G��z|�aiB��1@|��,�n�igc�mmk�aR9M���i�W��'@��[��51�/N��<Z������*�"�d��t�¿�R��@�T�Ѕ��j��*sV"o�/�m�%j	P���$�/������:����Dk��A�������s47OCC�! ��i�wX��d�<�⹫G2�N&-�UG��ޅ܎ٱ8w
T��;�f��ۯ�K�"�V{�}�K�`Y>L@�!AZ	7w��o4���Q��@Y�j-�<�ya��'���.2�$�?=�׳S��[�KuЦ�%R�d�(��9ΑOO�-���B�7c��P?I.�T�	��;�k5���K��fR�[4�f6Wb�r��
��\��j�26�!� 
�#��O���'����SA��t����-+h�dU�{�h-N�}+����9؍��Z�u$Y@V0\$������gb��8��;��,���9�&�öӾC�R�A�'��ֿ�HVt~.J���g?��B0�XX�`���xH���֭��a�aa��`X�Ba�=�$N�Ps�����6<����? �]w�^�mf7���U*����q�~�4"Q�e㕽KK�>��� ��{ڝ	pǿ���C��$�ZwYzL�q�m�(���X�]�?�i����W�r2�5�������-��xU�i�o+��`�b���)��6��$��� ���Rf��)-�2���n����3a�hm���-1�T�BS������N���2�_������w�vl����l�����a��ks�^1��=��)i���$��ع�������X4c�pC�4�Ho���}my�����+@�vB��.e�V{��(��
���ܬ���)���9�+{�any��B���_���+��z�l�E=`s����!k�Y��_��[\8)j�_��p���UE���s9zԑ*e����#u�2Ξ��?J�[� �	�kJ��嫪=C�\\���d��A֢�����rXረ���F�b:����%f�u�{�TY-a���,Am�k�@K�!��[�{���!Jԕ˚D��޽��@�oz� ��< ��Ni��v�M���	L���M���������"��䇝_VET��lc��;$i5�i*�,���g�mƨ���rڹd�v���i�Gͥ���������	�n�	�f�6��m�)�F�-�N��.��6�k�ҏ`�>�{���`�q�׾Qgb���|�`�$}����=���dP����=iwゔ�޿�}LGFhh��N&@%|�{�ZSq�ɬfE�D�$���B��+V{QU�����Yŋ \Z�#����m���0j�6�;�21�t,��4�1=������F�a�2�۞o�������+�ʤ�=��:�`�됽ոהȎP��ǮK�O"d�\�q�L�*q�D���Aw~�ugCN?�^a���I��oÙ*(V��ه��9'���{�j�)�<�;�_�PiM�P�MJ��ن�A�P�H�^��`�)%��\���D�1�C�،�`��MM���Q/�/���o$P��%5K��;�B"�ɓ�{\�*��_׈`Uc:B�L�\��x��HVL���%s��e�_�?{��Jb� ��R,��-� eS�э��&LTm�%o���ļ3����~r��}|��'�P.HE�O�'������#�B|D�6h#�)��
������/�L�ká�M����D)M�g�#���F`]������i��F�o���h���R�|q�%�|9�ݯ��j�!M�r����AҪ���V��;c/3!T?&5u\X�=����7�>~�	�)�0�O��5Z����R��l1������S�g�-����W�'�������Lw��~Ҩ���>���T=��%����X�C������C��4��oS!�kxn�ƚܹ���%@�c��"�,���W��ǆ�C�*&L���k���.�Y�{Eť���9�$�ۉ�dm�U�)�i�0`M����X_Ǭ+��GǩJ�� ]\����	R��h�`0��Z����a�H��F�\~�j[t�%B��s	� 8p��*U�"IL�+�n�Pb�ML�4���P���+�n�Z��[���̶σ*�slI�x�u }�/�9/�3qZ��EJԹ�A���bA� �9~K+u���Q�� �i��q��0��D���@�!���q=[�P�ˎ�t.vҵn���3v{�i]P\G.{���O!����f��E�Ǝ�*�lO�n(`������W ��ҁ��G^+�Vw	/x��͕��"�;J��C-���~Ǆ�Ze&�[9��rخ'����B�T�^��)O${���*|�ɋ�U>�(e���:W���܈e/�`X=Y����9���O�{�c�OՇ� ���E������2Q{��X����?8�A�����^(��)��p(U5�EWn?~��rP���!O>�y��a]��W+Wf�'�z�"hc�h���
�-�=�NS��J��L��;&FS�~=�Ϋ���բZ�I~���Bĝ����Sʦt�\�K[v��/o�aaB�y)��4��g�5R=ਖ਼=��(����I�JA�K'4��c���%�yg�h�T����١��\������h� ���u �t�s簹<�#��{TF��t�j��X���8�V��R���ȞY�ZU�R~F�ҹ�n{Yn_�
]�� b^�$������مCC;��c�+Jx9e�x��NM���e�������ژ�]���'T�({��_��e��|������wE��C��u
�Hk�и�o�O��z�Ğ��y/�*d��1I��ƫ~�P��o4����\�K�N\�I���Ι�l�c4�f̑�9�1��^� ['��]��l\����UK/St�Q�,�:� }�t�O�1���>i=�8ȣ�ؽ>�.��f�aX.��W.��y�-v���z�Gfn�d�+Aοo׊Z)�~�W�Z|L���7�a�Jg�u�~��7 �c���lNH$x���y>��^�#'W�H���*��jO
�cU9��p���RեT�f�00�l���*)�:��.����.�0��:��Æf$�7��Z��&	Y�.C�|�z^��59��a�	�J�_ꀻCDxk����a��iљb�)7��VApu�%�0e/�ӣ8{M_KV����������{-̥#X�?
�~;4�������-S�\���c�R���F]7tZ��1�-�|���C���؎�v@)�ե��!yJ��\���N�oD���r��`P�l�D���Yl��Q	�}x�1�(誻�K�f����o@��彖>�fy�s�Z�l�J�ʧ��xy#�	�D���l��c�H�}q,� A?���^� ���uZ��z�;G��ѝL��Sl*8'X���	FZ~_�g 5�Ju@t�,�Qy��C���v��A�|%��t��z��i�,��d���A�UF1C�7���E���ѹ����&����T\�:��AU?})2! ��~+Ԕ��3�Põ,��-5��BH-E�Iclq샑���<4U�&�u���6=���m*��^�:���$n��pKq{�}�S�b�R�����opF���"�K�(�?�;���k(bwKXJq�=c��v�}�(�l��ڏt��m�L����E�^�a��c����S�z�x�^����[B��ꦵ����ϓԺ$ڻ�Mt*������|�u�{�V�V�U>!}i��U�L�@����>%�kyv��}�A�v6\Ǵľ�A8��gt0�Y��F;Xu��R�kQza�%��0MZ��5])��֠�e��y�u �cB�ƾ�)�߁E��}]@���#m��������CD����I1Ih�!~{�3�;9��5QI�Ю��m��J��M%�0( ��m������7�?ʦ�b��/^�7����R����;|�lI��D_�/6I��]�������y^b�L���i��4����7qz����3���{�����{�۶꩜��*�Y��T��m��Hf�sN��,�%b���_Ӆ#/���S\!h��Br/Z���ngd9<�d �,�4�5$e���!W;?	[���H'+��Ry��{ -�:�*��<#��|�A���xe�KI�\���¢\���B���43��2B�V��>ZC	%�H^!��dbD�-9L�L��mEI�V]��>�A���?l�Ϥ=`*ض�LR�5�~X),�A�tn��ױ��kG�"��h+��*1�b���/���9�wʹآ�i��q�ҧ�Y�BZ�j�e	��ŀ�Yݬ���b�q��#�f�."������Np���toL{rߏ�L���[�P�)<�`��i���V���I�+D��³�4���q�o����"2GΑ�X�1�w�R;���PN�L����ϮV�����P��pv7�Q��r[�_Gn5��	At-�J��$tg�|~�$��k9�~�4	�w{69EMz���֋�T08���R!~$k)B�7�Ҷ�5�o*	q��-7^�Ⱓ��~��=C:��F�LVmU�F���˭�ݾq\bI��oz����P������#R�6{��;�P��{b�7Y�YF���q��e��մî"?�n�$�I>����VC�,v�����6�m��0������ Crv���e�y�e�/ҋ�DIA�t�k&��k9O�d��b��u~�#�`f�Z�OH�w_�#�CUi���w^�}چ����/�!��j1�P�p�PtG�r�i�S����hKG��/*8�� ��`��j��@���6,�|�u�u��P���?�m��mQ֔�1���!�lem��i������"��,�NWئ���.�Ns��fōa�6���ߛ?��tI�Z�IrV�yj��1��!6W����6���Nx���2�sD��/�b����nn�b
	q��Q�'��_�`G�h���o�ǯ+ə��ِ�y2AA��������ʧf6�iy6H���g���-�.��dL۳J��u���W-�ÄL�î��cR}%��-��H����#�-Z��K]�]�1�Ei�P��9���A`�hg�ۮ�f����VzGRV1��To��}�)�^��W�t����D��ޱ���]����O�
���+�u�P�nlp�
��ßJ��m�����]�{� ~�9I�o�]V=�wi����722� /�n]���[U�e�Y��l�[ե��OOY�[�[�;��p.�o�ٹJ̅@�>����	�m	s$w�*�\��i��p���Ff��[)_�P	)v�'O��Jv��l�N�EV�UM�*�;zӝ��.+?���iD)X���Ok_d���eoJ�*wV�S@�g��E��L%�߰�:�0�K��,���k�Z�랢
드����:d娎|_6@�S��G�-�I��{}�X��1dq4��� x&�!��=�����q!`e;�sy�b\D��;���^�y���&�'�N�(!cBT�X��mc��%-gQ�*��i��J�r���4����vр5��t�!L����QV �0F����:Z,��Yus�_�(f��J� Y}�O|�@�Q6�����!��!�	��66���!��y� ���Y>#n7{x��j>mV�u�J��$'��݁���b�٤��f�����~p�hn"A�=��a��1�x$E�G�Q{�/0�	uε���2�s�0��mPf-���BuP� q���ՃyA����#q�@��u?>��0�uެ3�?|N��,��~������6 �<h܏���<F�F����5�-�[�
=�/� ^(�7���X���_������'CY3�_þ�nYr��+F�o|
��O]K�&J��g�/=K`�wp���!�ƹ��:��k�FG�����\ϝp4���ҷ�'�ΪU�5�N���Ц��*��h���������؝���^g���0�!Z�eDk�& �tZ�[oIM�5Ws7�AG�=o�Qϲ���}#�@Q�؄�JIϷֽ5�z�3�~s�O��箂&5�'�|5��o���j<�9��lW��=�!��|�a�=�=�5��CI!�>�==ȻwX�i����WN&,}5,�!�S!�\<�`��e��f�����&X>��P��������;iG�3�ڦ�C�`h+���M�d�������F����cb����_��b w��,WDQS�������������S�����k��VK�aÒ0��!CZA�(G	��,��Х��t"�CF���М��:�>Q9~��
����m!���MP
�|D��ﶗ�Gy���a%�!z`����}yg)��%�0e0��<2ŧ�:xD ��_�����C�Y�����+�p���(W]�6	J�,p��?�<Փ�^y|@���p)1*s$	@9�Z�0�"�8�H#o�_�h�=~��7�F,F1%�xHd������	�G3{{ɜ5nV�K�Z����d1�b�׳�����$y��ݥ�t2_M�?-Đ� T�*����I�WAEs_����#��]�>��͖���wz$��|1�Ym! [6���a�n�_������?H�T�A,S��mda}��˃�V�ê�nt�Op8e�@κ�_�&�/�@����C=N�l)����IsF%O�&�O�.��9�pWs� �`�X��	�MHG��!%O@>7Zxv���t�7�32I83��j��a�_eM,k�(���}��Wz=(w�� �6b�#X������[�J�I�����Zu�}`�s�R0��̏��+EZn[>2խ��4!0[�����w1�=�������lL	��U�&�$�j�
I��gcG��Ÿ�3�Ӓ�{tJ����9i lD�ף�hε�u�E>�Ҏ6p0�&�L���joK�����5d4;�[�@B*M�-d`�� ^�O��,��%�R�1r�C�̕&��3���i�Pּ[����D�:�Ǭ!��o9~�l{��F:Y_ݶɹ����K�~(��[z�.��ɯ:o���kaa�|��+\8�I����"�R�?�xl4%��!�u��*F�H��7����s�w��%�Ul��������D��F��}�5z�XŽV����Y�7U�يS�w5uۍ�ڑ��Y�������.P! �$�9��Hu���UTG$���GxUX����2�h��U��3���c��7/��P�1����7����j�='�IL�ʤ���'��9���\B����P���6��q��]9�z�+����N�Bc�'�Pmj��*��R��v����4s�z�e�@�d�(���t�ӰK�	�N��b�Y�������v\5{���e�i�J�k9)Z����Zr":*���c�	���'�G�Y�gP�	7h$o��5���x\k	L&j�A4��2l��K�3���f���.�[)aix�2�h�$�^��D�4)�K��N@{�]&�a�E���J(HlI����pu3G��T�DK�:<�ʙ��|�`��Q��m�����d���Bxg�\4���4^�⥿����\p=�a�WD-{G�I��az��M�#�v ۝��kk��V�ve�d߈e�)��y'���w�@�b�%���ɡ"��+�rS�fj�L���U���y᳣��Q jg!m�M�����d9��2o�ԙ�,���
�ڧ݊S�I5� stA)O��]�sV]����ۀr׀�f���W�}I��1�Q���IYT�&�o�6�]�t-��Dg�AO�Ҥ	�ev� �	�6�z��r����.���[�ݘh�9��[�Ϫ�31m7:�X�"�g�T�[�}�A�N�#��` �a��ĽIM�I!�*��TttXF{lw�R�*��Yi�z�>`f�Rc_�^�+���H���1�8�'���3O��N%ƹ��\
�� %D�R-h�����,q'@w\G"���T�u����U�����m_TX7ž�}^xz^;҅�B+>5Dr���R�`e,M��ku0ǔ�� �.��0g��}���o`��οj���@��w@�)�9��?���ǆ��Oj��y� \�ꏂ=�F��[<�^�b��".��<���|�8Vmː.�Hi��{uuN��I���Fd�6�����ȉ)F%���q礰��t&�<Q��>p�C�n����͹+zq�O.����k�����%��1���VF���̓ʝ��I�(�1�����ND�1�jh��e���o+���X��߭�8��P3 h�xfGV���5C�[���_(g\��Ug%���܍�(��� �S:x�qP-�q���\���X�X�i�H�!�&�S�Z���;�����B"�D��c�`�?��</O_\��|�:���V��*�J��n�����7AJ�$G ͐��À��.=5�2/۠����<��y��-��m:.;`��r�|�=�\�࿢"��������)-]Kw��'e�!Mo��@��C-j��*-����:�SL��p�c
�\��	�8�CK��;�ek���z���ws,��e���Jf�fɈL�R��
:{_^�؅ǌc8 ��I��R#�T|f��$��gdgJrȉ*�j���~Tg^����e(L]����(5�5:���׸8�쳋e��܄����u�0;!���+ʍY8�<��ד��W�����t�͕�k|��*�����^�r�t�C��r�_\2��Ll��0ɍ���j�,�er���-��2�rׁ���T�c=:��I�Ko���<���v���/lV���<����I�M?>���$3����hPQ-v΅�,�ޖ���'���d���D���⺧�Q�s�0i�'S�f�HYq��V�E�)WBhf)�Qr����C�&����2�c>�S��gZQ1�3�'�OTu���z�X�2vIg�ef���Af~�:.z[�Q�Mo���^A��x����)r� ����]��,0����H)�hKh�^Y~�;�"D��c��ê�5ttkğ�Gd@��DB��*>�]�#��iߛU�t%���L��3	S�/6-��Fe��[4���\x�^R�J�/G˷@�r����x^�p��>Y�*�<,4ց&���Y�ʰ�'�|`��˷C=�1��A�5�ܿ�J*;���ĺ:��~)#��G "���̃�*�S�fCS�ɺ~02��.R8C�y����w��>[ZJٜR?T�\r�O��p���|��t��h[���� ���2\A�iVe� D�׎�
����7S%�N�$zh=u*�����:=��/���'NC�c��'�N�w/�+�$j1NH�_ȂGR>�4^�{� �ؾ����e^�D�����p�I���x��A;\^�YGk9"m+���.m�p���/��	��h�դ'P��m����y��v�] <�z�!�	�[��W��S3�QX�'����_�v`2[.j����'2����kG5<�ܪy�"����x]S�p.Ӛ����2`B-�k�m�	�׌���"̀����*�ݵZK�,k��L���U���~!�Y��6#L��W�T���K"�ӷy*�v���z�v�<�K�l�2BMygS/�E�ׁ���9�|��BtU`^v���h�)��ds��H�+*.�ER%q~ 28�	����������û~p�^&�%�?�z\9#��ʄ�,�J�u���0E���`������1�(c>k,��T�X^�WXl��g�^ŗB�X�>�Ԏ�Q�'
g���E����aP怷 ý"����na�:��_�� ���͹$�����Z��9*O�z��5l�6פ�% ��>Ɂ9'"gL�Q � �BQ >k�Q=Se��f41�Z|����/�J�� �r�߉�t�y�5��0��rA�R���9)6A�@���1���f�/q؁vF�qr�%�;�������دI+jҾ�J[�7OF�.e���@:.�sd�WEa���Mr1t��*�� ~�;��𘸗F) �p��>�h��d���c+��
�@:;����ֈj�li�7��Ej��� q!�;��3&A�Ob��5Լ�^$������&����>��~�ѭ$�>r��Zя^!W.��^��/fzJ�]�*��
�Yզ{�`$8x��<܁"|�,Q��L��+�b���t����:C����B_	��J^�9�ܔ���ǈRud�n��ڀ(���k�"jӁ���~B�`�H�M�D�>1s������(g��~AC�;�!�شN�htfe���r�K�0h
�j[x��S[Zۮ6 n�!ܵ�~eIAs�`����^	`n����S��Pq�g�	%��C��4<?Fx�dA�����WW��M��NG��8���'ͱDv�DX� 	��Ћ}1�F^�O�]vT���R��g�9[�ԏ���FY�W
�� ���4�4���/	�&�|Y���F�u���J��o��lf�O�U�R���b�n�B�>�Z��J�J�G�p@������׳�G�Э~`�k|<Z`�/�(�;Dw�=n�q�����SdF�6��B�s\����z����z��V��bVFق�*-��"��_�FE�Vc%c�+{A-7��FwG���{@q��o�X�?ϙ .�P*�n���¿R�ܿ�=<i���ə�\�t��L	K߼V!�����}�rO�ͩ����RD��<�)ڬŌ)���{*c�� �J��C�������Z^/�S���u?��*;ES��)`f�)�AR��L��[�Zۧ`���x�C(�֊u@����}�R�d:����_pu���s~vc=00�Q��4Z9��?��l`
�&̕��R@�#����C�aܴ���n�u?�E�������r���-8�����l-��Y��ٵ�"�S�����Ql��7;�<����+C|���&�[�L�=����%�L0!?���k��D�ǽb�e�l�v�abՂ�%�>��S��H� -��M2|���5t����L��3%4��np(�O�xX����Gt$�)�����J��WG�*In�M�g#��0E���F+�QJ�/FW�f撅cΪ�F�CT���|.|�r�u�c��FxZE��
:#_��[n�~����'-�q��xh��<.��L��*Q��!���<1`ҽl�^������hA�3������Ě�Uc�ڬ����Vĳ	��ɲs��Z�%�[8�|�tb4�A���<�\��y`�L Q�Q�mm���~����@	��詯�BPC��;H�v��f�'&��d��аnJs+eϗ���Z�P�Nñr�½�*Y�$�tz�c����	��4����2��lT<S���cZ�6�1�B"�GhZ�V�bv���_r1D�G�s�(������3�l��58��/���YO�
�ב!�#��c�V#�r�\?��)�W,Wn��ߒ���'�F�jO�s'�_�Mj�2�#LmU{Q�����k�a�ЍԉY|�~��T2=mR;��t�{��9�E1c���W���U"��ňN��f�����o%�y������2�1(�Fx�눩ȑ.�S�~���bЛ2ȉo�`׃!nR�����'O�I��;h!x` �/�-���[���*̲��n�/��w�&f�����P9l l�y��O/��՘����[�WZ���(�x`��,�s���!�;�y~��(����J&xh�mD�խM^x¦#fGK{n|� Rw:�����ܜ1�{a?Gy^YtC�R�����̼WB5��W�If��r��>-t��U�YfgA�ɣ���U�Y��k�DWP���\�E��c�(�����/�EG�P�p�	��������Y��Z�+�6�e-�+z��&,�?N�����3~��K/1 .��#��c�Xޮ��*���4��[���j����3!x �i0"LU+k2�R�-[�ͣ���ԠM�Ge�㌓-�wq9�}�?B*��ìVy��'�Ґ_?bT�l��zB��6�g.R&ae'J�E2�80�.Kb5�y?���h� ��y �9���]��T~�2F���c�~f���Hxycԗ���2q�G�P��Eԍ������F��C��m��Hж���z�v�ȩ����^z;H��鴽+X�"Dn�/#j���7D����U����5���E�%��?{���0��8����!���	�i8�3zL@LA�wLQ}wq9��2f�ˌs&>�C���?�R7�9�����q��}~���,�E���fo�BBw���h?���\Ҿl��Dt�pR�9@H��1i]ϝ8��M�ɋ9�,?��FV��){��^��g�[z=)��",#�`UA��5f	f����z��L��k���]p<N�l�F�0F��L.��!�Qc��T >�A|O���b\^�Ogi�ߎ�@Ω��)�6יɍw�}L̩֐sh������$�tܧ� �%���c�h��$�{&��f��ͻa��.�h�RC�md43'�d��?X�{R�ޛ�O7T*��yI����ks^�g�D�%�1{O~����� r���wI��!L*���Z�5����z[5�(��)�@[���N�Z�<M��%����g�X	/��9�:Kd��.�4H��A��՚d���@�~oX�_�<�?/�N����"���"bW�V��N��YŰ�XY�<YpA��\����J�'u��Ze��͑p���������J�^[f�D`������"9�pi�7g���0DS�1
��흰 �}�[�O6x�:o��n��q���(V��Ud�'9G���LV��:�Ȼ]�H�[�;�#(_�E;6BN�H���D���{ŗS�g��a�G�V2k/*�,C?�@�0f�#�������%�|�]����Pt��UP�����DL�[v��8�Zp@��t#҄?��5ѓ��vΪ�%(�f�X��6:)�w�׿�`�!�񘒘�u-�T�2S��ҽ�<V�Ґ��Ϳz��Ώ���ڊ�W{Z��D2��]��E����YDm�}Xcݚ%�����o�������ڥ�ڷ5]��q�Z�C퍻�5bVn�4�����E	0p�7)�l�
�Y��POw�p�Hْ��S�m����ځ�E�� ��9T��j�i3���V�;��r��K�n��K��Z{M�{��}�xJ�1��g��]ފs��G���ǻ'�%x��nF:{u[�| "����CF�]@'���H/��Zh=�Z�~�����a徙ş4�
@Sz8'h�3��}	_�^�KؽZ!ΰ����t-@+{ξ�,�=z�����j�-�r[�lۈ��ӓ���(o/�s�uyE�n��`D�%�3�Zn�DD?�/�[�Wz���
yg���*%c�uC�pϧ�Jޛ}')gF+q��,�#w�D�`�ZG2��*BxIĎ������������d�(�&U����?��2z��ҹ��PD�'Y��(o�)�q�Y�����+��*K�9ۉx��| %O>��YP���7�F0IH2"�Omw*%�S6�F�b0��Hs��K��=��6�������M����Bo9����=��-%��\WUX`��ݜI��Jk;�Y���a��4���0��C������]LNl���֠��]�,���콈�r�C�F��f;�n�R�"G�N�d���aMl������>��Rm�Q3ܙl�&[��Ѐd��+���ٮ��鋼�g�cOrO�T*YV^�\>%s^��:�q���o�c9���E�籭-�n������"��ېT:?���@7Sb�x�F�ƻn��
���Th܄�O{z�g.�@�AӮsܨ6�t�Ān>�딀X��8]7,<#e��@1W�����@0�Q��[��%@C�S3�߶�ϝ[�r�L��<m�*���ZV�T��b"�k?�n����Ŗ	V���������n$4(_��D�fٗ��Ĕ��n���E���'���\'���Y�m���.���4�9'��Z^d���.4���9��<��&�pG^W�B	��o�ȧ>�����S��X�L�¼�
��B�/��0����H��@I	�� ��K�ٱ .?�F-/e���h���~
�����������ݜ�X|�~ܧ"�d4F���eor��׭�
uhkR"�b��#h[��۾���I ������jw���b:�%U;��6����hը/�~&"�[��-t�.�5�{�|��@XcS�I�	q(:�Ƭ���w��G{�_(����zrӛ��Ajp�O�+�~O�`-8�	g55?Ү3S̜�]�wA�$xf�\K��c�iY!��.w'+)�ħ��dԬvܼ��#����AO��S΄�i6.�2���ҪX ��h�qHk.�v�ɓ�,)j>����	��I[�h;�[�ꔐ���d��!�d&"�����)ZQIH���.n�}/9W���ǒ��5�hԸC�\�}EBW�@E��(�i�Hd�ޡ�\�&�@��g4�J�.��T.�T�7;�e� qi�p7�*4�F��!��ܪQ�H�,h��-Ɠ����c%�x� f�r-��&�h�n��J����3�,� ��³v��[�Q�%As��:�
Ya�`�R`�g��i�����r�F�����F����R�H@�k�sm�.̭���+Sw1,БG=?���<~Vf�������d�F���?r7�/����T�j����*/�d�q��i��)an~��JЃN����I��3����z�����P!Z#@�zz�Q�Ap3�������jܻ�bob�FI�o^�Q�Pnj*��A�Z0di���e�M+��n�<3�j����dg��j���K��My뭭嘢5�w�Yf"���m�}����I�aj;*��<������㔷���W�7V3��/i�����˾\*ލ�8m���1�/Hb���x���r�a��X�9��t���Ş`�N�@�oh^��6p� ��ƿ�B���f�w�T2�f����D���R�H՜�5��}J�8~5�ZX�e�����B�f
��\Uz�r�v;n�T1y��"��r���~���%)����۟$�D�E���8�g_�}�/�h)>2�#]v�$��S�RA�1�c���J�X�PXZH�Y��*91�����h,,�'\�gJ|�Z�7x����ᲝM�,��?�/�g�݌Q��u/BoY*]������ �H�����"�\Ĉ���T3puj\c��F�x�!]O4��N�}b� W{��L����MfB�v/����2���5�F�{W顐5j��vӧ�w-젮���kɼJC'R�mj�g�i�	=�y,�����t7O	�6�<���Y~���������i�)\���c���w�ݘ�K����9�?�aWT/g�(��VT9���	��c�����݃��mҘʆ'WܟW��2��YU���U��	�N���������W�����"��i��D���x�,��G\{���o�7qb��7��ah�)?~��G|���}l��c�m����2d4��1���ZY�3�����g���y�,����#���P�w;�����&%.������4!
J�=��cj7�,
�SZ+B�1exPc*S�8hiC�,��u���xI��"Cn�R/m��N�f�U�^�MY|-N�!}?[L�6=K3��.|�E�����$��I�l��HPL}Aӫ��P�� 2I�XZ��M^��l,ʚ霃�䁻g��x�v�����݂���'�"��>��Y���ld���yC;�-m�[�؟s.N#?�t��nj2q��3�OVѿ���+� e���K������X$�<IuT��$<�D@� ��o)�(��Յ��Gr	����F��O��9e��*�ܽ��ۧ!��E��~�xX�5�Q��c?i��oX{�搓���`�*�P��et���g�0.�#h�#��r���;�D�c�L�f��0Q��+U�
�D�_y�F�<��l��`]W��@怳O`| �<g��Xߵ�����b>��:>C 9u�zS�ŉ! ی����i�;H�B����&y���SĜJ[R	�w�( s �=�8��jݺz�q��6
�����{����S��H��n�}-�c9Չ�Ghf�P��FuCd�2�������'B��=�3v?��ލ�	_.�+��d��ydDż�w5pմp!��12�EG�ޠ#;ַ�(�xhxf' �ˢ�[�y�}m*5������-<�g<�b�/+����^8��F��|	;��1�����<��ڭ_��&�!�ЈĲ��g׷6��9�*�i��X�E����S�tz���b��*�_AwxòY��&U��>�O��U�D�U��fY��M!��ۘ�T��x:Q�գ����{U����G�cx�.cZ-��`By�+Wo��ʻV�_"�Ưh1@�2�/od�e̋�5z+�z��Zu���<��HY�;���H�f���3 �@X�5�:��vU~m�т�����(�B��m�b@r��)�y	Q��'A?/���s�IK�m#ò��H@�<b�c@�_B�Dj���ry����Al�TZ�8HJ����/�*]f����ƌ�yGcYjCS5Ksa5)�=䮄�Ѐ��`����>��i�YR��pΏ.h��I�mz�s�)�<�>���Hu.��$�A�����_���gV�I�����V�n��Ϋ~\)����#y�d�I�YE;��1���N���R��(��� ���踹�sy�m���	dJ�{�#P�7)�H�(Fd|2J����!��/��DA3"�o����!|U�e,�0�ћ�����)��y�SY��Ra�U��4;��J�34�H��4�6�7��,�1em�2:��y�Z�,���pX�CwDsΕ�\p�8��u�;6n������%Q3N��N{2��*� ���&�Vb�m,߷�b��h����{�o���/:�ՉDI	��'SB��x��~ B��%�U�}IU�
�=����>�2\�䐫�Wr]7�ru��{ӧ#�tEbϑ�֋��,�"��~��Ou#Eg,��I��2G�ƭʢ	���6y�[����K�~�����Zf��b�ț�Dǥ?H���d�Af�f%��:�5HH�-(Kف��;{�W������t�BJ�_�h�-�>	Mǐ����^T������9Mf�@��ƶ)B�l1v�Rб�ߎ�R��\�}����߭���^!����M��ݱ���ŋ�1U�JI(�>�#:ls~ZA�4���\.� �ީ���2D�f�.F�����g��1-d6�hr����V�v،�9���2�� >4�mX��h��V�+j�����k��\��&�k�i�8F���oV���k���'��]�%�'���������l#8��aA�SҲ��n�W�R�����=�#o?�	��
�%}��.��{N�~�F�h�V�`t�������˕�Ԇ��S��%�R�lsZ�W���������K��n�
Ւs"�m��%iE�mAl-�G`$�!�Dӟ��a)��|����0�X�-�v�C{�����|�Pt������,��5��s�p/g;.�p���606�7�"Vr(�
"3f�,B����X5 ����	�l1�p�R�wM���~	&P�d�m���eI7�kQ�:Z#[Y��a��
g���8*wX��>#ya�5��+ь��?N��)���-pv�nhx�V���#hO�'NoFF�D���AYPnZ?}.}�ATg�qW��TG�$��=\����������Q_�.N��w�c��aέ`��~ѐߋ�ʕW9����mv��h��.�jNq�5��
A�&����;��k�GB�$M,-cE��_�uWԻ��8�Bm}6s�� x�1��Q�ͤߔ7��l����Ur�{�D*di:<�a��A�`��UC=c��֩Dn���2��u����9��
��
�{
仨%fkă kᰣ��v��{ݰ����bM���:�#�.�t�D��b,�ePK�-@����S�֬l ǳ0�?��;���.O\�$tQc.7)4�<���J�������ɾ��	ᄩ��{��g�[��ǝq���*G���F���S�(�M�����T՛����Q ������K�m')?f\l"
�~���0�Y�_r�(����|�0^�H�����K�����󐖮�H��f�4c��~��"�:b6�G��ī���L��[���rU�?�=�9N1 �z|�H��G����
����u�����y)љ������|e0�� �9�<��/pp)�/�a� )2�$�d�է#3G+XTs���p)�{��	O�\�Q�F"�I�:#�l�3SA5�^K/�]�-�g�V�h�Y�͊+��N%�~T�~��a��e�7ж�Y$��0�3�q}S?z�t��z���SY��J7k�5O��|\Et&.U��wM���V�j҉�QQ�n�����ȴ��xҰ����滘�xW*����N
=d|^��n�@���vS(���#y?r�RB쯧�F&�ZՋ�xM�y�*t��;/h�j�>N��a�%��K����g�C*d�ޔ��@#J�1.�;h];��Tlj�>:����+��0�H�������q���2�:��+Ib��ݨW"#;�f2Qr�����Z{��)��l�����_��� h⢒3��/ĝKټ���D/cML��a��LT���5E�xB֦&�x�,[�L<�	���~�����v5�)\�����:�/{�Y¾�e�⍙�S�������H��N2&�Mcy�}�.��t�S�y=m�g�9Sl�$��W�/��i�Kdb�����w�#�?U��u���}|�u5eR��uE�E�