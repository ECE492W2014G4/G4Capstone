��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�"��F9s�`&���a�oq���F�g�O�]�<ݲ����eCL��D���{�5��8̝DFI��Zp\m|Q��
�}�6C���UnF:<�jΈ�2�����<����sf�k��,jڙ�����2��X��Ss�HL��	�������+g?���N�Ż�����|�v7�{M��VNB
��Rs�゙�Ld\��X�'��R :�J���^�����kMkx�Q���3!P}�e���Z�Y?.�U{�RP	�)��lI{tI(S
7ZFhXg�wW���l���|i��p��:�������ƂyҚq�4�t�!��L���U����v���YR��8�9�s���{��E1�O�j��숯>�Q��B��r����LkJ%�|���9�J֍}�_��V��PW0�-X� �(r�iX�x��(ū{H1��������OD�7;&�7���%4�AL��@
oq�?�Z�~��	�V"l��Z�S!��X�~(�ܮr��=����4ϋt��$�+��>� y�1J
m�(1SOn���5`���g���D�er&�ƴۼ��ݸ-��i��ZL˞���Fl�W� H�1�n���enǑ˨�XK���=��?���Ք#z���ِ��7�W\�|���<	�ޅrQK���/��sX����)�<,��x��D�U�	}pP�I	��I�Fd��ԮFfX���.H�ٿd3��5�����ζ���ʡ�9���J�k3�X���vH����w�̚Ӄ�V���^�?b����6�cp�}��%�LHĸ+�KGt��J�^�)Q����w����6��_ji�you�4��X5Q�����O����͗�Z>r���B��I1\L-�
�a�������93X+ʡj��䍳�{��=g/�����0 ��+�-?ir`������-(?�{ �Jen##O�)��|ٔ*�i�}���S[�z@S��{$m�@P�7D]��W+8�0r���5.��>�J�O1 4��{N4��:�K���΋aQ<���*c�+t�ONT}�6���Q�Qo�C*�K�hi� ��#+�0)I��o�[�I��W�(�b�h�*�YD܆\����A�����4�8�rL�T�@t7�V��bfh`g��tY��k}�}/��)�/�����u�8=?�xxߛ�Ql3�@�*,T��`0�%1�����ڶ�{��;�B�75�n7��[��w^�~��[ai�0�/� ����{l�|�T�˓�J��4D��/����htF]ƀg��em��P.�L
:-��l6r&��1z�<�2��ꌦ?�l�8�V�6YҸm\ãT\iXf�k���!��O�%x~z8��s;�i��1)0��Nʡ�$� �S��C��ױ3����zVo5y����(�c�%���R�������eI�6x��x3��)��yn���3���:������<2�3NiM�pvr uc�̾:V�-��ߎZ�pB�,��d��~��*(���i1�a�ە��I��/E?��}"Y+���:�hr�3M�S���@��y�)�R6�{S~
I����S���P����p�48�l �f?�e�9�P�B�?���0���+�>[ƣ�ȩv{��W�-�<�ҥ����_e��U$	ǁo�������c�	?Ej�v��v��ϰH�(M�@c�x:Ct9R}�h֍-���*@�A@��aEu���h���Y���@oIx:| ߤ��P�댥�ou̜�p���l�b;E-%?�̱�@?y��D����6>�ƿ"�e�p��v�,�~-���^HuԾT7!TM��j0�YK9G��^�����͸����w9��Asv����{��mL�k=r����ı3~H�[�0����vz�&�Ԧ��g6u9�֫��{�y�����t�c �1fT��<)n�� 2����@��@�v�W��G~Kھ�⢷�Sq���>�/F@�
n�iS��nІl�1Di��o���ρ_"׬���v�W�u;����#0�� �[����4K`"���?cjF�"�Dj�)L�����&ly�&�#"{J�%2*=��ֆ8k�ix0�;�P\�uk�'���x�w��szh�8>{�b_��J�ӒJ���(g�"�s���V����&q{ۿZ�z��tA�����Ck?$F(T�f);93�u�a(>#X6}MT,e��l�Cɷ��� SX]vW�Z�L��%,pњ�3	����
��"��$����+6\I�Pp�Z��Ǘ�_�`�C&Z��h��3�)��Z�1g�s���]��)��^��¥-j�(�"L� �S��󭾿ol�玼�uh=��6g4��1�l���~�(3���@�����7�w�]/�l�w[1ju	6oЃ|��_&E����N�l논3xY+"%Q+B���Ւ��g�q� ��t�	�D��R�6~��Iџ=�(6$�%aE󠗔o��L�q3���m���7W���Y�~��y����-2+da1]#n�nQHP[\D��k?ˠ�n��V
aj_xu<`@<uǒ�d��)�J�]�_ �<�؋ӑ	��xCGԘ�h��m�T�6���US���5 '�s� �!��)��N���=yY͝�6Y$�3�^9���V���ǹU�s��0;)��@�g;�����:-��Z��-���[�BR��ނN��J��F��e�(K�/%ȁ�tO��q�i�ĴAZU�ǎ�J� �x)1�&�Y?����0d��P �A���G�jb��V!�J���0h��P�� �)�A���5:����������y.k	��s7��ɝn6�1u�Rul��F^�����@�Hv[�<l�����x&�T� ���^܍��C0��ʓ\��I���v;t�4³�W�Ъ��6J-x	��Ӊ��RO��I���{�����Ŋ�)���Q�rN|p��J@��B:����S�-	��"�ɩѹ��L����\'8c����#�YM��D��M�c��=awF4hðW\��e���ho���c4*/Z�dxd��T{�9���Zbac���Z3��5w)�3�n�M���2�]`VC��d��ƪ�;�o��"s�ّ*�R疋��O�i
�e|�n�1rf��rSgD1�|�%G���2���G�9�[���H�hurS]Ȍհ���g�
(X�Jui��A���瀃���ƞw����=�m�XMP�w�� !8>��Ii"�&�.�b�Y�%�����#�0;T1���ڐ>�d���;B.f��M�׍௹�����{��H��°ۍ��� �b����q�5�I�}�O(؂�pq��,��t�c#������T�e�PhfB�t�z���ـ\�%�f���͕�LӼ�:�VQ/@}�koz����6��\�j�h��9�Y�VZ��O~��/4�{Da�Ŗ{_�.��f�����cz ����TpM���tj�MwH�w���*Xr��Ę������9��)W�^ۻR�6�Mxp�.�ʡ(��Jw��k���+�`]9 ���H��}��;4�������9��gX��h�����S�ܾ�8(��$П����B?�K)}�ь�UE��	 ��M��:�ٱBC�@%
�VZ���1�	�����wO�K����/�l�.�� �%�[��[�RO/�#F��mV�a�����:n.�������pՏ��R�?Z��fI�)n��b�|f���YZ���v#��	佨�����L���G��ϫ'�8J����|�:��L�im{��F2-"$a ���$<ߦ"V�˺�~3�:s8�g��]���>�H���|1.tt��O;��bՅ��B�/��99�~�b�Q��OA�Ţ� �A�D[q��Q*'��KG���E?Ef8��xհs���a(��
�&0b=é����Ɓ�K���u���'{bX�k(!���^������ـyLU�O�O���hI�,[�D�'�ϫ�H򴣔#�z��������8�}}:?.����s���#v�봸CM��Ѥa�@_B��a4�?a\��шiZJb�k��\in|u~l�h������,�ud��f���L��u�ٍc�����@��7��	����/�I���5w֫���PpK?3�G�x�ȡJ�+7;��G+ם&�o��D`���gxݬUK(��\�Q.Nt*!KP�@M����;��\��GM2G}xm�%?�����PMիN:"���)�/�3T���v)���=E{�q�~YG��v��x:7���+LH0M�{W�AkD���Ԧ�v��r�Z�:�@�ZX�/��R���^�/��f*[��q��s�C�s�S:&�ڏG��097|��EK�ju?��v�z��P�.X��n�ʉ��yv'%r>��x�E�"6DDAܓ��r�W�k�?z�jN�oI�Z��2Ω)-��v,ʁ����^�E���(���3��N��b�a,��Y�/E�0;G^-e����^�p^�k�!�
FB��O!)k��X�^���~ʡ�(Z����l����� DJ�Ӽo�M���a�Io��f�:TkL`$�+(i�5�C�͢<�P��X������Ԋo�iA>$:	�]���I,%��k����n�8��q�O-lo���v���;��g�����w�ɕ@���q�,��p툌w5*���Ej��DmnY�i�W�4�d��U�G:��TY�@[�ܙd&}��F߿5O�h�(�6a�ab��W���������V�r�9�WsO��iӈ��^
�/�R3ٓ�)+�9m,��B����X�}*����*5d��TG��&��D0�q<*[��w�{s�����6�x2��pǢ�qeˋ��F�����A@����Y>dSY��$�޾�"f�C�m����m�*x����M~w2lxǛP�j] X�%���'p��J����ֹܫw�Z�e{�W���+؊���x����e)�m��R�C����%���d8ǌS��y��x�rO�י��f�X5S�tށ��h�_!����TB�Gq][L��鍼��YY,3Џ�OJ���C6�� ����ލzN3����S��מ( �u���/⢠F���(��n��3��P�ʶTw��E���5�f"DI{��u~�i��g��KBB���<��q�"yG��r����[M�ͤ�8�����!�a��<�R�o$�����i|6]���j�.���F�}u�W�7�ڥ�{Df9~ﲠ�vhd6��0!�(HDj�Y'_�r/^�d�E�q7%��:���|�F)�c�n��j��z#}f�N�>M$�o)�:g�J�S�Y��N��3���'���,vRo	�(9VX��y�|1l~�>h�wAm^]2��? ��x�6�(��9��4�:��ڛ�}�:qˠS�m��aq"�Eo
�*e��*u�,	+���y�w���(�0o;��h��5�ݓ�t�(�z����l �(��R��F�O�R�_%���As��&C)\1��#�,A�]�ϭ�� ͈D�+�6��B�+*0��/�<T`��%S���SJx�}Yli�|[>.f�OR���4��P&�FC��l4B�#���Ҹ#*��^h5_���BP�EU!��P"ӷ�؃�g=�g 8c�g���`��A&'v!ɵ�;����!T�$�N?Q�<Z"���:$@���=<-��sD������#���fP�d�/\��Ow�|_���R���	�����ɑ{(n�&[���%�M��{S��r�eiJ_&����W��:��wyp���cY;���C�Y��T.�政]R���y��ِⲁy���!�C�E��lV��f���&�9��+�F��8�ra��uAmg��YN�f��ϯ/��u��ҵ���+����F�:�o|q����j��+�y6%��"ܡirZ�L��#(~ �N� �{]Bx���w^)��cw��d�]�?��z���-38+�/�F��m�N���؀;���+��k��XX�g�2�S﹮:����Y{���6n��c��׃����e6a��C�v8��}QN�0g�\
���Da."�.��Xp0��K#8B/�W���6I��s���hhU�gy��*���z-��M�t>�hkUC%J1����"�����>E�lB?%h��<\��!ɒK\�[1%-+q�N8�8��XS'*aMx0y\�g����S��*B+
��|Z��Ql��;�t/�7l����}�dV;�OCW{�d��aȕ�&��� �f>Pk~���/۩y(/�&� 7����Gr`��ISf{�g��ބ2͠W>�N|���]����j�wj�K����%�ر�