��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�"��F9s�`&���a�oq���F�g�O�]�<ݲ����eCL��D���{�5��8̝DFI��Zp\m|Q��
�}�6C���UnF:<�jΈ�2�����<����sf�k��,jڙ�����2��X��Ss�HL��	�������+g?���N�Ż�����|�v7�{M��VNB
��Rs�゙�Ld\��X�'��R :�J���^�����kMkx�Q���3!P}�e���Z�Y?.�U{�RP	�)��lI{tI(S
7ZF�W+h���Jg�zoUB=��w\7���v���HO8���;�:��$_/�Z@x�*xC�eLg�$:��+����L��/(jQ�{����G���� ���##lf/^�i�\��2.�Q�-�8��-���Q��")�x��xxUb�e;r�~���	S��p[��,�]~V�,>�U9�8Oͣ�p]g����x&TLX�_��J�\�x�eZѣAg)���,�O�v�KNG_��~OD�b���N�4y���7䌭�`o7H���0���	"RC��[��m�߯�K WX��ؿY�}w��"3_�� #�C�߹N�O���-���(|�L{5ʱ�Q0�_��1��� �;Z�h��e�f"��S��Y�6j.ˮ_��;~:����ػ�5Ǡv�)]�[~[Q��U߬tT�7�~�P߼����)t�`��*���|j�M�*�%� �m��ڜ0�6`�;3��/�"�|B2ID� |�R� P�;j;F���	�t'��1�E2O��f�`[���ݠ�>��.�_�����C�sjO�=��J�����*M5ou���2#b(�u�| �v�j/!v8V�}�{�nTl�ܴ/{VT�S �J�L��s����Sq~Ǯ�,߃~�����3A��s�����K��l�\����q�Ǐ�g/���*<�U��U�Uq�u����<��iIj��"�ݼ��9%�;���Z%y/ۤ�_)�ym�tr�������N~�]�5/7{9]�j���" ӷ�;�vAX��|�^�W3�X��ّ%b�=r�^��U�X�y��r������
ѯ$$Z�&o��?� y�87:x
���z����r)����(@'�_�+�;��.���K��d�T'��Z,�M7.��O�ӱ�0��\�#�����B��I{�O|`?'pm�1e&��Bu'_��P�XK?�|����a�ь�a\��H��x�	Y���{V0�TbO3Q#�F6p�2O�FMU뿥���D�R��E�<�\^�?����+M^29��7�H����x�>4��֚5UDO�C�̴�@D�.,@�9��!�O�ډ��+N+�Z��Y�b�������0~�5�Nڰ-��~���,{7詛�9�B�99ê�! �a�.h��-�;yt�F�����f�'�up*.��6k���hN�F��Z��SKN`�����[ӕ��F��C�e�=v�������qQ� }ї�z��mgv���PF���
�JOrI�+��R<\m�L�<�`��8&��/�Zхs�B���s��]�[�FEV�
�~�ŝDP�Dy��F=��q8���.�j��Z8;�B����J�4���2�K��x��#I�MW����YfR���Z�(w?�(M�}�J�/t���#�R\D�������zqw��K	�`��\�Z�2���������!CI�<-�ٗM��ňg�4��X��ܪ���Ǟ�yUcD���@�?U;秌^ٽ�(�i���%ី�M�y��]�\�-��)Q��j�-�3i��&�M;�\ix�+�B)���76a�![}
�.V,�+���d�^3��&0�`��VP��pl����%�xv�~�'��?�wR/�T;���%z0��l��YP�HH���E�(!,sW�CΏ�,o��1]9����������A��Pʌ�����mH�__��Ut��源��.B�����N��4e�jh<Jd��G?[<BL�����~�.R��sJH��pe^_�R�qA��t�^[njd,���z����\�T�����OIO����l"G�l�� .Ռ|η f�:�.�Img\uIB{�������  25��v����g�}�uYޯ�Y�U����]N@��Wο-\��D���}d���e��j���<A�R-X�Q�s2��������f`����n�9@z�@,�r�����$BZI$2O�M�J�L�m�mu��wg��P�����������GP7�S��$�u�����r���������D�/E2��𣗐L��ȍ�	$�1�d�������[&UkR2>�e8 lV�"�2?�
E�β����52@��7�V$\�݉�F0����ɖWᗰ�������!�R����Qg�K�5�cKV|m�!J��N�f�?���@�<�C��-���S�Kj���2���&٥D����,��5�k�rN�f{����5Fw��i�����l�F~�u
�N������.�(����]�QD����C��!�g�����D���Z�g��".shq���T�8M�RG6~"��gM�n�o�U�9\�c��,呓�ӊ��v���  /�Xf�5�*P&P�^�n>�g�`�}�޹q�Z�Hȹ/�=�f��Њ-b�7��Df�
c
JB���S��Geζ;�����jN���]< ����Cq�����9�`H �ιu~�U���B��z~ �'F���q���۹�%�U����oNW��0�$/U����R/'Gi�~�
5�j\�/��;S�:B!ƴ3̠�ť,�R�凄|��KI'�o2��8�P�2W��WxF]�x#D���bx�d��S����Pu��vέ�%���ݺS�9!+�(�6V�c�;�M�+V8RC���Ml\���{� VF���!hN�j2'!Ő꬞Zq�������k��ǡzh��׫�%;����J�ӓ}�E�i�&��G.䉨�Ʀ֏ڲ�>|%/�BSMLq��@���R�\��ⲗG��a;����ݕN�,����`A��ޗy�[w�|� ��i�B��Ĉ4���߳ib^Z��b��j'�2��X���$�A,���,$C;�r1Γ�#1t���u1�w���+�b��N����:��#7��`d&�{�i-+^�)Z�:NWE�����z�,�.�8����=�y_��"��u�x&�G�d۔�eL�	��T��0>�(�"oQ2u�/���ھ�� %���^��iJ]�%����������4��8!�����uz�v��1t�%�JQM�-E�K��Y�p���]���I��0ь���$-oL���
O�ii�q]skܠ�s �;�VR�g!2Y���M�ڷ7^R����W���*�_83�qbV���%�n��zp��n�A��4�Fs���Y���x03�k����V�_��^w��Lz�}J�_xw�T*�����{���8��&�p_���#lM�$K�r�I�Ma�o�E����-^����>��͆�4�[/�(6��~"���Ϗ��yʚ{��	��@�h��������\v�ݒ �k�`����R��N��O���N�F��Y�ӝu���Ǩ�w\���SY ��)��"+�eSZ�dz�,�V�ŏ��ۥ�뵷QԪ�M�A1(�g/41�n�!���T-�DD��t�*�������h��Ź��ˡ<�vV�RS1P������S.Dy!>�IX�ѱ�����o^��h�M,���8������+J�
:V<Zs��N!'f�p�k�����3wq����쩌�����ڞ�,hA���S�'E>S�O>8jo��z$t̸xZ����b�ϥ��m�y笞�R0?3���u����.�� ):ݶ����,���!���j�9u�"H�,P�BE�����8�,���]]�~��FP�)P4��Ţo<����iIO>J$��)��S�i����C�)&q2��f�>�$���]����/#�b�����os��,(�mA�#\�2��:�Z #NN=���?����֏�\���<?M��)#���=j�bzvUX+?��ն�w�?P�LId-�$wb��T�Ϝ�j_�G\��F�c���(7=�S��YseFtoZ�^������.�95�x�2c���x����#5T�6���܀�bv�&�O1���잻��-��ֽl��W��Q`�Q�*�������|��m��Nz'}�J�����8.���;>�v}g���كl�)A:�쭵:?����br{��zjp+�۔F���rHz�2��O��Vʝ��r%��fy����ۜ�)�b��@�#�G��b
Q�S�٪��1׳�J<��x�p��ۈ��t ��u�9����07ȦM��l%#&BJ��qՊb��'�\��>�Ė��.'+)���(V�]k��6߽G��;!*EK?NŞ�3�o�����Ř�Wq&��9�:���~/=�8�,B��^n�IƴGXὅD���x�W��% �<l� �R�b�ś���"�%V��\�4�����d�ҹ{ >�@C0&���y5��О=�m��l�j0��Mc�C�s���i�m��J�YI��qO��	�K�z�B��|���Tز�"]nO�o��1o���%�l��Z�{]��*�H��ra(?|8�Fx���x��
�x\����7�l��!���� \���rĻ�
��_�ې��� i��..��{�]�
4ZZ�S�5���tZ��H�v��`���J�D�#�yH�N
M�)I|�� )^���QMw�;��������.�㉓���!xPLu���C���)6�y����%���
g���w\�ݤ7�Pݱ��]I	��Zh�څȦ�Q��֦n]?ϧ�bDe��tA������`8���T�Y�Ը�t�n�.T4��'?�q$����dp��$��L���ǃUh9G�(WqJwd��y��o=[f�D'n���/n�3�K���>�bX����%��J�y��pE�ts&x���­y��A�"fa����&f�F�8��0���gIF��p�+P��t���8]{��|@��s��]]4�j4���� HƯڶ6��7z�8�� J0@p����r����Z]�yݬ3�Z#�f+�LU�b
y��$�uJ���|�zL��կ%��&��@��Df��E<�	+���b��ɹ1��
�o)��l�����'�jJ�:��W�m���rDO�D�H�E* צҒ�a%-�l��U.������W�K`�ս�Ψ�P�����a��~\A�I�B"�C� _P��=��H�����4�k����څ���D���"j�ߛ�̍�������B&aL�շnQբ��S�%�L���0�v��W��	�j�
�LA�������PCw��/;�9������ᤥUh�5S���VH���s<�.���T����d�S�����r���,�9�	�ȡq_I�L��8���-UC�%�:���G�o�_0�ҥ��Y�W���ۛ��$/@�9��`���ȯ�/�)��}�\z�T�]nG|��FA���o�i{H�¤��
$�8b5'�n_�9P	�y���v�0T�IZ0G,�Mn7��VoYm̷�H��,v����=���%��t,�	�S�񵤋,�������9��g��׳��R���]5�@ǣ�j�]ʚ���8����U�m;'��*�o�hYY�%��g�V�Zc����AY^v?5��7
���1����@����/5���kW�#Z�ΉG��H��QO�k�v8��W}|eeN�jԴ�v���Pǵ�(v� y���4Yw
��V���,G_�ѱ��)�����ّ�b�����9TkT|��`���`Fb��Mw��o�@ER����Kp�����QHB���Lm��$��S�y���gcD��/N3	�'ʆ�`��2�]A$ �ĩi�t�v_��))!�g���z����C�彼���#��P�����c�Ƥ+*
(�O��T��O��6�u�3��Ez�������R�3������r��yx�t�A�c���ڏ��V�A�s�r�AƘW-Y%g���EQƲVZ:����t����j�[���h+E�|��Tà,f8t�/j�<�㐧^l��]6[^�]�e�D�kUC�e��/X��<.3��G���A5��>ʑ�pR=���-��ɳ+h5��&ydd�=�ߑ���]�FO���2�3|kؿn<��{4��Wǃk���Co\(_�_cyC Q�[�_����9�|#1�Enm��
1�rǿC3u&r.�I/D�X�?�>��*�D�z�ay�_��o]�܌P�����ӗ�V��߯!H��;���&�T�ì�1�Z��t�����zKb:��Ĥ��m�5���ŏ��T-����!q����~��ߩ]
Xo /����Q���_敛���7ג��T�bRF�rSF)5�=�<�G��|(�b�:p���`�ȏ�?��@*��HM�t�/�����%�p�kI/˖�[�f�m��C�Wp�rv�� �l<L�����8R��-�N��WO)� ܴ�EI�5JB(�.��#����g���e찎*v��	�
��{7�9�� /��]�Y�_����!Hv�l�C�iUi�BoH��|�0�u3���q�	n��F�v�Z�:�5a�{Ʃf�f'e�XY��P�D��FDW�R������|��-��2�av~��;�O��OytoΗ�o�,UE��09���K���jl���ڿ]cmz陚-�φL`O���}��Wi�j���݊�2b��;yCj�5&�Xu�U�iZ�0�Z���r��@X<c���>AE��G�5ލ1T��f,
4�g'L)� K$ln�w���@�e��(�[�}<�X3W���";�n��$��k���מ�^Q��ЇQ_�A��>��d�{bq�cؓ���S>ε=� �0���(!|ώ�JZ�D]�{mPP)�H����v7:TME�QG��9b�Ť���X�3a��ߧ�?��ƓX6����Ů�m��٧_Jk�Z�Sf�T#~��$T�! ���T�C�$�J���C��/r�~���~G.ڿ�2�lC�(v��r�4��B�٥�Yb�Ĩs�{q�;md\�i�<r���Z�ĩ��C�5Q�"�Kh}��T��:0?�<S��ܸ�&����k�H5\���ˑ���cb��XY����;�C��j�A=��8ң'����!�^��Bzs�� t\M��+�'ﳗ��7p��;$Ȃ�U�g<ڿ��Y�WPn��Ry�Ґ	�z��6�܁�ocC#���/��M����X�@R�vU���e���ꕛB����h��C��9�#���Z V���7�,��<&D��,
2�o�H��ҙ�XE>*�v�z��i�@P9w��(���7yO��T<���r�1fP�-�):"�Mcה�̶��Ş������Ώ	4��Q��i�x�����:Θ�Op�p��&P�ᰲ�=Wp	��f�PkP#89�0�	�nR=�y�A���1�q֊�0���y�o���:X'�����y�N����p71��L������Ί=��J\�CO���H��.�Ҷ�g�騝1 y�3 ���Y��Й'K�������>�:>���;��7�V�&Oqݽ�����$��d�镗�\ܴT�8��<���22�{SG��]���JE�5����|\���m
�f��iS��Z�LZ����+�v����L���xof�P��t?�7�Aك<�[�ܰ���׆p���j�_5v���������W�D	z�;��zX=wp����.sS8�b�s,�,[�Hf�}x�'�'�/atQ�}$�oy+����ˋj``�i�}binR��/����w�Z4cFகnb��B�
o x��}y��l�P�5��7����J��xrDe�����T)�>�90{>n���Ԕ��A��J����8��ք�ma���J  �q�c��3��9'֩�Y(�x�����׶ҡ�e?^��3<i�>
D*N�,��W[F}������*���|�E��|s�yGF�{Z�_�O^�<����W����;(s$���Pm޿�G�#$�*1��`C�t��Ơ*���=)��<��=_;g���4��o��Pɺ���z�V0�:<i����8���X��%k�`vE�)`T�_Y�>��WY/3%;�:��'
�V3��;ӷI�ݻ"Қ里��M��a�B<����'�%�PS��m'v'��"i1�#KI��E]��� [Hդ"|"UN�l�az�'��2�`�g4��|��X�z6�ݎ����A�WF���י�-�͹��
��`C�"�S�@]:�=(y�Z��4�����>K����5}Z5Xs5�W�cs�g[��G�u�����K�r���z�)��6&N	w��|���B���%+�z��� ߀ӧ{�k@������m��ոg��s���
'�ñjP���Î$C�_4��'Kk��^b�%��!���m�鿌�S��Tt���� �����h[T�� U�D2�$D�8	!1E�THƦ�u�>u��{��6'���s��`��S�]�r��
���j?'f:�bl&KKY���e�j������1aE0<|�j�,r�\^B�N��һ�����V����9���k:c���؞tyV$�?]zs�Y�k�-�5W6Q<_z�Y&b�;��Me���ɺ�_7&����OA�gیL�-��t,��7=�e��)�6r�@�	�y��L��M'�� etՔɤ��D��x�۟r�,עy������A�|��x:_���T:@�zU��(ď��,p>��J��ٝn��j��L4�Z����el��F��n>	��G�-ݚafL�M�A��]M���8�]�K��Nf~�,���w���G�yc���!o͹V�k���	?c��d�*�X��$0�������.`醊
%��f�.pn���:����/h�D�#3l�}����j������n����h0n���#��\(�؈g8<Ծ��U�bipQ�4�"���Km������+*sw%
y�����EV>P��ϥ��y;��Let˘���?S�B8�`^�	Mdxd�	Uf�$Du�4���$w�w��"�Dkȧf�T:��`��, �!����.���JiF�:`���z^G��;�<pX�yN����dS���k�ت��`�I�t�	T��1�Z���䞝��b�d�;`�Y���ʬE��|�k%(�Dc�,U��gN[��z�9�\
d�R-���io�g%z۳L�I��o �*�g��:�6w]�����G������k[[�H2����i�R]u_����9-A�O�$Q��4���J����a+��2�dV���a,}�t�uHq̼����X�ԉ��=EF ����>�	�~U���ݽѱZt�F������}ě�l{�ɰBrg�s�]f�,5!�C�^6�[s�d>������9���ƌ�]�*�.�+4�0���o��N� �����ZTA��n��O<��&b�ᑉ0�?��n_��)5���Xve>�@��Of2�o�͝�˓F��;�M�f�S���V�ȑ��Z����س����u��(i:x��R4�?�q��쮄�׮ �o9~����Ĭ�P�-�߬J����3��:��ݸ0p���6�\3�o��Ө-���\(.O였����q?&����we�V���c	%\gm�|V.��5#���. P��Ř#�7b>ç��r�Gf�q+LJq���@V�+�Xx&֟��9^�R)a�$.<�m��d��E�
ĺ*�$��ho��|���D:S
�a_fC])�2�����mP���*�
�]��MdG���<�-��%�����+��W�Raa@�oy�h|��˲�a���K�q+Y�#���(4�ٗ��$�J��k^���4�:��c-�o^DOl1F+��˷�Co�vGm&��FB�F�w����%*c���*�叁s�⚳�x��R�GIE���F�� �h�A^P�����vE�7d�) �%>L���9�>t�	�d��~r*vǘ�2�K��?��яL����S�cی�6��~���@5U6�������w�1�'��/=U�+ZC��yYWg!0�Q�"/	�>�t�㈱����ɾŉڌ�<ٚ&^�|huė��Na�At�N�L7e,�T����͊A�{k��ѷ����>�q�������Ey�Z3�bzX6�/\|u�RQT�?� eժ�>��7�7�M��\"���]��{���״lp)r��Ɖ0�j�5$|�t�@��&\�;=���0�����"�h�0�ٜxﳷd(���>36
�pM͹: ���.����QS�S4z$����C3��2<�;�k�
lw�r �߹&�6��L& �8`�@΃%���,bQ��wCy� dDV��V�}���oT�{DA��ɵ �<�1F�c,�#@ά�"�'Gk�^��?@9��z	D��>+79M���?#X90�|}���>�:�	{�
	�F�Vn��Y_u�P?~����O�,�&�E��&^���,�ɘh��`=���n΄֑�e����{�oY� ����	ی�u�,J|��M�s�T�6�Z �0���I�b�1�m�(�Л�]��)�إ�8��� �s�_@���A̓d@#������UF;YL/n���P�]��P� �s�&�B6��w�<�=<$W����s�/h"](	w�����S����ot����g����v���MԩY�?7���y��s���@��4���U��u�%KN���T����Z��[G�o9���B)�&fX��Zd&5 ��Vk��)�XO0� �|�-��}<�t��̈��ܨmR���f=c3�������!��AE��M%��ͻ�j��{�������	���T
	z��	��T��s�!ǹˇ�;���L�us��<X��F��8�4Yz��)j�t�~�%!����\�F�2�/�=����/�U� .n5q��'�.6]��槩�YvQj����߷������PV��i�T�I�B��"@jġNyj�כ�z�a6O�MG�r�����&{�R��Qq��;�Kݍ��V����}T�d۶�"��ެ���}��O�N�6_*�����;y��|f����ЀSw�5n���=^�,�'f��7�kۦ!MeD�3�``nX��Ӯ�R_�(�|:8�u@3����.�g�t�W�w�]�m�7^�\�W��E�Jrf�� �g����X���� ��tFs�7Z<r��{Y���f�i����o��S���	���Cz�js#n��ƛ@�����ax������M��:��eJ0O�{K�?�g�\Hλc�,��[�����Q��Q�1�J�����=u��;Rda�PP�1����ҖY�R��ok��z�{��A�f��;��B�K	G���}��Ñ�h�Y�W�gml�����Q�$72N��D�v�U6;�QBUWw'����qz$[�)�k�@�o�5�Xy�4���1��:bP�I��JN�������Ƿ�K�Hx�4��܁��Z��4!䁲�iO��?��ӊ����ߘ���Εk%tO2Xܱf	5[k�ν���TjU�vW�����q��w6�ᰌ*h�����I?.$ nH+7�f@���F�W��aߜa ���Z��	Be�S��O|J:M�gz:�D>R����(�2�o_���`� �)aŎ����3ɳM'�/�UB%�'H}�Յ�:�jM��[X����c�?�E�G��P4��y��B/EP��l�N�r�<�Gu�S��~5Ԥ��?��������ǖ��|�ӷEH3oS�9
�h�q�i$N�(d`�
������xn����L�!l�c6�R�L*Un�l@��/���G� ��W&M�2�n.L��+�HWO������� �~�j!��5�����b^�R��^�Xr{,�O4�E���ڠ��A��a+��e�Gt��o4�Gt��t���T��jhS�M���a�w�DR>G��J�2�Xc%��1N�(G�ѡ�J�/�xh�_u\W��8^��'i�hx��K��s�!�K����Ns�wj��A78Ĵ/t��L�76M_�ї�F�iq��j�;cX����O�kI�b�$ m��bQ��d�ߪf�C�	'��.�R8����C���OY�rcy�Pu嚗� ^��L��G��6u۪Ϭ���%�8�h�����9d���pԯ%�{���R�-�~N��i׻0���<��k]2p�H���l
�_mT0��X�GW���`P���BF�2�l�w���x�2��a��e��͆�,�+�5=.����sT����ba�eYOHp��z]{�&�$͇*�$�	�Ta5N�=�z9:�́��ȼ3���8�p��R/J{|�\|�3ײW2��v?��˞Vp���&�*O�,�V�� u|twDi�d>T�`�W�Q�h�dg��ND�G$���x�six5�X�N�G�ae=mc]GZs����e<:t!�s"���.�}Xnt*���]!*�y��[YO�:H%�M#��� �1�Uʏj�<<�c*�����^�C�4�v����:�%���������Z��ou�M�����I�9Z��e�ڐ����2���Z��E���!�C����$ �grx�:N�Db
eZoT�L���m/�e�Tx"��H�U�[�V�8��g���ؕ�c��#��:�e1`����r3�Sq�^��˯;
2WA��1�����L��M�[�� �jǢj�?���S��w�Ek��k��a��p����Lt��C3����7��0��	��W�$M�c�:��+���?�˕������Pp;��Y\-8����﹥�3e&{��H';�p�Q4�y�3��!�RM�l����n�O~3
��-��y2�h���/�&`|Il{�F�k"��O ]:i����N����VKO/�m��+�>�k��V��Ĉ{�-*��W	��4�N��5��f1���R�S:��J�7>+��6�wC����uu��%ҳ��ɜ
��r��]���b�I�?y�0v1��/�H;�j?$)�S��c0�`c��0�UU����k�z�C��R��Wib�P`��b�����>�*�n��ݵi�q�<��������]+��O��%`��}�WC�	��&ł�.�����QsT�����E���Q�|�[�jS$�4F���8�P�B�?I�q�'qpf�u>I���w~��?醑��V=U5�N����s�!FY���?��Q�KK��cN�Y	W��1SR�)y�V��~C3�LC����q�<N�`t���Ʀp4��E� ���Uuw�_��E���=�9d���~�Sit� �����!���e��B����=ΰ!��A�kn�.-U����7h�Q�
��-ڈ�V��s�H��5/I$��zuY�G��U��cB %�с���I�#G�0roQkV�HH>8ϺG,.W��w����9:ú���չ�!!�L����}hW��7\�ĐWF��ĀS< o4�O#,��=-��u8��4�ǫ��)od�2j���޺Y_��>xҋo?�c�,�������N������Γ/L���AD��	�̐��S?��PB�FH:��8�	P��}�E�)=h![Oޟ��}�Ϡt��K���&i?g��"�_���w�oUyH! a�i/��#����Z}G�OA�����wɌv�W˟�}ȯu�JH�9`���U��c�6�n�H��sj�]�ax�hI���{�%T�6��F#��Q�NX�G�f@Z���H=Y4"���9F�~;D6C+�(T���$���v���:e�֝o�J�ގ�눴 �\_�p\3FE�;���*�g8�[{�ʯ�s�J�a5�1P�qQ��7
&A�-���U��]�� CZ��A.��v�SKro��a�HSЏS�뛹򮪕ޚB�;v\�P���c��� Y\[(��31�џ���d��>`�bӏ+V���I�,��ByI���
.=��ֶ
���{l�R��yr��2���_
$�����[��W��1(c��=�Nd��oV߬�'�>{�.61��(j�;�<LV�
p�� �v��J(�I���,�������&]D+��o"����MN�Ye��;�m�:���4�P���[��gȶ�"���}*yWY��QX.�#� �[���9��c��l-�5W�7_�#۪=��R��љg)��V�ŁmpB�#ٳx �*;FT�5u�^�m�9g��cP�˺�7ze�r �����:�b����y��I�P+}_\�gQc3��Q��Uk%=�P���<x1r����:���"�
�kF�.	�kâ�P����C_�aݿ�ΰ��H>4����e �7�ł����}�S�'R���-e��[ ��s��_�b�gc�p&N���rp��PШ+�Ф�f ߚc��v{"Y�KHY��K.wd�v�Cf�&�q�����5�%b7q����(�f_kX&�F� `��A����t��D��4ܝ�45�5�ܶ/��D�2�w%�j��h��M��t�d�p���"��b����>��V��<q�	���L��43���ao2O��V+T�����d�M�Z_�Kq7g���^��� 2y>�G��b׈ �*#��*��B%H{����c�c@��K�|��l`��m�P����}�Id7:']ͤ~�Ω{��kP0l0���үмp�#��W��3 �o���hG���"��S�	1�`�]�-�@T�N�Fn�8e�R ���C�~���GT���A����R0��Q��s��W]O��;�P��j?�Ȭ�_"����S���70-Q{�/Z+Sf��Ѭ��Wz5�;
���[f~��{����TL/�����gz��f_��%
�+��Bɰ��,��g�
�׍�O�����O�=��$���1���O]8H
�h�~ՙ�u�	u�N����ǚT�ߨ�\Z�P���"��^b�
4^���FuE��(���n�P� �Bl�lbK��}e�CV��ۙo'�=�<^֋U�*�>��L·�x���̛�����N�-FUé�\�3A��%s	4"Q�o�t�:��N[T_�a�Z�}��AZ@k�6A���۪L>f���%R��:��6\��&�׉�G�{����>��+�
�É1�����*��qG�FE,�L{ !A����,]&,�|=�s$���j�1��rB�\"f?Rv/ �-�c;��߱;�5��s�CU���D3���tP��H��*�܃�L�肩��5JI�M���baۅ� ���F��J�.��P�|�	>y�Z���:�b��.�$����������O�%6�7/N�a_��zo�z�q�"F:I����� B�� �L���'�Jcģ�9���h��#��&�J���^�ǔ��3#��*�� �A�ĝ�N���]�th=i�b:�����T@	���������+e��ߘ�������MU��34q9�����N��Abs� 5�lI���'Sڟ��zȡ�2�G�m�I�irs;bj���>;:�����U�9�S�!Q����f�AZͼQ��������{��Ţ_������J�[N��`V�( ���j���z~���\	��܄��ʯ�|j���5���|�ͪ��N�8�;�Y�6%��y<�L�_F���@�ђ
¤�:�E���)��� ?&�"�H��r��U݈lcwY�a�9�ڷ��SC�/�g6��&_sr{�%�����[��H5~��qC	Fa4����Cw>>j� Y�`����k�A�v�F���/ll:��j�#���Ӹ��	�A�'z[Ŵ�P�t]�L�E_�d�g1&�Y8VU'������UH��&���R\l�����mS������#�ܺ.�����k22�0�&bW6�t;@���E�bG8�&���n�%oR�tSV����~�3Og ���!�[�݀�s9��	���.���'6g�5 #!�:�#3ŧ�L��5VApOz�N���s&?��陊y��RSL5��~~���{9t�w�����9�� ���B~,}��� 3L���kW�JHo��� g.f׳����X�z�1!Q�Z��d�$���+;�}$�R螼���&U�gȔ�(V��~�#�y���ܤ��T�!L�-��z�V�$��V���6�*^�A��7���L�*Q����������a�<��~Y�4�5�J��_�\燸vJ�
�"F����u�T�|L�G����Jf�W1�2�W5�ˍ�*$چ���՗B%�;�xȽ�{��灀.�L�c��QD��u~���0�������(؋�����dd�U���ק�.0<��l�h*�K敻Z�-�5��<��j̇.�;k*1�߈x��������;�j
�C����-��WNR��T%��>�d�GK[�p`Q53BstEWb`�����FL����]�ԃ�{0���(��6F���ܮ-{�b�խ�&鴕U|aPSk���J�W:�zCD+���T��9mT�K+��|R��v�5e#?�%Ra�V��;��W�X��q��",&u��a�`b3c�{1D�:OII����C�JӚ��<KU��u��Sq�(�J�S8��v��������L�4�X}�&����DJ-C�Ȅ��v�.(���+���>t�؈Q����ǜbק^���� �Cd玀�L`ՁO>���
#����䅐�Xa>����Q��f��ߙU"I�y�H���OQ�]�:}Lo9�wgS��1��.Ҿ.�����(Z��4YM����'$�j�t?P�*[�;�N�6�T.b���}a&�je�&ɍ�E^o%�pK�V��Z��6�E��q�˲�zN�������Ӏ�������vG�ʮ���a�#A��i.B,?�Gu2Ff�� ���| t �z~)��^ծ�%�b����Y���}��jܝ��	�6�_�� v,�mn�J
��q�����=�.�,}Vv��-)R��[��3耘D�8'��cq�'�RD��X���^S���$>6���cr�w�/�\"S^T��ݸ��z����U��_�+�uS$��$JL �iRqxM�]����9�^ݩ�]~(o����w��׷����s��b���yDI�4L�(�f9޲9-�e}�8��11��[q7&��ǅv��Iw�!Ě���i�Ѓh�{��5o�Aj��ձW
70���E"��fn�����@y�6���	Unٽ�z&�GM�[�TO
�|�JK�3�ЯF��}�&7���s�� 5���r"X/�
+N��܏�g[�De���D�"ܫ���@# ��-�n3m�.�ؙDuB�>�$/�F=dԎ
�B�x+��j-��3{\�p��<�E�����zܤ���[�Q� �VK��֋�����ek
}����cL3�
�;U�v�(�[vx����+А�!/ѳ4�>��f�>ތ��_~�_��BW#ʿ�~�_�O�sS[Z�ӺǞ�?��\�'e�n��d ���5�u�M]s��QܧinR~jZ\k7��'�9 !u�J2TT����D�
ߪ�2��i�r��]e$��՚�P淴;�@��cH|�kN:�	r7�I��z�`Z�N�Ö���"�Q��#X��//��ᑉs�!��2B�2r��:�	�:\�;R���,	_����5�
:9�}%��O�Q�o��r���L��]~��l�t&l8�*Y����\F�[f��_�E�%�f��0�M/�I����V8v��-כkIjS�I���V�M��=�����yr�"�DA��Vv�Kue�5��h�,�EO �0���}���jٴ7TZ*2�&������)��^���*�T���w���J��A��9��@���vh����DLG�*��:�6�Іeޝ���o����!٨CJ7��&�dX��?�y�4�A��;�ԅ�T0��dq/IX�o�������J_)���S5�����W����^#77m��R���߂���%���B�L�Ch-��h�N�ٌ�p���O�+K���??b�O[��%�W�J���&t������'���	j���������؃��N�c�?]��{Ç�D^fǐp�����+�6��Kmp#�Ə8��*�d������R�7�mMI������\r"}���q�UZYr�g�t6���9&Sŏ�ߩ=��u?ǧ�����7��߃u^�y���H�������a44e	.$b��	��UJ���_CN��`CFD�cC�2��	�F����`��\���(٬���s��V��d��̛��Ynڙx�z���a�'S��7\����r9�ۦ}ޓ�f���$�H��K�r���l}�;�#c�1��]�77#5�Nf��"*�Y�ˇ��e�0�,�	TCѷ��������&��>Z~�?]cb�j'��65�kT�E�^gC�n<��V�M�:��l¼o�u��k��wV����";gf�-P�Vꌛ+Y{���s�"�(87�F��N@��cy^[���@p�#پi�!����j�<����R0.`�;5.	aY�u^�լ��I����զt+�f�9S���'ҹY��i`.�S D�AN��$'���6pL�b3M�c��lh�G�1�������.��_<�Z�s���z����߸��t��s6՚شt���16e��nE�ʲTB\V����&q����?�g	���@Kp	��I�kVh�L�����S����KX�V`����dڅ�)�<��~�#�3��;��¾	aU0J�8�{��]C��-�sO5�:����>��1��8�<{�D��V���E�Ƹ6�C�Vv�n�!�����l�8�j��c��ԫ[}�h��� �-?�54a��"d�����������ktl����������E�x
{C�Δx���6��˗:�A���ڟ��\��r����Sz���9�[��9�2mu
�͛��&�R2�ʬ�{�%?�̤R� ~�7&3����쥦�����&>���ւV��"ˀ��q��������l?��z+�P�� �=��~C�fz����S�T��]U)���'��0�����ݲ�LE&YU��۴���"v�u��Y.*�d�Od�@ H���;b%O�#C��4)�'n$�HS�[v��N*W

����x@ͼ779H�����,b���T��!h8h׳kE��mF�k^'3�,�Z��X�&��d�<ꔚ� ̺u��a�?4�˦�?�L��0kl�#�Y=T����Y詠T�m�$�f�t�6ݯ�e����2��n��&���r�ی�$y�
��+�mZ���������ܪu9���^~?l�N))p��K���_wy��@�d!�E@=K���s1jC�� ���+��[�S�_�j���g��̇�3���3�~$�La޽~]�FV��}��W;�RYg��o�$������C�ϙ��/�=
��n	���p���SU��A�E
���'�A�o�F�T�l��7EG��M ���gU(�K�	�DgU� {$Vicn#A@����=i���%���X�''��:V)7�'
�@Ax�r%��(|����;���6�X�����J�Y�x�"�r]��}�KV,"8jdAX��I(�n�_�X�я̞^�w�Rz�����|�]����̀���}X/��Z�������ng�$���>�Ƞ/ߚ����d'�H2w�V��*>x�x��W���(�P!Y��5���aD�����f*��L~ҥ�2�
ns��x�|��C�*�����s��`��Ó>b�佑&����3����6��]e(A�`��� ��{!�s�-�`�jPx�TFT
��c����y���4h��9�l��{��ޝP���T����J������d
�������[\�S�aPch����S0~&j��Z���*T�P��<u���?��&9E){��n9�L�����@Q�gWtk;-a�4��:ip���{�K^�ZuWr������v_�Ц.�h��;Zז�~ͧ����Q���|���z �
��z9��,XnI�7�*�K��Y@�Q=�s]*',�{[�v�n�CO�z�^�c��j�8�6�橙��L8��֢��M{?SɃ�� ����	ӹ���n��ɇ� ����D<|J�"�|��F+!���kE�X��f�,��*�)'ƴ{r�D`��;Չ��'f�
u+��n��/�VA�*Ie����d�G��#Bu5��p��cvH-�֚��%nd�ca�K��<��|-�V���z,�v-܍�
�P@��.R�f�.D�m(���w���Ĩc~�}���dסQf9(�� ��'X�;z7�W��[?He�/@˾�n4����~�2o�̻i���T2B�d��Ԙ��E�5"R[��:xihZo����#������1)�P���b����K ��Mh"\�A3;[K�TT�é�7:#&?tY�yQ��T�&��^��P̙�Wpn+ �C"1<W�z���=�q��_��4F����R�蠦֞��Z�C�[Oh
F���_`��=T4zk�w��4�#b���#�+ ���+��uk��VM��=(f^�lv��ʾ�_���T=yiVZ��H��� �.UP���<Ȉ�].EƳ�U�ez�mU���-iՈ�o�K �._s9��x2���d�\f�،��.����{N��ry��8���KArn¯T=���I2�|�{�ӌ�(��vU[ǡ)1�^��(��a�2O$p��g�L.�	�[�g�g3v���2UĆD�>�l��:������QxA9�iӮQi5�/�����h祕i�M�I+�M��F��?<h��=|��8����Z�k�-���������|JS���[���=������gIqm��&aM+�����y���X<- ��&���TBs!�_� Z��J=�O���?���Б؜�t�� 鵨��(ͧ�Ăʤ~�����d�Uj+���SSh��i.eF��/�;6��u�f�Q�+�����ǧ _(���/o��<�+S0�S�E����!�Zj��2;�U�郌��F5hB����4BP݅����~,B�*GƔ�Z���F�8��7H�쬼��������W#F���~��/�\|���v���]���p�c7�4�DSd1R����"[���C;YNzYڻR������~R��m7��kTN;c"��7�������/!���^I���1n0�9�	�x�����
���+����7e�m.�p�a��cVe���/��k���'$�ñ>M�P!���'b-6$ɸ:UV�l�Q�&�9���k������ٌX��qPbF��@H�)/+=�KcB��,4�,TrF�{w0�a�BR_?�<��[�����řx}/��賋;݌4|��\2tu��̗���[��g`f��&�e�JKXSuGF���۰�%�w�QRu'� ��tv�&�GGI�{~Q�n�_��e��Bx(�k�i��ͽ��%O��A	8���h�S���}�K8O*B)a���/��wA�W	22��5tSt��=��]�~���&��Y%��ӷ�L��R��u�<��]�g�-�Մ�F1�F�j7�������գ�Q�l���'�nN5��;�I�W��jǲr���1�>������y���e�ܨY��$U�e��}p�(jt����.9�c`��P睢6���F�������vR���
,EhZ��7;;��%3k[J�jC]���f{�5|��o����*Ч��y�0s��F.��xjk&~�v��(X,���,U�ywq�&���G���.�l}�7+o���%+��j�e���K��F��q�n���3 �Ѽ����5���#X5G2���H���tmoP�h�:6�%o�er���PC���(�0��m�����N2!�б�9�K��T�8v�EI��u����r� ^� #�Dv�u�u�k0�(���V$�����GL�ޏ~�<%���oI�G����::�>*̵��2؄���ߜ=�	�\�3=����5*���&7äՍ5&[p_
���_�i�<P줢�b =��c�@���`1A�QǏg�a+�;��ᛡ�� �*�O
�ެ"%�(E�6�����l]����eK�G�C�d����KRa������>�0�ivJ��FM%����>�`�wX)�~����Q�Y�ű�o|V�i6��S��ڠ�s�J�h���@x�a�n�5�p�Yk�+=�n�#7��L�EJ��\���j�����>������o$��؅�gj�����I��؊w��JX��	�[�p�2��M
2b�'׌��%�:8_k*Gz�f8çs���Hu$Pa's����Y���)���W s��徛��7ǔg~7��9��O�=B��5�r��;qR^c��~�����'Q��R��Y�w�gFn4�ۯZ2%9��f��dbVoh�-��c�bN�X��6�r��=$=G���p������?햮1�(Ϊ+��1�(�1��q5�4��n�H*��6ͨ�����n��m���-�̴�5���ͥ��~�L���@LČ8�D��.�i�Ě��Ojg�<sC��(pӑ��,"�`U2㬓��r�Jq���D8�̦���4i}|�=s�\�~��=k����:EhQ�K!�2�t�jv�'��I��t��������-p��B@�W�0j"��b��_���`�Z��Ԥu��#�:E1���c��?��CXȣ{�����y�a!s�����µ����ۻ5���M�5J�2�R��|BТ{��<�֘[�2�5~������z�����f���")�VVv$�c^=ĭu�Q��ʏ�KV䵙�ݚr.��	[��]��r.r�B���4L�� Q�6��ǐ��B��%�.�t�)K�.ڇ�[=��5�ה��6*������j�����}�5g�Q,�c8Ȥ"�;�\x�Φ�{��b~l����.�$��Y�|yf��z���5֡XP���2d,
��K<`��szfh?�׳p��Iv2.f=�1&��=Ü�
A����V?���8�J��>Rb	t�K�:��"����I�(Vs7���I�����)^�b�#YY�8ö�Tc"�_�n�KΚ�?���$�c�e���3C:"�F�v��1N���e�E�,�'�g<>��>�ƆE���:3<p��7s�L�ߠ��ӧ26���X��B��W�M�WL"W%'�0�=��~<�H�'�@��ԉ��h����g:=���D�y/�S8L$�b�X}�_0��h8��.%aa�}&E:��9�T��I�y����O;��pi�(y�?O�Qf)���c�ds��U��)�lmE�*#ؼ9�9�-��z>���d.MB�E�u��E���!�&�[wg���}�OS�:Mǋ9Q��5�d@T��Sa+&�X�~�h�m{�z�驯�C�I�f����D�Eq�X�u����:���c��V0������a�Y%@��*�
&	MtUH��]_�x���oC��o(?I�^(��&~��/���%[)]����`��R{�
BL4�{O��zɫ�D&:�]P,���K��yQ���}6�3����=m��Q���;��m3S=riMǯ�heͺlzfc��h��u����\v?���@��ʢ`!�4�	�%�pЁ��J�֏n���dr6MN#��y�M$�-����0��ˈx��$o����']Y����Z&�������}��X�hvƫ����p�ٸ�NY�0ݬ=,��I���pa���ݛ�h3^Y�s�ʛ��s��|�.z�_��>������$$#��O��Ȅ��c�+���������.��,6�K�:`d���]}t��"P�9��2��+��F��{M �΅J8�[�R=��)�ee^	�]�Rݒ�c����wa��L`�C��Z]u�_��fY4)�?O�e�j����v�,n�����R]}�i��E��wx_�ir��$��Kyofe:��������4
֫Yݪ�l���F��/����Y��4.��S�l*~5�.q)��
 s�S
���쏉-�@��T�m['�8��>� ����@E=��>��0#�BCN��9b����V���Mw'�
V_r�&�1�+�n�5�MZ�Rs�n��"��ܞ�oSR){m8��N��|V��&43078C��I�-������!�l����u?Ў��Vf]d�;;�,_�v8�t����A�0#y�� �߶n�~!Z�u�h�i�߁TªI�s��pw�	��ک� ��>���Յ�M��+<�	 Ld�*bO���R=d�yx���!��+b*�깆��Z�M�{\ٞ�uh����cX��V�ղ�6;-�U
�
�thؕǌ>�9����8�����Ȍ���}	^>`(�aB��I��i��/�#k�b��A�GHV���C��oj�Vy�D1��U�P`MM�F�l��Ԟ?��;��wk��o�j�L9���:�{���$�zZ��Q7w|}���)а���3N���S"�3��ˀb�+U�|��Z� ,h]1z��5b�Hwc{�^w��*;�T% @��Ή���ٰˈhU�O�r\x�']$C:�lf�BiY�~�Cn�ͱ	-M]����HC!��	4~���o@�@��)[|7o/2.݋��E��1U���V� �4��<2#Wf}��'��I6�o"�7u��<�����Q�P#��r�:[8Z�k�%��|$V�S��e�h�8q-܃���B 8�&4w.�́��.f!7��l̗�(%-q/,��	ؠ6�o�^ k!��	����s�E8R�p�����B��q~\�ǐ��Թ��#�%��w�76�SN_�M/`;(�k\o����+ G�;��-���-��ꭻO)��Mڤ�aJߋ���1?)�!L�ڗO�s��b�d�j J�����%��CB�R��~{��v���0E+�￙����c��B25>�;��DOV�ڈ�O��h��03�Dg%w���)���}�����J��ת*�/�������{��9���.��[� P����s+���t�2�7�fͻHE׉�uƀ�L�r��
7'��!ʭ�)QyT]��1�Au?�� !�z$n҆=f �mB��]-\e��B����eh�L'{*�u�K�չ�o�t�J��S�H+W�O�C��%h�\Z�?��v[_��T
P[���K?Zl�y�a��n�Һ�����zJ"տM���}�7�~�jrZg��U�g��:3:�U󸥕����e�\�l�n�lA�u�C`�¾Z��㽰������Vq`Z
���қ��R�D�k[�A�^�]���3D��~��uG�L��>�E��;�z+x�v��� �u|1;iPXV�=���%w��1�G;N(p����2��p
���B2S/ʆu�q8�_(��;��k�v��u��>����#�,�шY�]����Y J��x����(����z�,�or�G&�w�!]Y�i��C�+�\u�?�7f�%J�7���+�$<�eҊœ|5j"���� �"������:/$A�?��U�M؈(����N���l�H�l>�R����]1v��e��q�E��2����^���p��v6�^7�N��/��t��g$��-����9�'	���2����DK�����'�T���Fr<���{�4:)�x�n�Xf�"�Wͭ׃$&t�*�����Pj2��Ǣ�/�:���H�1� O����J�c�L�C�V>�®��8ZuJ�o� �4oO� G��k*�@��Y��*Hn�w`d$�,!�oO�`�k����jJ�ɜb_A^C|K�'�4��5�l&8��������DD�.5���sV�pz8{�0�>T�pZ�>Z�*�?��J��6��E�G0}�?��,���l�-/���t�.2�=FV1~��u��/DሷDE��^�?M�$��ՋWE�H�k�O�b@���1��S�wj'�m^��h����(�K�kn�t��]��iI<�lb�����{z����:�8���vsKH�f��*�J��4��$c�o�~]~�	-qi�n��H�Xu�ֱ�J�'�sv��.�$�d�/F���A؊6��灠:���-{� �jw�C�ŮW���N���ӑ����O{����9����u�8���e��� }�B�o6&\лƦ��r���5FI����S����h���C�h��~�Pzɾ|>JN�f(<OA'��m�9O�[>�u�Y��7�0CG��k"�od�M�&j��-t,kX�C�v��#��Y���o�/��L���8(�\�  ,�q�{&���b,��d�#��-	���p���g��wkp��`�Ҹ�Ҹ5��c�By����Wb�cT�0#�UNF�O6T����Aas%c�(]	���g�*A�����F&�j��]�s�%�J�9�W
���om��c��6�P�ܱ���!v?,l�\[�k�[��Nݤ��ſ�UDP��r�zo,1Ha���Gs0`$�q���2��{�"Caّ֩LФ`#bCN�w�t����䜘�tGP���m]��>/�Ҭ�0w��j6c�E�`�(���/�Oڙb�\X��&�C���b��EP㞵˓�Y/��'Fy(J�|���i��%���������O��c�ۖW�>����^N��]��R.eEr4 p��ߊB�Y_�Y+]�^r��pU+�b˪��Jk�:��xIV-��G�~�V�L�\��:+�:<r�r5�!�Q�A#�jt���d��mŖ����)M��Vp �>B��g��TN�U�r*J���Cs+%	�kn�C�^�x�V6�+7c2s���h)acM@�4/8~of�u?Nڰ�gD0~��V�z>T���b$;E+�Ll6XR�g%YD71�/�0�=d�/aV�4���J�L@x�[E,}e�ia�]b���3�{lmg_�=�U{�@�#ik6�׊F�G���&�'��pR���h�d��+�!m�\�*9G3�3��Q��A����~��3��3g�US�L���ъ���WEs�!��Z�B�N�cfҾ_�B���������e�V���@�i�Va�{+�Rn�w�g��"���J�^R,�*��WjG?�V�3�v����b��R_G��O�����L����3��d�2��1x>j�O��1}��B� �aC2�Uб�߮������l`k�mK�*�5�W�=:��B�]I4�WR[�E��&������ g��e����	��8���e!2�]<=�Ȁ0�G�Y-�)C�q���z�������<գ���p+��>8j^�[j^8?�t��Z>��Pc�H�?��z<���������Q]1E�p�t�Q��+U���d���e�OɹjB����л��8R�$#������!qI�9��'�5!���c�nu���	�EF�.���Qۄ�}	�s.�`��8EՔA�[�f�H%'��Wn��&�"����sk��u��ɞ��{�9r$_q��ƀς�����$��+����ՅϠ�Pgՙ�C:�Z3k{W�D%MW/�Y8dXkto���X�Y'��}�<�J�m���fT8F�ފ1�V'�E�dM����S�����6O�Y~h���rdO�+Qؖ�TB3�����:=���͎����CٷP�A;�;%Ş}�dD�s�-Xn ��D6�l�8җA7γ��@��u6�@�{�Ppy���������{��&At�5�m��z�y�2J�`d~5:s*��h`�O	� ����5Ex�rԡ���C�|�Z�6�Ȏ����{v���($�ha����*��T~0O(RC�Fq��_[e����8�r��Ǣb�	T�e�s��8f�鐸�(`w��X@��-�պm/���Y�X���o�:���i�[��)�*uY��(�����)u���F��C�S�)PH��^Mm����.ˏ;SU��f�����X�1�$:o�7����C�S�jq�Ag��`	�'��Jv��Z���� b �K�3֋����(��q��D/H�{]�8��M �w]f���=6�M��vd/�LUP6�P��]��Z�R�$A=8��_��m�OM�g�	"�S�.��Ü�/�/����z�_�uLZBЈŲl�)7���,B�h���^����9p/�/�D�%�}� ��4�!��M��V�J�[5�ʾD�pt�)��G��b�X������bA �=0���[-��G]��-�Ϝ��1��Z�s�ǘ�[�����(���;5��:7�a�2;�����J}n%ڮi��Wt�Lq�el���L����R9IR��&+/ՏW�� X`�S��e%߆�$�	�BO\�s��Pq�Ј�L��É#{�{�V�e��}��([�_|�i8י-]�n�\]/7X�q��S��]t-/�S�Ր���E�>T���J�ͭ���qZ��q�^��V|���0�G�?���ʴ��{a��J7H:�W�_�D��-�_god	8`������ћ�-fņ��Xn2�������:�F����X�f\I�V�jQ��������9�Z*�����	�aD��(�R�M5�&Wڄ0���lԉg˼�>���fw�<���J���<��e�h�Hi���q�Ԁk��������q�{p-��C,��d������\U�zx��)�Bt��<��z�]�#�i��>VH&��ƫ�d��� F�2�EܱR�F�33ki[�+��O G%�gw�d�M�S=Z��Z%� ��oG�9�3����$D=��1�l1����!`�o^��x�I�Zy����h_�<�܆]);紷����5��vQ�-iE�xɠ�7�H
}�* �Y<�n�b9ɖ���*#��۷e���0��#L2ݟ�}Ĭ�:Xe��`x?T�yF0T\�V��/J�ۈ�]&g޵pn�=$����e�2�(r+̠�� �L�:g�ʋz~��9����&�?}J���%$���� �%k�t:&�z�;��D�BEJ݋L��{�y.��h���#�Xd]��$=�^�0bL>�G�$�_Do�s �>?3�g�fzwQf��n�(^�� aU�A���������o`[�]%	l���Oom�O��g��"lwn�n�J�AO�{T�w;(`�w�su�E�Q�%��O��n8 ��0�B�)��bW�c4B]x��4-�ٜ��ҵ����@�N��]�$0����eT>"(���!�$�y�}~rK'06���2��)�����aw��	��K�x<��P����
kl/E��[A�My��+Q0�d������'w
�޼���a}Ƭ]�����fa[�Px�"^aN�K��5����U�;|����#)�e�ɀ��a��
Wvq��a���+V���@f]U��<��ew����?f"��?x)<�Z�
�]��S7���_c�*�5�Q?���͌��G���޲�͠m_~`��e���,�F����
�`�d�Jܰ��%�u�O��ڑ�G��f�h�i���>&��@<��yM�b>�������������I��@wt)S�%ܴ�?��i����_Q�Bd�L��NW1���9��ް2��48���R���T2�l_�n��;w� җ�b��#�.̟q��6������7�\�.ٳg%l�,r�Ij:���/��jKp���NcJ<r��`B�儃ACc	b�g�\�	��""��@Ԓ��m�k����~쎁��M�oP=���%	�`��Q�*@�N��~d�x`�1�C�.��-FٰX�S�:��ٷ��R~*�f�iB_L�vw���O�C����JjR3�܊ �����p�O�0�'�q����HI�n��E�P�̍X�+te�fU1q�.�h/�F:ƥU:�<�>P1�O�K��vqڏ�!@��M+�a*��4.�J��3����@֋@�$��WS�D$0r�b�O��~3���'�G���PLE[ L���h�f�k�y2M��j�}oP6�0��˫O�y�y� :�7��\�	9�817R�����o�q�(�����}�(��t}�'��a�(]�GQ�Y�hh�Z�mB�
�y���q�X���s�������;���1��e[[�7�m���*��c�r&fٱ�Q�j,|�K��, �-+l�"���q�o�i)]@}�GY�b ���0�4(q]ȄNRS]/6~9)�;zYj��֪L�q���\;�1�����"d���~�;�5T�����뎒�(�g����dNzVo�M��(���j�	*߬_����%?AP3�O�i���)A�o��RwJ!_M�f��/˭T�J�=��r����3Tr�-�O�V�b
����m,-h> ��Jj���u����"��X"j�K8��g�B�93e΀��U:�5a>yjrQ��
��A�������V���6�D��<Z�/حk�	a�XѠڱB��uXsD�pz��5R~M+K��1$���{I����}YgR×L���V�3�ѣ�e�����)����n"�x���mh|�%�G�w�
	�S6#@c�Y�.d3�PN�Eцi�N�'-ˤ���A�Y�l�p(v��rO����"i[�|��p	�g�g�ު��.�h8�d�I�CwzN!~x����b�6�
��Q!������V�����̃%��,�����
L�%[���)TN��.���Uj��&��E:䢬��)�]L��r���.���u'�,6�p�8����\���\��qqyN5�:#����5	�rmGJgV�����?�E�s#�����Fc�0<�=��n)��ku� �E>�,��cT�5�E[�p����=�N2�RHn�_J����>M&*����F�賠k:�DT���+C��`�H{f�F��5sF����L�$Q�ɜW���&��45!зQ����Ҵ_��q�zSߺ�`J����,�}��\R�8�ܺ�|�:nN��2�os�	Ӯ'[W��t?�/�*f����Y	Gx�z-��B��8do �F��gC��Û~pwZ�j���4؄���.���Z$���n,tzδ��+����SA��gR���jb��B�B�6�(q��%8g�b���O����*8C���3ͨ�'�en�������b6 ��@ZX͋k�#
|3Z�7�W�{���.� ��j�ߠܯ�S����"��9�f;�͙��za��GY�x8z*���vl=�h���ߎ���d�����v��Z����V�q���3!�r-쁺8~����C�it6��_́p�ըQb���0��<��5E�.	q���k}���`�3I�ߐ�A���K�����*��)wX�������K�l����6��O Ѣw�P�t���"�����\���E3Ӳ�e�0�
��Q����D��+z��PiG��]wt_O>a!��x{�)=6D���E�����t��i����O��AX�#�9�󼰥��%�D��@�Kx�A�z���Ю�>ۮ� �`���xx�Mf�ːkǢ'T��gb	�s���T�+}�'q�b�T#x]S���
#�S� �:�z���m�3N@��#��xt [���Y�6�0���B��po�B2�7\���G�* L���N��8��o ��ڊ�1KX�����O��B�3�p4���,9�@0@��]	n+\�4�$��/�d�=�Ԇ6�����J�ph���"ޙ�a~�ߗ&���,�b�x�@ �$�$�ɑa�cM��s��Ճ0_��q��;�hNDtr���xi��PSAK΁l�TV����'�y�D5�b�E�n��Q��Ҽ�YfB��MeVM��O�{��͵U�!�)�5���Q~���zG�_�͒wȏ�/��'U����do�-i�*��������z�^���t����������ռ[Ip��G�4n,�$�>r�q �G\6`yh"!9Ւ�M�����������7�e�~6��X/<9̒� Jq�ZL�JV�+q]E���:PPO��Y�I�12l���薐.t�&�n.�yQj�ƛk��Nf~��V_͉��!s��p����GK�>��2b����l�Bp�Ξ =�ի��H�v}E;�ʠ�z��F1�}'q1�l���a��~1q���Jl�,�~h�/'���"����*NF�L�*��7��_.��0��1X1��!����Ev�3+��Qi�q��\Aos�W�|���A��p�:^��V�ۘ����1��;��&;�g��'� �>���q@f�irK96/a+EW���Sy�\(Q
����6HF������n��߿FɂчD'��s����F���U\ȷ��Q�}��-<]h�H���И��%h�Bs����5;ɒY����s�=C�'6��%�M��D���S)�g�o�:����u:���8�G�������Nqv1�v�AY|*��y>r2�W
����S�.Q8"�2U� f�ڕ���3Ur��0X���5*F]n �"��ԇ��r_���ma�d�7�!�z��Q����_(�%t��Ԃ�h<�K(�mgm�F�������� �����~k��=G�H�}K0�y��g���K�PP��֥�ī�1�>D2��mZQ]��$��_�x��@���+>?�Hl��H���~Y	�K��UkG/C��F �s*�d��W��=^�æ��e��N�
�,�
�q��p�@�ǚ4��8��^C̥��5���
��	S6�c7(k{q��|a>�G�by��4^�(;q}�ͻ)� �e~����H)ǯ��:"|�E�O��7b;)�s&xuS�wִ�5���!\�'dKپ�l|��!�̙٠+#5�ҝ�1j���񜗴)�*N�O���ZAm3���3��6�d���OĜO�V]8G���{i���p��/mŊ_�#���?-:�R�4�-p5D푳*�,˺)���;t�R��r���ߐR2A����~|>�F�m����<N���,�t?��#5G �l!A&>$�R<x^�㿜�L%x��u�@6I�/+���|�m��������wm��"*�<\�O�O�9X�D�wZ!h�������Fظo����,$�%��i�݁���A��X����0ֱZG���2����C�( �\��*B:A�$"��.G'�L-)�U���|��n�n����쀖z?#4_uI�֪6!���r�@V��;�W �X�ז�]�C?����ho���J��月q�Φ�O��P��WZ��EqkG���8��V�>!��mo��0�����[l��L�A5m3�W�
7�� ���,�Gkg4"2�״�O��K�Sܹr��9f�A�E�
3|
$�pDNlF�����?#���0L#�C��ȝed���p��ֻn���.o�LSi1n���������*)�P�)
3��b�p�k��W�R��|�d���<@�/�������K| ���<̐+���b�W���V�b��*tPN�>[���gyh�vd;6��+<(�3��rSX+t>�k��Ap`Ľ@ʞ_�ˀ��N+��I���ě!a#x!m��Sr�����=G��q�}Im�H����n������2p�f�{1~C�\ >��o�M�P�O���.Wp���#w�Q��x��{l�_�HPP��`�^LE�������u�<���a��J��c;ե:>t Fu=}�����^fX_��a�Yd��Ta)C� ����<aK��#n:�(�7 �U��U��8]�P���B�4'r;ح��� �ޭz�E�;�,���ɀR�M�$���;��Y�j�:�En˩ޔt]�od)u+}D��\+y�չt�@Ig����I�`��4���|
��=i��o�'��J_��i"���͡.a��Ӈ�$ܙGlI�H��mI!j��*��10	�f٥W�l6]���nb�,G���5��P�M��Gf���_2S����/ԥ�caÐ�_r���l 58n~A?k#�|_ ��rLm���u��d(M�P����	F��7P@�(w��3@6$9�5�E�H4����ָ)�-�S/
JA��r�s�~L�x`�������f�6B�ulВsv+g�0�� �8㼾�i��o��WdK^
D���y.tK	�TF`�`�a$I8wX+�Z��}�ԳZ���ʪ��<�m��'�n
*��l�'�P�$��%��E����Џ�٨�Ǧ�����$�(��GU9��)�����WS�P��*Jp~;�z9^iފjʫ��"Z��R� 7zT�Vl/��<�2�MI���� �OҜ���g�"�[ɑ�c�}��|����:e,M^�Z��F���W�3o��Ű	�C���璤�)�3���^`��i�O{׮�k�$��tF-ٖ�\3b���X�A�2����Vz�@��E1r�����N>����ii��?��u��8�;�CJyb{�h�BcnE/�Q�C����.�|Q���1����PGz�ܜy|��{ �v��ʷ-�zD�Q�����6DohΏkEb�&y%�03���V���a��|�i:�P0xGm�h)�>h�"�Nt\C�;�1����)�=҇s4���\�
*���ۻuʓ��(w�>|I�d%�Ǒ#'�o
M����uA�$ȰI|�5eP#�L\"E����x#%cC4�x�J�uc9X�����A�QK#�����^AyA�`L;H�D[���u��X eX5h�Dן�:c����M����r�!�婞��2���P��!��]��٪x̨���3��
�T��U���6X���JWg#��\��r	���vcP�e��\���v��G�C�,�ۛb���w
b�Z[�+W�0�̂�
���,��!=83��x	�p��{�K"Rb;�X����&�[m��Q:K_]t:Z�kV?ۉ���N���_ku�E�*/����9N�>N����8��a�g�s���2��ac#��G�V�|<]�st����gr�$��*�!�
 �W��o���p=���:���w�Ĩ-d0V�ez����l��:N�%��[}�(w,��5�?_t'��5?x��z�#n0i����Pkt09aJ{�>,����|]G�]KTr�s���wX�����{��׉�(\���Gk`�K�� ��
���m}�l9mL�>^�FDq��G%�S̔���R�[hO��7�j}$��be	s$�'�dNW%םw�M�~��u/0�����Tt��坍�
�F3k�!B�<߈S6�9UGU�/�r	���9pU�2Y�(ʯ���K�y���Q(���`�dr��u!��7nX����|�S3;-=�5r�%9ꚶ]��eM���]�
&�� �@$��q:@���{�h�Lf9Vl�+�CC^��kC��|���ݐq.���:��S���{�YVX��5"�����c�[cfʪ�7�;h���x��ir�#�,��9+$�%^�S�e��zY�H�s���0��
brJ6\�������"�R��`2�\(��t"��(jΟr���������ӱ��J����I�,����#��:��AW9�:&�%��?~7�?������R��R$�ZR�q?�F�x�Y׀��G�K?Q���:d�I�D9+�ƶgj&Ʌ�0xjU�E>������3з�yEV�X@'Uy+���9\��G>����?��@���;;,#L�u*p)��}��bH{�X$8�kKHq�a�����@K��2ʳ�F�M���t��G�>���-Wr�����[*֪3?h�r�uhL`�3�D��� �Lc��4<�S0���	a׷ �u�t��\.g��z�� 	�Zȧ�yL��W&�3��~�1�U�����nju�beXm�~�'p ��y�$��$��F{�Zŕ�SI�n���6�hTF5,9l=Xj����"	u7�2�n��������},ڄ��j��@��&]��f!}�옟��~|����39c����W�i�	�qM��w�à��uϝj�7λ�\��T&�ǖqh�y�.���)�{{�Ԑ��tnv'���9dO|�i~�:��},�i\!��.�N����;���j�о�H�w3�$�9�'h�ga�y�j3�ҥQ��
g� ��܋�<ͮl�)���iQ�	�u�:�$�����bi��:m�o�}]��Z<SC=�5� -4���EBK�Utں|� }W�7��'�\i��B��}�I?�_�ny��p�ݒ���4��4�S�����|\q���%�s{��o���V,>���s�S���m�(��O���5Bl��ۘ���q��%}�.8�n�r�D��J�YnV�r�=.z>ƕ
Mh���:�汳�=b��ʉB�c��d]���=��Lt篃���W/�A@�h�{�4w�:Y5���"#�d*JW6�en��q�2d���k�X6�e_U�W簗P��ϣ7�>��#��6��l_��yCm�Ki>\��2a���,�檻�A�|�����'�O���Y�h$���|���'�d �l+ـNb�!g_ּk���5n�'D��R����٩������_�4�X�4�?�o?�����\�� �-�W��@�5�T{�`:��Ŭ�|b��]x�c�k�I_����8*)F�t'����]�b2K�U9�?�*OTҎ,�-`0��m���y�)r�=եp�t�Ŀ>b`�2"��78����(�pR�oL_�@�Bg�	���tcF��I*X-�>��$�r�1"�_�����+c+L�8y�D��^�Pō�Au�'�w:�<l�tq�;b��mB�	
'����ko���Q�s]]�(����/(�!��i�,�8Ѝ�7?p3A �3��y��\L�EÖ�<"���&~���]?b����5~�0���(�(�Y��[����$î��wjx3�g����;EG���C�.c��o�֮Y2B�N�+�<f��MD�H�x��Aժ����yw©���±��ձ~�-�&D���8/=�SE���3&xt1���������}��i��8n.WǮO����2;;���j��B�3��O�nY�֏-�����5��a��k�As�c�u,}[SM�o��/�b�6��Y.�e�K����w�{؞�S�N;�fƝ���P�:���Y
�u꣼my3��#��t��-���xT^*%�e7m\�܌)���Φ)-�rBz���3�r��,+���4�l�d76�����.% ])a�E�C&��cg�!��Ͱq���o�ܠ{�q�U���x�f�ܨ2/k` �]�wal��5��y��.K��Qn�$�]���/�h>d���u���1�iH�J���T�8J��@�GK�
���HH;��ׅ|�G�m+5u�0UDeR*!��=�^EHf����=fO�V�Uf��C(`�SuF�۶Z��Г4��6�HS���f*ņ@�Lx�qT�k��� ~l�&���� A�=U�G���x-�FD����5lt�J׊�q�nڪlF$0^5�M��u#����Ė�t�є�r�-�;?����.~�"nN������L&�Qʥ��+����o�:?с��`�ƚՌ�;�cD�,��؅v-��{Z�9��%�<2�V�%:�qr;��!��K��ںz�e��N��"<��qx��b�Gaj.!u�HlxЉβ�k:� ��aX�v�qU�.V�D�,��%#t�)!u&�&j�6�j���K���h����	�F��0��T��=��6��顺Q�ϝ�sA�?O�:б���V�@�p��[�=��z�`E��ⴼa	�?:k0w��ˠm�s!��&H�k������� A�=8�&�>/�� �E�갶;f��U�����z3��X������k`+�����J��7<º��+�v�M,*��̝���f:`�7�����3��7��r]h�]K�$�ն@%+s"�[���2��'OuH����������a�n�gJv��ߞTiw~�Vid��F�N��xЈ:�1w^[穉���w��Q�Z?nﭓ�)��MAZ��j݋)���d���n� .��W�3e*|��"Z�6`􅔧`�WZ��d�|+�5Ђ�d�o^��7�s:Q;�سVW���qT�����	QHaed3�`�$�R�Y����ynO��֝?��/��f��f��%;��sVl���/Yj���Z�y_�|�lw}x8�0:����.�
���nD�V�O�-Gsǁ:X�Z��FR(��؞Zʘ����$+��b�Y� t	$�����(�P��g�B����xeg��{Ms�䳎2�./��۟O��Y燼꣇j�p��f��r�}�o�1���,ҏ<�N�2�1���W��Ð����g9L���A:O�c��Y��d��[����혎��d�f�n���iL&J8m��ޝ����id�fg�U�&��h7��Z��t�U��&���ҩ�%�JQN~�1V8�ߎ�xy�� {�+D���������O�
oY�A�0��̥�|=(j~���](�ꌕ��/?I�Qx�m8���[���Rϓ_�s�*&��=ǈ@��24D�fS�3qL,}7���jn��~?(G�g%A�U���|0�U�K;�?1�j�2+"��%���m ����H|��f�nUTv&�؞u7��M�?��J�r3d��Y�͏[x�%]���!�4u�x)��lM:E��T�rD`R��2�ߩ��#?��!E��Z�,���e�Q�zF͵�z�-�I�Zt-P�-���5�1�*O�2��^��o��cӖPD�(�ΥѳZ$5��J�Q�[DuV5��6�����@v>U"���.#
8��K{���ڳ]�\�O-Վ�n>e��T�zxb�����L$�~qa���j|hJ��ω��)�����#L�^�8�D�l�"sZ#��~*�K�O��r X��$B�V(�`���C��G͂���4��n��͸W�@�,�*}���9~x�ah�Ƹ��71+�b��U9��V�{44d(�ui��
9+ıx���^QE�_���M��o`D��6� �13�T)K��	�V�T�3�|���klqh^�z��`I�)�=f��xw
��c�	ss�Vr{�G���Z���6�yL����&f�[��B����\���e�vTP�v�_@�wLC���Mm�X)D�x^ź�|f��?��'N�'�ON)��SR�U����4z0ͪ��&�c�{� ��E�*�~I$ ����MW	���B�	�V�O!�ʌx���B�v��x�7kX��S�VA������ƕ�ҝ셐}�an�?X�e�[�y���]�/���H��s�u|H�9Q�����[Vx=���ʂS:9t�x.�mT��uOP3�˧�}S{V�&LvJ8��L��~�/u&��Z2�^7Hde?Vaǹ�0�b|J_c.b��f�ӻ��X}Pi-#�O�>��)�]D�@�
L����jjHzv��!��75<�L�s�}fq��hcN���>ِ���ҵS��xA���(J�AJ�1፭�%z��M/aWxE0������F�~�-M�5[��4T�1��[�#N�~�\)�&mw!.˺�%@�^lǫ���N)��x};���i0��"Q�s-rG�f9���M՟U+U�.���@�7-��K�S��c��#�+���]k��_|~F�ŘT�!��v߁2;7�k�,HH$��`<M�{���h�6��{�Ȕ��;�jie�PL�@���L%�2ϛw���Zd`���!_��5����Pu���<<��B{�WfФ���+�\��m
S�D#�˹��!�?�q2��إ��E8���=W��eb}�#۸naߑE�&R�]IC�9,9�'7��U����	!� ���Bږ&Pފ���%4p�H6�lG�@Qd�����7���P�Z|I�Y%������1gM���wo�����ǐT��l��p�7K ~��O]��q�&0�����Hk�MF�t��{Q�E��]�rair��E4�H���/'��C�
�j	<KKb����T�RP�|>W<2C0[�e�%*N�p<P��o�l�\s!��?�7@����������3˅��?��2`��{ҬlN�	b�D����a��Ud��xޔ ��#7��!m붩*�g��qm�Q���W�X����n��M� ����zէu�S����M߰�E��<�R?�ҥ�t֧^Y�j��N��>�X�j(���O,��y����
|G���	�VL���W(6lќ]�/�}ǒm��#�Q*���Ar�0@����!s4	`5�K�L���N9���Q�EH��� ��iy�Ф�gv��:�q(w^�]�%p�Ł�^���\���_"W���
�h�D��*|�e}��y�#x�T��O��q/�p�B�Y�cj�>�Fd�5q6��	�Τ����h缼5A�4t��
/�A$���5����#�������{��� y�HR�˛��Y�FN�1v`�5+�ѿ2,��+6�TՌMޔ�ˢu]���IĳCR;�[\
H�s��yE;��=C*
�r2t��J�-w�k��9���p�m�8]\�"�@gx����9���cK�.�~2c�Bf����wgM�T��z����;�3f ����s���#� /�#��˖�`/�a�m2�aBe6i���-�I�;g. ����t�ϑ�E��$ �խ!���9��U�MXM�9�q�Ϙn�cѨĘN��!�P�k�R#r���2Z�,E]��Q�}ܵ{=i�E�Uw�����p޶K0w_��z�F�.�M�9,{��׹U{�%ZH���pPu���K>�5� ��\1:
�k�Q
��X�1~�ʘ�۝�!*��&��,�%�����6�ݝ�Y��"�I2Aн�!ǻ7Cn�~B)��������o����(�-��f��LT�2�g^����I�6�m�c
��\:��
�.)�V�� tve��`Λ�6�NN�+a�B()�����of0E�,� ���[�FJ�)oĶ�|O�{��U|�������%{�X�:�4�Bg'u퉽C	�v�S��(
�.�fO}ۺ��Fi!A4�J�bI(��̢Mg�2'��9yB?����TKK���Cw�p\�xd|M����1�F�T� �^��KP�Ԫ�⥁Q�X��]�YlK���b���[���n��o��݌���ՀWShd�.�~S�&�tɦ{�`�f=�Nj�gTi��['tpk}���(�B���c%�~�!�VZf���˯��XP��T��"���J�ID�:��ak'�fɪ$Bؙ��X�TGh�D�r�y�e�*�����	�g���/��v�w�Iu�|)�z�&���KQ&A��}~�x�YC�����\'iƼ5<w8�Gx��@]y������1�W��ar� ��k)Ρ��ܭ���8��Po��Mυ�x��\�}}�~��@;g��j97�}�6Ou)��>g�����Qδ,8�q��?�Os]\q6i����\�d� *	 2��`��r�a<__Τ�5u���:d���Wa�;n��(�]#�?kIV�R����Au��� b�s a]ǫx������e�T:�l�K���u晃�4�l��<��?�Sۛ��/%�YR%�T��Xs}��ʝN8(���7�k���՜��f�$�#�
d��A/�C&0Z��Lw�Il@'E�e�NC �����"��f�H��+\�#[D���P�q\�*-�����x 2�Fgz�jt]�:��y�z�S��'�W��g���mj�I����Rͧ9�q>���Μu�j�K2�d=:(Rƞ��9���m21��>Z��Ão�a���U�x92�j�kνNPgd�jy�����>w�~��.�y��ʑ���C�_�FqP>�'�^��q�l�&�%3��,��;�T(6��yY�/V!��j�V�:�X�̥����	�3R��������U��j�Mߠ(���s�:6���-!B�+r�b��5w_Z��Ӯ���ͼ���*�9�´c��g��|\XW��Z�/6���}��hY`p�8�UUp���O��x��ߖ �����Ѽ=W�I�G7�@�XB��M�M��-�z�*p�x�L��T��'w��W�x?l%>4~�oB�ܥn��!v�(���W�t= d@N\c��r�[b->A���$��)��S/Y@����R�V(ӻb�A�8�~���[Q�1w��( ��HS�+U�x�E4�ܥ�����w�d�X�M?Һ��m�Ғo����Z���>,U~wE�ZZDR�Cu�E�0�&��"���I�h�d/s
o\ �t<(�u��z��.~��b�%k�|G��isn�Eq�1]��W��\.V'>�m�	wA�M\y��0�
���|��m�Sq�$����H�ݴ��oq �/�'���Q�v�|c����qo��e�v���W�g-���`lZn6i��8|t���fuI��������\/q��U8HD2�`)�����Zf񫕐r�t��PTХ�;U2�oh�e�O_1��J{$���5/y`�����F?RRX��z�r!���	���ڭ�Q�e�?8����sb�͋�<�޻\��.�2tB|�A��/��=%�)p!���:`o�6�����'��i3=����C�"I��!M�0$y؞Um���wY���1��iL�}i�W�r�H���%?g��S���T���	��
����?OS���m+�i��v�8P2��8�ch@��𽪸��mxY���L];"�"�0ɸ����侇J���Q0~��îI�y� ��_h��QO�ʂ�*����|����?����l1P_�Xd�jcԺ!=;��鈀Á;M���;��}:���u��먮<"K./�z�Y�O�ЪOdd�v �[����L������a�{����FkS�x]L"��ft£�؎�Ҥ�[E>fjvy���)���φ�<��������^t�q�v�O�D��ބ`g���'v�^y�V|ř8"�����3�d�����3C�S�5�q��8>����1$L�')�0tߣ�Ā� ���m�g`�K�O�=�Up�ʘ��S���Tg�i`¹�ઌ��c�H9L1ϕ�Xr����LB���Db�<��h-��;h4t�<0;�ه}���%\�Y�P>�T���S�D}K��'����1���y;H�}0�L}�3\H��9p��J��� N�k �N�q%�<�oތ+$�\�wo���,��5~`�|��j�!8h$iX��jʜ%zѯA������1��P؇�-N��I(I4�r�#�؂��+6F䦴[Vw(L��d�|�5�Nw��Lt��������I�����2}�\���xy<��w�Jo�s=aSf�!�s��jE�C2z��'W^R�^x۬����b�_v�O���<!`�ON���a���u��B�Q�)�������D՗������P1a���KN0�������	ntVj��D(����%Ive������%����f��U~cr:��<_��)ߦ*����p�c{���:w��U_s�]�_�_;�1����h��xj�`?w{�<�K�1!�CH݀����9��׈��lQ�@�O�oE���ק;P)^����L	\��2kmh~�Y���Ẕu �P �2���O�8�x)I��j�C��z�K2B5N������6+c�{j�����`b��,n��nb(������lcj�!�J.Qپ����zr�)U'S>d�8&(�Ze����؆��W �۵��~u5�Q�Ax�����|m��hGTj�E�>Ú���^��S�~o��5a�#��En.���^T��{�z���2��c�� %���:g���@��m���"��p3��j��9�Cϣ��������ʾٿ����P������7�٩Z|\�2`��fr��f�3��Z(��ض�σ�6����Y�QX��0/l���Yl5��#p:[�D\��b�x<��u�a�=��yQe��L�4~y��	����O�Ή��a�m��#4��BUC~��*(��q+��<��S�8�D�l6���n+�_%Ӯ�3ĳ��%u^K	0}<lƞ�0h���Stܖ.ӡ��R����W�$�$>9�~����l*N~TS����Y:3)#Օ���UN��>����}����~�������Wc��e�km�AX��ӻ���� ]����$�C���oL�0`BvXt�������͆���(c5?޼ړR�Θ��o��q�WG]xyH��-+�\���d�������[N��t�t�U
�bar�U��5P}f��}w����HR�ˢ6fB�g�ƾ�4uPn�qh�4��[��0o�����o��7\�a�3`�����~ex~D�$��,]¹�S���(��r��ٵ�b����������R�R��}�-��WTN���}A��m�g�ŞA����u�`c���U=\���%�o��u���)�*� �9#��?+H�*K4��������l��EKQ݇10����.Z���ֺkt&ro�LP5���ew���0��l�g�e�v�ȏ�q�>�<W`�*J��.S�rEL^���3�I���խ�xq=��P�\ �E]u��v+��|�x��O	���ݤ�d�y�{LF�5*1��ek2#��	��oƓ�)�a#0�G�}.�0�� �T���(+���V�>S!�rԳ��s�k7�hk�`8ϢD�3�?y�a��UJ�&7��
��5/�/'O�EJ�� �I�����'��[]�m�݊G��]�����#����U�1|����:`��ï�e]�*u�vZS�����/w��˓�e~TCP>��t�����_-�,g �-!�WM]#e�I����}����	'WDN��?Dn�:�wl�W���v��_+E�Bs�^����2'f�Sq�A��`�)�S�K���$�J�����ڊ.�A���+ANQ�ʬ^�|Z�O��z��-\�f� �j(�Y�
��ƣЁ ,�"U��B�S�xQ:,��?�>)���Y�_��^���=y?���ؤ���
��Z�_Ԏ�D$Z䘣�������߶Ɇz̪�觰��ܵ�;��qDei��J%�@Q�+~���i���& �j�u��%G�k�Q�����ᐞ#�ե���&)Y6N5!�F��� ��9�#�v$����ӄƊ㎆�El/����Z��uv�1����W�ȕ���qM�$fj"���t�S>�*�y���\�5R��m���J��>�X>	�o��3���ɬ+2_z��$�i5�
W��6Ng�M�������ڬP�d p'��'p��(^r)�(?<��y͂iz��_o�Llx$�]<U��I�]��'oJI}�i�.79F\�#�I�"�0}ul5O�l=�!ԉ���|���{���[x�ŏA���GwM�:��Uj�rQ �,��s�RI�T��]�f�}dQlމ�[Q���_<l��=��8���/*�ń),�,�=�$���B�|s{�/�Gw������:�Ʈ2v��k*!=iv��p��{8��T4�������$;�����l:lܳ����fsK䈼oS��ec�<2*�,÷�s3�I�BES���8b�ݰ9$�X��y���0kn�.c+2p�<¾�2�a�z���BF����c�"_=�h�ny]��K ��{]Č0I �-��ö�`Ν�C��º�1�!���8)����K(��S?��r@1�?r�i�i� $��<��3uP�6=���$�YJ>�ݕӣ@��
_�"n�$Wg%�,.�Ƌ�a8�k�aw+)����3�8��������_������t��^�{a�(�K"-e�X���c��e��&032�+7����F��mn�"�b�\�$s��2�j�N�)�8$U��|��iP�{t���{LQ�4�s�Q�G.�@b����9m)����l���{�a~����[�6ms� ����z���1R�0��7��W�^Wuy�+�g�1�f��:�q���陀e{�j����=7�`e��e{�É��MS��t�b�z7���ʨTG�%3�����	r�T�W�7����۶v�d�yd<p�j�f�����s0�zqޕ2��N7����$:h �lA���}��5Yg/�3q������"�#�U�?&?��A*O�	?�k!P��0B�L��$�Tf�V2�@��l�������1��5Y��y����!yL�ZEi$��I�&s��Tq���������:
h�����N���,��YT����ÿGW���o�]1�~K  ?��c��!�Q���%3�8��ϣ{1א�����.�_\����h��U��=����ʳ���r���Y��~K�;�G�Ev\⼩��M3gɠ]tN�`�⨜.���[o���� �<����<j k���αT�_�7��	љ�8�d�%r�-�G�V{����'@��L E�97Y�Y�LI��rxeU��G��%�{�#z۳�a�}�����+��>9<J����8���#�=H��;�A��vE�M|s��/�l���vE܆v�\k�<ɴJ[�t�Yn=F�������.�D�B�tʝ�Tk}������,MN���"�h�Wn8���ƃ��4����h'�'��h����S������\M�Q�D����~�RVq;�k�$������z��|��v˸xVY$���Kf���p�1b����*�'ح	�MFW۾�M��ӄx�8Gj'z��G��
�����o��E/�҇u��&���S���d��Q��o	0�iU�Բ(*!RC��F�����J�+�έ����%3���4�/��*Hn�^q9m�n\�N�p��b�[�"�A;���`#&>�C��-#<z�/c�	���p�U����v
$�a ��Y1��{}��b$����3�#A¢����t�)g@��0�T����E@����)%��:`�z�y�ϐ凨#��X~��ܰza�7"q��;��e�(&���:�fנ ����x���.��^M��=~���T���M�-2l>/RQ{��yG��V��Gy��S���3(X%�wpU�T�;VC�����=s���mآDy/z�(��<��Ͷ�|+����r�(:ܸ����C��7�#��_�$�/;h|���AxB/��}U!���h�ɍ�fO/��F۝�ow���.}Se�R��A�9�m�̺_ɶ@�@>[���2�#:�L<܌ſ(;&��#M�O=��C�I�2(�8��ي��>�{�'��0�ֿo\�=�˾HC�VZ�Bج)|�N��(DyF8}�"��7������I�Y���?��A�'r�"� �D�掷}�E��L�� .=A�iA!	���v�:a��gQs��wӜQ�Hk�<�x!�Ӿ�>�<k�Ve�k�*����ph�5t'޿�,`Y���A&�_�^⇨&�ڠo�mr/d���<��� ?�u��5��ؕJT��c�˓;��z���*��82�jޱ}�E!z��æ�u��|M��f�6N���>�?�l4�F��q�����|�q9�#�	����ҙJ�	��d͕�om�<A)�JI���b?�F�P�K;'CX�2����N�	�!��j"���z8��O���B�6]h�v��_O������'����ϟX$��Ʈ�%�� &�W	�'Q<b⪅�mʦw���^c�o ������O\�!`����O��c<K��!G��ҷ#���68R���V�c����`Ud�D_\?3)]�7�������n��ΦN ������0�`j'��oF���'�܍�)e!/�>*�.� ��*�v���4��ѕ����C4b���U#@������-!&����ƽ����Sn!����CD�Y�޻�mKw�J�Ufx�r+R��J��@����h4��uB��\�<ɯI͵O����a����������l������AqW�0oM �QPE�6�i���]���֌����v�����H"�yFi�C$��#���⠻���|���|,����4��zl�YϚ^�E5��9���y�/�iD܆�p���W�p�!��ՙ-���զ<U����g��|vV5��'^#m9��2.]I����a���V6�y��#ꢮƈ �"��m_�JG�UN2��I�:��K�,��{[�(%�S���N�40Bb��O�ڽ���q�¸����(S�����o��a�u?��/��N�i	��)B��}���˷�2�~�}���љpC���߯KW�=��0�b�I_6�4�����k=��޹/O�>� ��������t�cEi����^��KY	���3`5K�{d2�����(es�!���~e ����|+G؋'���>��8��&j ���tK�F!p�臬c��0�bh���¬���?�d_f	�z�kd7��QenT��\�`%{K����K�O�&�ZP�/�p�N��(B�g���=�����0b�O�mB�?�W�aJb�u�rek�1�ȉ�Z:�9�3I��	?�K	�Ǯ_�&�!����4� FJ��!��o�E��\�_Er/D+ӆ"/SY=�7TV{*��p*X���Ln0�c�$y�B�QQ�!�$�gѻ����m�<;��H$S��T�$= �~LWz,l6b`���<���OT��s˗��7�W��Z�ڜE)Lr�S	x�+\r�����E��������w I\���v�Ѩ�=!_�Q�;*�x���iM������ևX;��
�]��y�������&y*�g�%��J-�k�b������*t�J^��F��(t�@�V���l�\��I�]b�c�J`�އC�	��G�$DPYR�b�n�e���+���]���R�!i_��y�_�m��[p��z�@BzDěx�;�Ԥ�B��cc�%W5M�����D����^)���d&�����2�u� ��ФT�����ARk�fZ�AH�W�9��X��j�[J���B�oKt'NZ������}��_�*�Kz��r����� <��p�Qd;\���� q�T��{���E^Dґ�e$k�7��9U-�V��C9������2=����ƑB�Fe�>iMw�\��B��9�!OF��mD�ʟjk�	�� 7%vVPDG�8X���Exۃh}�����Xl��P
_���\%�C��9�\#x��L������΋kH�J(���x�k��o="$�E��A&Jl�:�t������
�Db����#��ث�9��D�L�ښ�j@�%�l�J�mfM�Y�xd�@`K�M��wI����N1�L�h�o�P#ެ?���d�L��eh�Zzt}(Q�J�{��K�����7��L7Ӆ�	dA�%=��cz����$��P`?rb����FN�%�Z��>���&���2Q��H���&��v���|�y�/���\UC�{�O��|	H��]��T��@ m4�k�á�:��Uf ��K��~�6��o�f�-�]��}"cx����ɢfRU�o� ����K�'�t��Lӌ.J��7Cj#����{���w>,���i�D���G
�JI�7�`���ĝ#e;m�3j׫�p��h,��EH�~LI�Gm�t�EUSC��4�9�tpXm-�h��g�����O�|CV�#y9����쑌h@��Ӆ��?��>_F�b��gm�X!^V�'���q��!k��!8>����IߔKR�z��#W4�B�J�hƁ��2��q|�"��"AƑ�QR�:�ιq��� %�<�1��YO�����8-�	�CM+��
����txv��;vbM&��=���Ķ��p��l��Iao��S�� :���<i@]A!)=�y ��,.� �x,�,�+���9�nKfq��ٴQ�q��c��G��z���)-$�6����<���:KY���{F$�!�$�vb%�7Az�l����8�����n&����hy�E��j�	%cÈ�R��l��k���-� h�~Lo��3`j��$���P�v^M_�x����@���(��.-����3{��a�/E2��=;�[\��Z��?�VD��+��T r�1P�����k)�z8q\���r� نq;J>��)��)F����Zr/=��>�lt&�����pC&��H��XL$��S \�k��!W��J�R�Kx�81�l�UGV�	bI��l��g2u��jԹ��=�=��@l%��(���NP��_�,٧\m+%��H|���4˜�?{�C��j�^����7��?���~��90Y�~U��UXeI��lr4�T� �����V�l��v��X�M<jx*" GP]�0o��J�8�肘�Ce�_�ϨyPL�M���I�2;zuy�j�z4�j��� d�Z�W�Ϩ6�����J��{��T@����F#b\�)b�7�q����'����P/������ұ������ţ+�5��(� l8���ؘ��0��EP�ߜ��u�?6 �#��IAvlm�>����>E����%�m� �d����zL�Z�H�T�*�u�M�X��lw�@�Q��y^R?��{x�$9y��yᶄ�ڃʹ=������L�yz? �]h<���&�i!���P�`��I����-&;�[��O#�(���ۺ�Q��Y�Tf�AO��o[Z`p)	l��>oUalԁa��*���+��9n��Y"�#q{���"�wV�w����l�C�T;��t�oB����]dn���'��=�����A��}A��;���֨!���3�9P=亁Hwb�Q�k��1R�/���a�9v�$�Q���K*��O�ͭ�	��s��E�[)w�$���|=���!��enU�A{��Fl� Qg���#�^r�\���C�{^���A��~���[��gu�*���QM+v/�:p��;�!?�wJ������h7*��l��'#�n\E@���j���MS<�cU���?���3矍�Y�-$D��#mls>�x�"߫�d�>��y��%X�S�>��� �E���T���[���s��ï�F�_
B���S�%�ľv�p�}���dO*^V:xY��%�pc��e�q������@�<�@/��p|��M7��o�ӝX�s1%�ز|��aA�7�g&����O�Q1Xt6��;~>Y)d��ƞ�eqd&���#�@yy�8�\{"X�1��I�8�R?d���r�{�y#��G�{�G| ��:�V�K��ȟEܖ`V}	��Z�&��� ���I�:��սܝ�4� j��Y?�\�����l��ZWa1
���Y\�&�%�-Iӂ��V�>P� ��t�DL�o	��	���P���A��$mm(�C*�I�9�z�z�=�����_�� ĝbI�83zZ�v�EM7]=�%6������x��T\�A�1p�3L�@�Hz~K� ߺ:U���3ti�����:��Ho�[9q�&��~��,:���/Hg)�fq���fE�W��������?b��s~ze~#��)>��,��^+�!n���v��$��$����~��x���� O&SF10�d+{j���<�]�:�zܞ�]'�J�4wx��wI�R���
��U!^n���?v{���5�(��,��� _9@�CC,�u����Ғ�]�@�w�~%7]�iu�!�)�=a℺�{L wYN(R$�0�u�w�~���?��⨸L.��,	v0`C|��5U..Q���u9H�Q�⩢�a� ������;������NZ�L���-��<��o�̝�s��hy0=�h�a��b}c���5*_2p���tG��{O���]~CF�^=�Kx��2 ����	l�R��r9��ˢ��%�ƎP&��_T{$(Y2���i�s_bŃ/l���D��S`�ͻ��&�j��܊f?f��pR>3))�?��~�r���(uC�!m�D�%����U9�T�]�Ȍ��j%�m�a���s�9��f�>�E�7�+Vw�O�߾�#j�h�c�W�b>�����A��YWG�V_T+p����j�u:b�Ҁ��?u4B{z�')`}Kva�PƿU�N�vnʏ:%4�B���r����w�XV�ѭ������3�Y����?e:_�2�s�oςn�:���s|��*z��ZO�����:X�����D���X��5�+�[�BP2�m2�� ����?�D��" ����;�J̡JS=�5�2D�z�>�e�t!H������9>�0�q���c�6@8_���c��z�88ї��ː]_E��f��iJaw(+�u^C�i�}��a���0�y��M���?=��-���ߢ%�bY_�Z� �R� �p5�w5�����kO-:,�^�����vk{�oq�T�2N�ઈ�k��G$9|U��/�T��3T�̠8F)`#в�#�s�4�Q*#gf�]͔q�2�m�C�H���W�3����VCbEk��l	$A���̔wȈ
kӾr��)�'sL,��!��8̈Vl�{��}������V���:Cb�������?��k�S)��!&/�>'dF��%.$_a�3<x�y�(��)���t�|��ؕ�"É-Ggi;�~
w�i㏸QG}��>=,;m�)	VY�?,�k��ڞ��)k��U�^�NpZu���5���$$���KY}A\E��G��v�6�������4넉�=yE���ҥ�L)A�'	�R#�	�p�)&7,׵���Y~5��|di�B��<��J��X�.�ϧb^7l��J��wV�U���k�6f��eF�"�M ���K�?%o��`�>`�B1�:{�j�[̘E$ⲽ���'��q82����y��T��0)C�/�,����n�/�ek�,��x�;6���^s3�!�W��h�J�=Fx�8\/�^Q�X_G�~�m�Ru[�2�ɖ�EsX5��г��������U+��o#B+�v��ㄶ`p�М?��hT'���D���]f�!t�<|Ml�/M�Y:_l�C����1"��T�
&�:����{��ڠ�Ƃ���I6~-��sC���>+����ex��R��L;'*��~�����F�&}�Xz=��j?��W^)�~�ǄS_X� a��h�B�A�1t�^����:���Mĳ7m��r�;gUDLX9�o��{N�r!�Ҿ�w�:��ss�XPA��_�1h�e)"hҶ���U���E�dYȗ�I*s=��_�K����hC�D���|�M��{����D�&�w��1Ξ�R�"��ˬ��|�a���B=7O\�[���`��ku���т�笫�����C��C��' Mz�x��H��T��^��<�r�|p�C��	�*�'p�(�/����jg�o�o��a��W����f���y�e�)̚��8+�����J@��컢_L>���1�Lw�?y��H��̣]6 ���٢��'΋�G�4�R��>�����S.Ӭq�����l{�K�&k���IӮ�Hmup�;�<���37�5���(�C���9n�1����}DN��2 �jk�J��}��Y$fo���E�U���C��D{�ǟ��/��;��=��&��K�_��6"���$���|�rB��y�U.�͝!׭���B��
��ُ����it�_�k�d�֭	-�l���h�!KSҒ�;r��̬��g67.l�'���Յ���b���@S�+͡t�ͦ�o���k�VgP{L�C	��	W�c�9M��/5 ~��J�� 6ZF:"����e>L���{�m�D�?̲W�����>�]�	JZN0=�S��oi�r#��vJWW��~af1[Iig࣪M3`���
�u�����E^[T�{T%$��Ѹ��l�ZƳ9au_E��z�Nqq��h��%�*-�F�?��e>�JDF��te��5	|�-�U�h�I=LH1(ek����9� _��Y���R��b,��($-�ݖ��{>PH���;�Э٭�]�]t�sh��y�N�M��U��s��b�E��/+M�6Ya|���/>l[�>�d��'iZ�GnU�c���1wO]`�=���Pמ���s5/�a
������_<n���@���\ε���l
�.�Ph����$ۼ˽�=§��{��e�Ğ�p�!�\�F-f9`��$��'�)<�n6| ���[�4�.*��-�"�-l��"x�uD0� �j��d�<m�5R�St�K�b_m�R�M�q\!�\�� ��^�����Ͽ��.$�����r�阉G�]�h~��M�㿦U�Q𑉆�vW��R��r����|e��.����;LrS���qm{3��Noų���M�������A�U�v��޷IR4�?'����ы��s�~,��|�8��Mz
�9�Gd�<��LhnE�	T?Uwb���1�"3�0��`.���;���̢��
��9���Wv���L��g���IybW�l9W���J���RL2�ُ�?�g�9ǎfE�������x����{Z�cE@�oY��{�$����+��^V�5��0������I,bf���"X����+Mˮ��L��x�cID	VYN_ؘ����-G'���6���*�a��O"J�@{�x)Y���;}�$��k.�$����i��*��y�,���aB���]=?K��P���}�%�23gz����
)��s�|{(��!!�K@�����'Gv��`+����]vD��{��s�L��̋���8ѨX1�JA'��� ��o�$	Uf�؅��:~�9����d���j�%���o@��{)K��d̩�e�IO�;54�ků�����~�yL�[������"���6�V.�4� " s���\Hy̩��":��ώ�_�l�9T"R�[4�Q�����q�B���$�$]h��}�����O�&�,UF~vZ�[ύϻF�p�>��'W��/�8raY}�7�gc���Gt�8Mc���ϒ�oe<U�3�����i:Z�ʨ�~"�e#��%�Kiһ�+�����J��l��z�幼	����}3�OHA�6	�ٹ� �Z�̅gM�C\բi�)� �$�`f].t����������|q�ߴ0-�N^!�%ĴnD��9*�A��I1qmG!b�;����Vk,�Ҍ)w2��UsX���M58��+Vt'c��I��Ƈ^��O tf�Yp��^�E_b0����P3kͱ&�rP��P]�I����Z'-�t��pu�164VE|PH�w���7�o��{Dc�� ��Q��͋3F������p�f:O-?;��tc�\�2�ř�W������܁3`�ٵ�?�D���z�UT��m����"�Q�r��:���A�r Z�7_�ÜC>G!	u���}H�D���t���|x�:�|FJ]5��A���[��q{s0O��_;W"y�ca��r#��<�2i(���AsKf����r�I�zQ�Jȝ	+0����~�hG_��ܧ��tB�k<*���)�`ͮm�-�
��t�����u��n|�\/6�6��{r��*���׬�?���d���2�/��x�#W��w
�"�K�� �td��%�� ���]k^�5�O�9+-�6�=��kH�LZ��`��4����Mx-���i����SsO<=K�O�����n��ƓC��G���=@�b�����ן-����P1�ܽA��>z�-��U���d����g�W?;F�oEt5�~x�	�	�G�� v/��nm2��>�葮�baJ!~./�t��a���>K1�Ʈ���{��P%2��R�
�ޭU�J�\��{��3�'��WͶ�	���#��{@�����X��)����k���u�E�@$�"��j��ARƧ��tbȡ�����z��\4���U�����5]u�ux�ӵ��A�Z�&�Ύ�4C"H ��I��E��%X�(���	�_>̓q�5Q8q�g�n��0���	@�Gٗa��2�AP|���V�2x�]�L��lǔ͸��k��'	��0'��W5�U,*O�*��z��7�<��h���(C-�2í-E�Ѕ��ר�y/~���v�T�HdM���^Y#�D�х�(�F����
KA��qX�=��1K_:�a����|(���ŋڦA���6%�RDY�8����8{�s�҆N�(��	������}�Gvj^v�]5Vx�ah������ߩ��D��A��6cʉവ�}͚���ǧ�C�)��BII�R\&��ԛ�X��o�s�\B�r��Vru�0��.����Wh� IT'M=(�V�����HkL��<�<�\kW��E5ƅbLcVfv�4[��L�բ�8���]'���	q�����g���B�o��~<�5DF%DQ�D�ˡwƥ9���#z�gsp����ډ/��+�Ў�'h����ָm�|�uE�p��FGlE�<H��t���NuΣ��U�%V�	X��n�s�9V+�(f��E����0�晜x7O� �f
���*��e�.9���Zs�����7Ǉ��V��7�͑�b`ȓoN4I��A�\�L���(�3���~�(��>���^��3��ARo��qq��r��odg�ŵ�\�"�L�3�r��[iK�QԐak儝�~�v�Ln����T�����[�p�6"�%?��
u��V�z��W��h���]�b' I&���j���$�>�1��wH&	��S���`9{~V�5i�'C3PH�����L|�μD��z�A5[X�(�
я�J�dzƞm�~$�c���sz:1��G�:���K��Jt���h)$�a=�5�)J�ta�8u����!������3�����5��D\�l��"���~2)��N�?/��`��z�M �p,��Rc��z��4�+���G[`*/v>&\3�.iH�� �G����-M�bt@|���N�Q���}��.V��󭹮Żbue+3�����M	p����$z�q4j�0��L�?�u���7*Fjr˕d�Dǂ)�������r-��+򦽘�ԜUqȔ�VIN�����g`C�=��9TH�09`Pڢ`�C!�/�5蹒P�g��aSLV[+o����ư����:��]���L��E�C!Y���6;���&=�@k�S���$ˬ��NM1%PH�����"ȹ��"j��q,}ĉ��� �C�����\�?��Z �0q��z����NJ�%�,##� �����vIel7�!����'� �c0f�k@򲰍���|I���q�(4��"Kh�<3͹;�@��+Ia)�h�|���E��-�69���P��>gNjR�t~J�k��P��� <��z�V�;�=��NZN�`���<��5%ɨE��:_��T�+�w�#��D9D�4��bΖ���e�9|Fr嵂�$�-u�r3QJM��*�Hq�z�	GO+��Q��/����88Yҿ����4LI+D�Y���v(�n��96�}�����1�bܼ
���7��0�5�5(�t�M`n�(-[($����zX�J}ܱ�B��lB�]/���W9��!G6pZTSo�yB��͙�W.�9?&=�����J���n��a,�6Rq�T�y�8smx�##@�/���aJ��EA��~q�C!�%{خ��O��=/o��mw��Dغ6�v�Gߓ��.iܣ�A=������K}CB���;v�ۤ�;F�1���n�L|ɒq�n�]�P>�d���E���������0m/ ^j�e#�x`�K�mb�5L.�L��_��퇺�4���b.���V��a���U��&y�E)��L��;�)�m�fN������
oE�P:��B�	AN��F��uth�
����}8�.��J�p-�T��3����W�T�J�2�P���)W��%/�)�z�l�N���9���h�'Όծ7V����U�B�|��bխ�g��yH���1\���+�Of���m h- �b��;�e �n�*8e�~�¡-�y=4'�f�i�#��ನ9��Wg����%��>��XWS��i��9�UL������q5Y˞������٤}�(��b�� y�7�s�+�R@-��/@��������*X,+��ci:�~BL��'����T9����jݩ�"���=p�Y8ʁ-�Dc�k�5#bj)l-Vs���������Dn�Jp��#�y;�nA;�m2�~�����8`H��Dh��gTJٹ-�2��G�\��)��ܟ�y�;Ix��(.@!3�D��i�EQ����K��VK�����g"��>^A���|F��Y�i�)B�����}��y�鍡J�m\���0ylWNCT��ṗ~�ߋ�ߋ��$Wu0�����ƧJ����1 H�<i��I$�4*n����|��B,C4-�s��k�S�����t��aF��5�ҝ�]�-���szD��zF'``�G8U)򸐚���L�V0N�'�f�م7�?�-/�rEX����c�[G���CPnyRڊ{eT��ұ�@��*_�!��
�·q)�� ���(&��c�����4I#V6K��i�"L߰l�OH�5����/�K��� A9�Ǟ��յ����b�)S���Ib�w�\��|����0��,��s~ת�(nq�4U�fl�$�������.ZV����rt�&��.Q/o��x�r��i��.�<Id�@]`L1�m�"��ˋ͐Cj��O~=켈&�u�g�Q�����3�ɯ͜���rL8I��1.l���������� ��5�� ����zw�b��s�L����y�X���+�׻a��<�aEIB��<dN؂��J���$�ʎ�D��t��Y�Y�� ��{�"M�.���L�-�{�
�yZ����m�����4xO�;nYo��4̩0rO��pi�nY����)�I��%���L�L��skԛ��)�a��)�.N�*�!M��1��)d4c�Y�aÎ�I�'}���u�����y��6��* �j7��{��mi�aCIvhF尃���q�J/�c�o��f��E �	u���^�<*�HtESwn����۞d�#nd�����㹭Z�y|92a�Ý���O'~0�8oj�2�W��s⃤��@�D�.uuh��i�]�|�|QH�ZŸ�j�% �?N(�͙;�]��5L�����3����@ˈd�ܻy����o��N��p��K`^�����������瞡��#1L��y�� �n�b�ϑ��K���*�5��Ӽ,A#W�ǯ��Z��ו}��C��]olp�2N�����"�̻f{�t)n-$�^�.m�>��nѝv���b��>U�p��������.Ȉ�Z�fZ�f����8��֍t��OD8gk+79����D>�}�:��#;���z�~꓇<��`U�G��8�o߀����V�l��Ct���6��`��ӚM{�*e�l섫$�"��-��c���S��9g�G�.jb4�e���⦖!#8U��1(�����h�� `j��Y�����I�kE��y:eth�KX�� dg�q�����z��t+��G�	 �oY��|�x�{��C�*5A�6Ȕo�]x�����8>��:���!$9����L;e%�v�ѐ_�#������4��X}�Y���%�)��!��8!�}�Og����c�+�|��R������j�'\��j�!�Ͱ����Fe�t�K`�G_0T��<�	cPMJA���HS3"�0*�tp5�9�Y|F��S8p�{5�WI⪝�ڹ�M7�S3�������:/ܷ���Me���QB+f�|GƲ�4ʕ�������)ʧC��41�I���w��=~�l�w,D���gp�H׫'3�[kB�⪜��,դI�ѻ�,QZ���߳Я���1��@U\el��Jϴ���P��C&��-{�����|Kc십����#��k3j�Dذ���k=L*Q�rJ��)y����h�����Ie�MB�3Q��j49���Z�J�椖��7�������@i�M#�)�ڏ�!D�XAi*��r��4��4���<��T�Z<O�be2�N�M�Z��m%z�z��< ȣ�#�E�I���|��c�Ba[�����i��dY Di��}�*l7Q^0s�q|q�q���� �+�g`j�o��ü_-ބ6��[w��)�ǆ��Z#��RN��T�ֽ�H����9��7�$��	[�k���pIg<���wt��0~^GW{����9? �3Q��\ʹ
,��I��J->�-͖���6�	��ٖ�9㘁�dU�.������Q��0��}Φ��A������5��x��1j� ��;/\���Y��=����Er����K���@������1���(�I�8�a�"?�죄��2��)ĕD�l���Vz+���5P�|��v�)7����m�R(!n�k�10����(г̞�ü���:�˥�$����@0���\yB ���-�H����z�� * i�u���U�)�ȏ:�.�L���M��m�!L�"����]�A�֑L��c���P�=�ػ�ǥ*!�?1��h ��	^-�����g�����1l���߃׏�j�6�;���uSoA^�%8�5 HT�aB�Q�@�v��c��u6P:9���t��l,W^A���}�X���O]�$	�©��<�r���F�B-J���r���,��qk�X��¯��ɖ�.C���|�����"���	?��7�η@D�����%�2��/�v������b!�<vq�Rk\ 9z��q*%;I}��b�m���X�%9	դ��l�(�׏��rY�0�BO�|����X�������>b�ӒcvBC�]��)u��� ^�\��'������7��1C��z�{��Z���e��)��m��T1k>
UY�/��IU<�e�aN�bE�ę�f���EBcc��}h�v�Tk�¶	b��*\ �E<W�1Ԩu�T��2�:�]�8�µ@Z�&G[����/l���7���:Ǘ_�>�_���E���}�#�HlM�E6ެF��E����3���
������Ì�[�6
����UGJ�`*)AX��jV6jh:�1?�Ӳb9١WPf>��*bӉ��ރ���;���$�� )�s����
������]$:�fƔ��
��6�5���.�G^��V5��O������a0�	�{�O��N���ހ��U��Y���,1�,�%�l���S�$@R{Y� Hݍݨ��ͯr/�'�H�~����P�f�	ЧQ�����q����ϐGB��z�����@"�	���m90�փe
���Y��XS�w���g��0v�\����<��d���q;�9]#�-��*�7�bЍ*���o.z�U�����;����O� ���
Br�6k��l(��F�$|��5��)���!�y_��3b��]��_���}�ZG
	{�~"�Vkt�i�5�l[J�m�	��DF�{a���H��|~�{��'�$�L��G.l��y5�r_I�S;?x�̺6�S1w�7��ٿV��7/�.����#7�~�a����q'��!Z�(�2��_��3��đ?]TR���n�&
R�`�Z��x'�SM�-��{�i,NG�h��H>��NMZ�:*���� }Y��7�.?��P�ߵ��/}��e����ib���^6�4vY_0�ϩ���]�%����;�F�n�8K�pv� �J�Z��WsW���M��ʼ)@y<�D�[Y�:dt��|^^^G4V����Tc����q�t�L�YP�m��2���e\3�Z���}��5k"fTl�����Kj�����c�3yK+{+���N�fbd���5@[�i��(�����-l����zQ%O�Y�7�F΍���O��LKqE ��K��,�-��;/cIe:%zw�j�1��2f�8���x�w8��I�z��#��?�r{0�FE�D�X�I�
5qy�(^y%'yRsJw���KO�A'� rđg��&�)SX����O�;#i9?6R�,��ni}.�XR҅�M&���|i�;A�d/�#�k�N����uD�F�G��j8�Y�qPˌ���d���)ٯ���U� B:�*�J�6cfR*�⭘,��}�a��ã��+^���v8[�ð�^_-�7S���g}b��D�R���L%_��?��xCvD�3��%�l|Z����j�h2�{w�W�����W��q�L�N������¤����Hb)B!j[�exKh�D5��(�d��Dh�ʤX�3�	�1�c�����AT�O��~��n�I�f��L�h�u�|n�<�Y(d΍�u��@}���gW�)�+<���)\���`��"w�p�����+��+���R���Hd^>�Q���!J ��y��.���J���7�YpQ����M&�p��1b�{~J��K�W�ԱQ���	ZGVmi������?��R4�O�=�44~CN`�ac��gC3��%����Xt��}�Ɨ�p=�����>�@+�&�k�D-B��p7�\�_�WT��;�$.�fc���kp��pYE3�~���oF��$s+��-���?�^Â����k3��N�H|����ƙ��:��Я�}�,�,GR9V��zU�����+n�����zl%� �^v����wԚ���0y�t���
�4�.ʟ���K�o��%>�I:]��@��EfQַ�כ!�Yw����v��0���n5LL7�m@� �|�}��I��X�s
�΂���tH��H��I�j����6��C��N*�p���J��fG$Y)�_�ݲ�!�*�s:3�j0[��3�<�k�d��u$2���DQ�[��Xr^�j�X?s"�.J�֩� �񂏰�J��{�N��	�ib.~ӵ���Ⱦ���J���Bs�)Ӕop5ؿ�_���J<�J-�~֘��Q'���S<��-؈z��x|�#Iř�{�,�ͮ��*��8T|�4�):`ӏ9�lI	��D�.�M��I�ۓ����q���}�K�ↅ-)���\�b�4���R�Z�w}`tz�-5+�R��H�p������<즰�d�J���葕�b��Eb���4�Z�r�w哏�v�S�᭻��s�/�C�H�V��Cy	�~��qs�[pk�ǌ�)�a�X�{C���Իo}�2�uΊ.ܑA 	���g���N�����R�)�s���y��uپ߲{�n��u$-)��M<A�,�!1e���:fF���O9�Rx��H��)��-�N*<�``4���Q^j�
�s�,��-"cn��1q5��ڈܝ��
Cy��8��Б5���D��e
`�U�f�"�Xm����+M����/��.�羛�}�D[����mښ��z�3�Kb���I�(8Df����R�wϠ�8�ϝP��S�ߵF�x�pyp<�rGg���&@�+4I��=S�$˚��P�@8������l��H�`ʣ��@%�4PD��C̜@��r���QM���x�7|��n�q�"b?$�nw�e������>|�}�?M���Ka�<��m}��k�р�K�����e�=�mR⨱�ch&Q��б�������6��?(sxť%`�CR���E�j֫�R]�x& +'���w����5fx�-i��ӃM���ݳ�����^5�uT'���M)�d'2�,�uE	�X��"|��$�䭟�
�}F�	&i⨡��'�<J���!P�q����E]��&�ZF�Dg��[S����Q�&IC�ҹ�4���<B��yR4e'��Zm8#��P4v}�#��_�$�gT�|e�P�8�fhQH�bf��^�|&:S������K�B#�lTW�$�u�B�x��h����s��J�~RJ�mJ���!?3p|�LhP�'�\�dq�=�/G��* `]���ާ@��2� C�K��Ǩk��{ i�>��%���N@@��g��/}`Oj����7��J�nI��M�Ԉ�S-`��T���k������%C[,�h
�@�!�!��� ��V�C6a���	 F���)��{�Z!����ƴU�e��kxx�弾�͌�C�˶�st��v�nE�XZ��:�\Q1��&��o�j�ԏ��\��)j�j��PD;����0�\:�L��'[��%��\�=�c�r����-��E�_v�1vn��a��A�aT���a$Q������ )C�[��d���m�<j]<=���cϰ ���K(�[��`�N�8(�	c�������K�6����!�; �3��{�g��y�����,��"4R�8���g�Vǳ�����O����Q]��z�N����<��N��E[0���X�f�^� �(���w�:;9��F�W�/����wj�yt������y<��+qPԄ���G浴N���l��0������]��GMV�y��>����K��2��ӌ.LCe��k.�2q�V��Q*	���Hv�W0XB=yC�(���4�|X�}i��ǐb��@Ӊ`�34U��{g���B�%�'ƕ����ipC*��:�f������Uĩ�B�]�_lg�u�6��	�D*��e$�������K�|ۀ���o�ڊ?r�O<�do�F�s:������.�#��`m�И`mE�!Xs��#�:�$+)�#��?8& J�Y�찆Q������s���q|u:�D'7��� ��^Y��&�.�v��q����c^�9��F�R�g���@���d3'
la���@�u��骵&���Y����'[���Hd�˞���{�N��!����0����H�I3G��/���Z�w~� 'F�s%��^]d���� ?�®�U�꒾{�ČF��CFɬ�� �t��V�B�/ S7�܁\νRi�w��g�~��1����b����W�R�4�x�2�7Bti1έ}d�?)���5U�#�8���al՚�&�ê^�� ��/�ڱka�2��%y�<ݞޞ�XKe/�L�U%~��Rs��ד���*iDnx*��?����M����A�����]�Z�6?m���qZ')�Mͩq���Qa�Կ�"�zA�]�SQ���1��9�|��ٗ��hxu�R��f��C���B7���nw�(��*߂�p���ħ��2Fx��U�{E2�3����m��yd�2S��,,=լ�W�P�S����+����R<�y�f�w)�Zw�l�ko*D*O-?9�bO�	��}���X���G�J60���bh��\�]0�vTL~���;̄h�7��T�L7�9��_��q(�r[���ڒ�A =M�1,D��FmZ"�P��(%ݼ*�\��n���L�=���q`G�/f!�����K��s�|��&�e�[����μ���d�KH����f
�"5�͌�c���w���]%�&��H�A.l(#%�wn�b �bs��.���+�ǻA6�A�����&"P�o��\P/@+�%����)����G�s�A��h�!LΦ���J1ޣf�U��["" ��q�U�.?@�-�ɋ�9�:�I[�:�1/~�S���:�kY�=Ձrۦڒ��F�*g,�N�=Z(GӞ+FWR#"���]Qj^�(��ge���K�-�f�(����9�<��V�Z�4 ��\�B�B����B�ɛ�ۛ;��k��Y-�U)�E�d���[��ˍv�D�m0��aT1F�h�pSzt���aARp�Qo��ޭ��d�.�3��,��!�`�g)Ge�V��W?�2%,�z�b��~��A9?�Ĳ�j��D�gj�hAj���_H3/�v�}z�W���G�Y�t����}�?L8!Z�p��T����8�Ʒ�ky�V��K7xc�
i��2���҄`3��������� �	�r*
\�댄�fX[����|��w�������,����l�߲�}��ɃPDl��e�	�E1!>�*|�pZ�
�����*`�
cB>�G�9��GU�b��S@������_5Dвj�0�s��ڳ�F$���(�g��u��ɜ��M����D�O�A�.I:kQ7�Do��9Q�-��=�@X�!|V�NO|l?�L�c�=��g~KH��Q�^�3��>�1�%�DW����r�U#�V�:l���V��| ����o70�A%]�u�
xfR�<�`�4B\��4L{����G`%���z�=��r*��bQ�= �9	`�P���?�@���@�E����.�JW$�OP{�Zꂬp`=(���4K�u������K�!%�a�N�lN�]
����=d��9��/��2F38|�qNS-A����:Vo2��B++�5�ɱ;t#<��%t��d�[5��:�皘�Zw�X6��9x@��k����`������ҎH�'������+�b]���ُcP�M�u$�i����b�p��ȸq�>��c��mm���O�&�]@�蔹�~p��Y{��.T��Ӈ,����m?��(N������GnOy
V%N�v�\5�W��~�����Հ���큗R�WU�T�2����@Aq�gf3�hJՋ-Qw:U�"!NOo;(�BW���9��gV�vWr͝S�s)�z�ɾ߬`}�����"����-�r����g�1��"�����ow����鉶�J�b�8�/w�bu7�����3�lx�XRȖ!��`�[<��Z�f�(��a%.�N���b�U�2]�l��MF���:�����ԇ�5�S�PB:�B���%��H�ϓ�� -��ӌB����-z�s�F��f�J�3-�4���\�u���l�-�͙i�|�D�Z�I]%P��[�ؠd�!���Ho�RMT�4.������Yv�q��������r�X��=z��Г|A��}�
�	������>��s����fiyO?:���ݐO6P��Uد��q�J�.��P0�/7�-�C4S!�Т#�'w��PV��w��~0d�Xť�	ExqWR�Cg��:2����6�	�p�r']s���.����Ӻ�D��7�{)�5CZG�,-����V��<+%�?��[�\|D���[���O� !�o��6"��ةu9�ϻiR ��aĪd�P�-�����������R�m�V�ќ����3Z��&��y�S�q��p<K��~Q����g]V��,sW��˓jgh��/�?4�ONUew����x�)��U1�u�>{vf�p�dPJ�ﶸ��!�
��=�sn+�RA�����3��+�>�� ��b<K)��d[��O�~�PN����`8n-���ʏLB(D/*�)o�Z#�+�2�i)�;Q��\�����Ee�-���Wp��ЌTUi�RC�B�l��Tw�<<CXmNk1m��
�/�;%�Ι����c_��,n&�2�O��m�3�"=��u��CB�+�o>�[|�c ��H N���^�)  �y|�N����TS3�C�i�/Q���<[�ab|H���\M�!�|e
զb؈��J��[t�X��1��{�L��t���#�쐊�4a#��+{^���Y�GX �?���q����e�����_q0M�@�eag��F	a�i����Ϻɚ3���n�,ӱ41pE���<b�=bjF�#�Mx���b����
�	.�7]��b�Y���!�<h�_��PE�n��^��*�x��-�Օ!�#/g�lTD�d۶1T�.�Z�
X�m�@�q���$T�zg�j�v�J�t,B*��|n�$h�G����MMj���<P V|:�,*,>�u���(�Bnm`�
�tM)��w�_*:fQ0{��K��c�ڈ��u��]�gWk������֩�؛��� �o�5�]���"��Y'��¨���o8܅�ü���]�%	�5���E.�������u��E\�]zKW��ځ	�[N ���	�|�s��1m���c&��e�����*���-�&�� ��Ϧ_T��J�P����=��߉����R�����t��݃��'s�I����H��'~nWs$��Nf�����.BiH�1��M�9���(#T'�N���GtA��)]�\L�%k	[�~�t�I�QsQ�;�u͞F�1�RW6M�z(?�w���"qg?�/�"�Y0/N� Hyɓ�d��.�ȡ_�K� @�L��'H�+��MR��1GAs��d��n7ޝ�����}\7��W5m�$ȅ��Z��`P3 qP+�i%�:o:½ʵ� 2N�t� ,����	28Q���oe��ɑ�jAq�~P6{Ǔ@Y!%"đ�H�W�ٱN+Xn�L�����@�t�U1�>���pʷ����'r�i����l��m!�n����C�,�	h�в�����?|"P֚H04a�Cޘ�j:��\SĂz��2��O7e2��դ���<��X�q�c�}�.�}�a��!!J�S�t�浖��\�`k�7���V�- ǹv�RbRt����anx��'N먈J�INk._XYfY�i�y�Ɩ[����6��Բ�Jv��s��
2,ԏ����=d�2��_>��d�W���~y<�[���Z����Ū�F5�z�=�R8V�݂JxQ�c.rH�=O@�*�vc1�]x�>D�M�|����݃#��2����O����1�ړ"��bC����]��� �BU�C��Ly��7�&�1H�H�W��	@����g��9�ݙlPϪv��Ĵb������p5/���c��.L�R=���BuW,�D��w:)䱨`��l��,YeU΃n�V���'V�a�(I5���>�^I"F�n����z�ƺ�R��Vzu��/Hl`<��1e�$�&	g�Dx��(��^[������;;�,V�$��С�#�JL1�\�b7�]'YM��(f��B�7���⑟7S���`Fu�|�U��E�Cg��3ȴ�=@���p��g<��6Zm޽	���폢%�����5�U�ОK�'dV��6��ʩG�ĝ���@�P�z�3)��+e��praBH��w�gZz�(	E=%*oQ�|��^�F�w�ISC7n������Wx�Z�N���:�&�S���`�۬@��|~?�=}�]��y�@u�J��Bc#�lπ[r��+��!��C�3?�rA��E6���ACCi�ΝR�;����Ԡ�����JNb�?�E�&���[(��EMUZn�� ��wk�>Ł����׃�^�:�Pi��Oy�6��H���.pJ�ר���-'X���HFS�uYʗ6��U������PY�RY������:�^J�y������8��%`�Rf2G|e����b�a~��#m� X
b��tU��ں5���@(����� ��;��L�޲��G�r� B�C�4�zUM��6S�ދa�-T�0�����cb�/�
�h�:=��;�?~�F���h�)�}OnV<K^}�ܼ��Ƶ�(e���Ѡi��w����z^8�P�ꚺJI��E�b�oF?/TZ�ak�TK�J�zLԷ�G!�[�]|4Iƥ�� ܍�.��d��v��*i*����o��"iP�����-Z����t/��oFv�*_K Ϗ�z��D��l�V�s�7�s�Y�3����2|M�G��O'��6X��3p_k�<:���C���:�wa���_�1�C���F�a��;����v�fmV���*���Kɛ˥}�����6&��ՅG�� $��L��zK���\S��� 
%q�6���@4��?����s_o��T���=w��d����F�H�^�[�<���*'e���Y9;��v�����%����-�e�!���ڸ���849��M�fL��f�R=z��m\�{_h�^�_�T���	z��x߹��qM�A��WA�q��ɬ�s\�՚��2��XE�F��ߪ�&�h�i��L'#I��� nxc�t��9�Y6����ߒ�׻��I���^�j�+�>�AdǇ�}.�5��!><d�:�IS�[�d�9���#>��O����~�@�{��|?��ڻ2H�y��h('̿K�
d��k�;L)4�#>;�C8�������6S�P�����q�`r��`g3���c)�U�Qi��Wx:Y�m��r�7ʇ�ѩ�.%�~G�1��>�Yk�<O%��D���Ǭnj#��s��նR�NG���)f�u�y5�(��{� ���`�����i�q�Q�����¤�\k���9��P��?����0#�f����%0D��N6�?����tWT�ϩ����.��b�ϲbo�kӂXv� �� ��T�Z��� ϵǧH|Gq�us*"�$�U�lJ_!�^z>R��!��Zf��+�(��l��!SY:iwC��a?VJ�|�1 �Y��1��*�f���KX�����c�4��3}H-�E���ȖPx���Ȁ�p
�%��tQ�'3v�J괕���(u��=����.��E�Ip�t�8���hS٣.q���9��}���y���Q7�[0]K4v��O���0o�3X�c�1��ulr{9��?�Qo9w�B&PN�enKƁ�>�_eR"b1�e����p�������?R`L�M�T8h/�ò����ś�ϏQ�L�@`|���$Mx�[�o3%z~�wH�H�fZ8Y�i�w�3vʊ��3�y�X�	N��%:�27�L��ĵ̍��H6:cO�%�cL�f�]�*��:�f#�]a�d�8o�dh�A45Y3���7á lqTt�	��
��zֱ��Y>�r��:��ᴔ���k���c�{��#��W�ŧ�O"b�b�kE���?6t�W��{���\����\��z��e����O�Sg=��Bׁ��F��5��0:��Y���!����&�u�1�H06O����LaTZ�p��l�������U�&J��� ���Y��*F�'̾煼޺(_�T�������@h;1��q
��YҦ1~�j��A֊��Ӫ�<+	�f, �_ycfR3f��Q��N&����^>m$\�ElF �w�5�z�Q��V��~(����;�@l,sO�Ϣ����h	.]�$����!D��xy��kY������jg������p,pm�{�g_��u��D�p�]��~�� ����t���:7_�s&;_!�����h�\IN&����`�z7V������OOkZ��'G�n��ȑf{���q�I4��D.����&c��k%Zj���3�����Ш<�SQt�"���u��#���H�W,�)���b:�Sx*3���Jsz*ىv������!�5�!��#.���v���J��V�6N�s�np2����-���2�`���!w]��K��������J��y��
���I̕G_�`���c�w(M[<	���S��͝İOX�c�v�ğO�^�yf��TD��Qs��`D^�p�_�lft0LSb ��;^��#V�|;�G�2S�����i� j����+����6�"W�k}���@�~)�Dˍ���}��/�0����g5F4;$�>���q�("�n�,{�����T��Cz��7��I�[7"
�92=�iP	D�`�_�$U*R<�.�j�����A��Ĥjq�+uPNրE�ܔd�C� �e��\X�3��OP����|тS	-N�� ��0��(O���c,>�RP��ٯ�w҃����8�;c�n�r��/�0�'��c�F��Q�3-��]9���k����f���|O璛U�fm{�ع������3��|L� 諭��9� �7I��m|j������e#��J��������0�
������Z#B2OYz�SS�(*a&e�ޗ[W�C��5�,� W��r{9�S��~���t,�ԏa�3�҃76����-�b}P'���Y�GGBk>"�WFhzU��,����W�3q���u�����-��dZAN�"xj���C ���$k2�&[^���Zج? �JJX�����Z/W���n��b��d��n`�Oެ�ꓥ�u:Fw�XO������lL\�Ni���!���e�������_�^���^�
��j�Փ�b�I�ސ����d��28pb��ߔ2�R��{���������r�V�r"�I�H�t?�n��z�!+�8�] �f�md�oFYu��xkB�GL�� ק�#ˉ[Y(�t�-��Z:�����8�@��k�I���J��C�p�jX��'���@ S���Û I!�z�mb�ӈ�_��囿w�	jүg�\��p!t�\d���h`:8I�y�Y���,6Y�����m
IK`�����=+��.in��]�g�>�X���I���b����Z���S����I��7 ��0fZ�y@%KL�`v�%�<���0��g�S��P�����3�$$�'��E�u
��5�4C\�94���`+������J:�#{J0�d>��%]p�'~e
3�6c1ca�l޷⋚l��xX��6Ԉ�X�U����@�^Qg������ͺ�7����=f�Z�r�v�K��?m��� %�>�"&m�_ m�ya����ْV�����S,���m��\�{	H~R���P��Xȹ)Ɯ�_��W9�*ezgk�A����$��k��P�(�iynEl@�	M9��m��1'��ǃM�p�gjܜ�)i����m�\�kp�;��C燐}#i�"���c��Y?��^���C!a#A�v�jp��h�c��ǘ�!eT�ŉ�ꐚ�O�,�a����"e�F��c�`�2�W�����!��:(�|��R�a��w& ��V�:,k�����a8�LC�M��v�ǌ���{��2g���3�"���Īۧ#{jS�����rU�:���X׆��q[�[��"�#ґyˎ'Pܝ����#����&�oU�g"�O$�EEH[OH�%Gˑ����t��I�ɿj;9��=:��`�t�u��Y+�Y�$�TP2K�g1��׺�"�og_\�ς94iZ^���5/�/�?��aܡvm,3Nl/'F�!W>GI���S|�g�Ɉ�B�5�_\���͆��������~�Ur�M�e�B�j�Z���$�f!$��䳊����?lin'�%�b"��*^���(�"Cw*f*�}K�|��g��fQ�Ր9��WP���Z_l]a��n!|P ;� ���jҩ�מ�ۯ	Y8�9җW��e�D����H�J�!�W�owT�{�ضÈ @���E"�=�%#�u�X���m����=_틖ӣ�2u�c4�"a�i9��8��ڼn��,k�R���F�}$/�2j=���AwD��R���%��7�V� 
i��f �ת/���2B� Y�3�E�M�|��!��#�a�ʏ�9$��~k�tHgS�0kz�ֲ���g���]���KU�-����
�:����#�j����w<i�5�0!�SE_+��kU�Or�a��ɠ�"Pj�k%��6�d��KB��~�������z���跘C<���|'�u�pk��@uCߐ*�߿Hy0�s���9�|��W���f:���2�����f�6��"*��Cc�K ��$	I����I�Qg_��F���L���k
p|YN#p��S<�m�}���^`V4�����.��%���as� tV���s�6�1�I�l'{T�8�l#�$<���0oT%�ZH?hm�Ԁ�P�A8h*�����^G�]��z�%[�V�h��鹈�=���F���8q�V���L�h�0=S�"�����I5a��X���*;�$��7w3m%�kO�o:������p�b5�gK�[cTC"E$i�R}��LT����]��ɓ�5�+`��i�H�`��y�+D�R�Sz�4��/����j��]���,�w�p�ф�������`���Y4�(�,i%���=����\�6��s<K�Έ��GD2( /��
����R-˹/9�|OhUI�r@��1�^���xf篿^�殕ٲl��f�/E��E%guU�)J��e����^%}����S�%���ntByBܚ1[�MY~R�e��P�1���P��Y�=�K�CW�}�F�T�c�z�Y�[�ac"��]�[X��B76�$P����z6t�f_Ș~��O=��&���S���4
���~�s�E�"���SR�珹l+���P`�4�w%��aR���[
r�p�'!~���s��\\0D��ܑ��+Ʀ��O�:�u!���.�H�>,�$��2I�����$+1����)|{�u0���эd&ak�k�v��Z��IF��V�]b��:c)K
{�L�:�h�����m�?�%ebNi3�]J?8�_�L�K���hᒱ�X�;�&��<��	�g*�V�ѕ��0	r��{�T��@�#�`ҝ5X����A���Z������$��l$SG�٭I��&�$�(���I"e��1q�!P�ו��� *��N�8�#��� ks�.kdգ�5ڽ��]9hpYk��1a[ L8舖��H����n�j)�Ds�M���L���1��n�?�<�[�X�uҿ���.]ˡ>uƀB������uM*I���rT�i�v�����6l��(��\�FK2e�E�U`��P���Nb�N�Мڀ��NsF~�G$�wi��*`S5���lfOJ6q�ųi�g�¬A	A�G��{��K���z���q�h�h��h<�|Rf�I1�&_Бn�?Ճ��q��ըXM���C�<:$����A�B�Y�O-4_u��0���}����tr*#��c��(�"�u�ֽ�ƅ�PL�إ0��r?V���?-�5)�4�fUI~Z8#=ޱ}�(�U���6a�"	\_�)�e�߬�o6�̽"FE#0��9�+mUL��TrI��J�wMu��@�+Ě��P5���o��^�m�j>��"���I����?��} Y�p�S'4{�У[Gs��]h<�t!�4d�noa���P��DT1�(�M�&�����c�D��'s��4�ѕP_�el�y��{b`���l��P�3�\�S}�S�ʫʹ��+������z��(�T^��^���ɡC��Z�NP�]����L�ǜ$�\=	��y	0K��� �8qůlm<�y_�eI?As��
��S�U���Z�.3�7Yv�0���̼�S���������\������Ȉq^W�W�����������M�v�����Mɴc��6����`��r�{擳9[ S/J���:��\�U�c���0�|N*Hs?�dZ�\�E�4.n����Ko�Ơ�=K���A��K�+<1d�]�x5)���O7o���bNh�˨����w��3���"B�44Q�Z+쟚9��`�"}�&�*!9������=�3��Â��Y�W$xՄq˅#�RM�	֒��5.iM��f�����RK)������&��oC'�'G�#I�`	#��2��C�ڪP���T�璨>��?�~��&�б�8��5�Ӕ�$Jg��!��q-�:�X��Hg�D����� ���i�_ɴ3���Y8yt�gʬ���C��ͼ��!������{&����(6|��T2�����@σȾ������ڂ������پ���`���?Y_D�+�Z�
����J�?���N+��ƣ}�၌��I���|�S�q��_7v#��nVd�o�d��f�����#{;���;W��`�3}U��'�"� V�9��=E����l��L��ozK�?�ܬ�/{K����wm��öǞE2��������o���t>e��(�sFn�6�>��[��\��2F��<F{�`�|����lԹ_�.��F4�g��U��w~���O>�0�|�E��wϵN+Dn��Z�݃�߯�v��| ��K
F�����y.�1��`��+�i��$n�Ųr������x%82��2�2k�a�|{��L#
���F7�Y9����̀���>��
���ds�������k���B�@c8�zѫT�E�+��;#F��w�ߍ�-���L֎v��s����=��p�A|,ɶAXk�U\��cMjFyiePg��l���LrDˊ��#̐,>�3�ER�!<qc�5��N�/����������K���ŶV\?iL<�b�����I3���d�	�)*KHǣRg�����lS�1�RƎ�!S�p�72&�����?�� _ Rʼ��S��{D�|t��W�l!b_�D��b��kb�T��[i�q�u�
�
�U�'t&t$5(�3��٠�F��ģ�j>+'����)��KQ���D� 2n�l�	�2�3G�";!s$�I+?@Ť�!���A��#��Q&��3���r�k��]Z��"/��\#�����֎1|WlwƓ��������o�����I��N>
yr�����Br8~uЦq�Sfi�t���5X�_���*��]W��E���̚�/�!�^��O���PL�{�C�B4X���ѹ=��^��R`w���gݧ~���� �:?�p@c���3̂���0J������;GN��գ�ٖ�/wI(�{R\��y��";^��m|�9d�!d�����1���6����R�f]��mە����ɹiA�Q]X~o8������O�~�[=���QuanY�y�Մ�Y03?��+�sC��g��_�����X��\�G����r �͎X�e���L�׌��F�5�?ܠc��8OV�54�A,QO� �}��#����?�/�[*�됙T�[�޺\�ta&(d+x�z5����j"^��������~"�5И��wB�櫰Q���JAI/�o�����Iy}�A%�K6�h�q�8��'���$�aU�c6l{��ӏ\����6�φ�{�2��B��Ț���Rta���S��M#��LP��uB
���[�n�ѥ�g�.�Y�:�o�������G��3P2yޓ	��Ⱥ�g�~�o�`�H^���'�;���v\�;|s�֒����2^��D�C��W�ΗI�L�3�d�O��)�`�`!���
���t���}��d��[���o3������~�j7�E	@�\n�@Ӟ<%�$�Q�P5�R�6_�����:���
��x��9C~��]�l��ħn�6�AX���)�N��\�#ݙׂm-�h]%�"���KPqz�s֝K��a�Ӷ���_�w���i3H��0T|�C��N �-��h���ܧ�����a��_�(�jF`B��1��)Pt�
�G젖����R���j�E7
p<3/Y�G�S���Y����s��^�CI}i�A�D<gD�a��/�?ꟂZute~���l]�.X7k��p{������m��ݭT�|H%	j��bh@�<�Q�c���^�m�����,.w2��}�_���S��r�i�,�e*oJu-����4~�d/�"�0�^[���;���C�Pc_$y3�JuIFD�H��Ʌ�:G�J�p�))`�?��8����َ{~p��N�� ��3�hg�����Ӛ�[��"mm<wً]�%�<��`M�ln\�>���������D/|�_;Q)�a�/�OE��f�W�R���Zu@K����p��MЭg��h��,W��+TM�q+�[ns�!�4�]����
�?sgqI5-���ut��<�I���'�r����D�I ��_��Lyc��9������֩э�6����Ob&R��I4�4 4�KOH�`��%1��.vy��K"�H�F��HzC[Y�<�J0�{c'�����Q
��N'��~�����EMC�F�Vg:<@LF%����_�d�V�P1��2��6G�e*gt��zz�R�����A��)Szǈ�#Q���V��=�������X����8�X�����q��V|5��(�p�I�.s��r���J��2��	�������%���'��sǬV�e	o��*�}7���>���"f�=2�tx�B�&��7y����\�bs�=�
��I�+v;k.��TO����} i*s��҈2X�\���\Hs,���LT�ܦ�&!�T��o�~-д��C�9�@|���J4ђ�&�l�i�l�~��E�#:��rY_[z�:#�0���j���{�����%��b����ɞ��?�S�z�@��)YK7�+<~JbU,6V��#����:7�2s!��S�M���#�9;��6��!z��"�T�ǵ�j�L��f�8:�6֪���Y�>�����k��;
RZ��#hĒ�f.��:���7$j��x��'���=�O���*;�?@D�6w�h�f9U%*�O�B���i,p�C�����V	��NPS�6����{6(BKx_�l |i�6����� ���]u���sÇ�z/�N���xڕ)��LO�����f��fA��ob("��,7�&B܀Tbh�]IVqF���O�����h�Rb��av��@�N��k4-����	��� V��ni(�gr��/����r�jh�%u�%=o��*K��?�E_R�[+"�	f��}5�۷fXo�Z�a�3��/,V�N�l �8��)H꿷R��"9
�)%�<2װ���:�-����3cq��kp���M��{B�G����L������]B���'�˞
�v���p���|6�4���m���W�S�ӒW����\��]��һ(�3��T".^��K���=�6.�)i�5~�s�OQ ].g�&�8�����c����j���rpK���cd�^�;gp���onҹ�<��I]����N��>�?��|fws�fY�L�K�㱻������*�n��� )��E���/-��=����@K)-Xt'A���^倥�zWF7=M�`وy7�?��W�����5����B��ޝቈ@�OF�~�d%84-��n:�>�*B-UF�{�ű��ͻ�#�TeUCr����qr���4��B��'k�e(���uQ�Jr�-ck��~��/��v��<%����u�$�rЦFY�t�\t�]#�J�&f��<K���Z�&��������#V?[��^Q!�t�݉���Q��0]�3��k�E#aC<�o�%S�;&�D[_8û+һ��<���2[�?MN��%�����÷�,!��ߢ4��S�2�=�^����A.��J�o��GlxZ��i-� �C����p��)�[V����K�,ss$�h�����%���u=�G�$F.24뢣yMb�ș�l�g�n� Y`f(n�����O"��3z����ֹ�Sq�i�gxW:��YM���rg���1�����L�?����X�9��;��hgF		>ߤœ�ǁ/���O�tV��������6@�P���i�U2pp����=|Zc����3[�nn|>�|�Á�~�^;��z�r�����0͵�F�1�g���$�9�bn�� ���`8�SE��U�	�M�2������8���"�bod�&#�e�f�ދ������Ϳ[�2ZuO}���I���
6�9ٱ�ƹ�q"w��F:6&�B������%�<(1t�(Q!�i�*˵�	��ϕ�E�*; x�ץ_�)��g�w��]`eP�T�O�$�Фo�''yv�U�b�h����N�4�j�8���x�����L���,�6�����X�E��� �j���oO����2{QT�Ɩ�C�8�w���wA΀�<���b�G��j}6�Fk��������,|�������s(�� �ƇZx�����'os��	��j�����S�����pw�ֆ��Rv���&�L�*��S��gYu��ز�M~:�=dӆߚ<е&���X!i�z�R�h�$��w}봆e�ױ}�m�?[�;��C������؜��9�ʐ����~'���%���帍�8WL��)��e�S��/(V���od�~��ʺyh�O��5N;>Η�r��+�F����C"
���Os�bzp���u!R���QZ!��:.{8�@���� Lt[��a�_�hT��A]�q��K��l �Yo|]�׏G��O;�at g꠵
�� sR�N^ؙ��UJ���[�sl��W��y��Ȧ��'x��B|!)r ج���1�b:f���vu���@e9�'�%c���iФM��?"4��"㥢�=�ŴG�#����F��+��&��)��G;������<�h��hOS�#�*+�� ��gXvF֘�7hMPX�x `�.�q�i�S]�+?��R�����B��[m�i+HY2ʯ���*=S�\��^h y���e %oFH�#1aL���DCc�BZ�rs��|k�$�ډ	(MGyRI@��%hK�)��b���9C`X��`F-T�gIS����_��~�ӑs�GlW�Pzsı>C`�Ԫ���A\�u�����h-���>a:� $wc�ZF�fBa����&�rG�π��'Z���mJW��~���t��
��f&�nul�TmR���xU�uJy}!ы��f섥��!8��tpj�t���3"��ݭ. Ra��<`J�1�����P��O� ��_�P#�Z�%�q!�	\��C3��l���l�:�+ҳ���(c�xR*�G��ת�k��"��:z������+lG��4�ݤ�Р���P~ꢍ���R�ڿړ�}>����Y��O��>CzL�9Υ`],��Cw�d�k*�W>�{���V�*}��?�t@X�:=����bff�A/o��r����C6Z)��)ț�I�yLl3u��G�eB5ӱv|$Bأ淍D�X�۟��1�jR�;5Vy
F���F��/�YTM~;wx�XYG.)�z9v���m@�o��NȒ|�n0�֑��#��C�ǲ�!�����2��kX���5�����f����{\[�a5����H��.���Q	��66�f�G�,��E�H����Hl)6��/�Yj��uw�~�'l^����_�>���HJ%��,��m��[o��WQ$7_q0$DSgM��XkN!*n�~#NvJ=��$v�U%s��z�a�C�E����2dj����}����j~u'$����S��ϸs(��$,E��]�K���->e~� �Dzp�F�tů���Ѥ(F��A���_��Z�ȫ�����m�)~4T3>�eS
�z��q�w�����=�_��u�,[�3;�!�=���+��R�_�n��5�q?}/�n2 hi����T����d.^r����������$5_)������.�A���ϳm,i����ݓ��2��?��Q��.8��/�L�T�N>M�E�)�'%�Z��I	P��q�7k@m�hbV�ѳ�\��l����~�����+^\�L��1kY�\&G<�V����pŝ7�@�F<b��p�=^�p&�z��Y�pMD�q⛢N6Z���D�$������&�ZԔ�D�7nx~��q����m�6���9�'W�n��_0ZcS"߈.FUd�����saA�8�>�ks���q���b�Կ���*��*}�!�&wj�PF��GSG� ��7Q״v#::ޖui�_���kN7�N���h��,�s�L���<r���慴s9i���	+�8�Z@���K81J\x���.��d��U?�����ú�!��{x��e�t���PIi2s�_b�����N�~v���q�2��V4�e���kQ�Y�ѝ�� {ުb}֧nO���Y&-m#p�Ï����bB�-�j�)AK�=ջ����V?�C�^#�,{�kt�#��1���q�eE��\Nx'�|-q���tD2 �@���݀[�(�o��?�`�������;N�'_����@W$�������;t�-�*4�A��eH��?�e['��S����-��GC�wI�ND��ږ��V���݈��2ς��e>��3}�9XDÜMO�$=���vq�����$�rN�E^�X��d�.�Ft��o�q��0h���I��#��84-�T�Q�)�h�a˯?ҍ�<YrB��*���ʯ�w��i.�638Fc���������[h>�n˫�-��J.E�c���e��]��>��:Lϝ���^懫�pQ'�,���{�>��Z��S���}�|']�������O����G�����5r���?ٷH�"��3��zU�0�uDx������� �����&�I+��$���Ί��v/�M��z��~�����z�/�5>�Ѭ0N����8~Lb�Cu�Y�>�{G���аZ�לp}Ӿ��rJ�BR��5��NG���g���˽$�z�U;�^����'w'����x�<�ꂽ@�lF��[��y���Ҏa��7��9��#�;v~�ht��ޭ��ncQ��ѻ�O~�' f��?*r�C[�b��"Un��%4�h|��\� s�Y\�"��1w=e��٠p�;�o;�O�P	[s�~k�^u��c�Yc��#�:����	��"%ı*�6G}f��4d6%w�P��Wdɂ��a(a��'��QV����7�Y�k��憂�<��!"�P��h�@/��][��}����ֺ1��kGpM��P�N� �#FO��aW������� �W�C!^C"vr�lb�����)b��7�I[hƚ�4*�{	J�?d����p�L��`!�iˋFy�5��<��Ĉ�|�_��aW�eOtG��E
)��NH��ۻ�V>+�r߹y��u��ƪVU�xI&�兡(�My��Es�3�?�[$7.:�R���T:y{�{C�G���,,i#MC�r9uoCT%�n�=Ix@�*n�u'�0-�3���n&����C f�zz���
\z?�蔉��T������R�n�nھ�aLo��Ж���k��M(�c�%��	���D�H�\�V�͡��+%KC+�����ܒ�#3@���&�h��@Vz�׃yp~pS�n)�J�W�2��ճ4�i�%^uNx��Ud��}��Th�Jrb�J��-�m��7��� �\�?��*�˴i&����e�٦@��v� &� �ma;f)������gi���&#�y.�)�au\���cõ�^f}�H|Ap���E^p�C�X*���B���XN@�x-��/��	)�Ѝ��f޳@��R����t�S�=Q��=h���^gekjӬ?�S8���8+�znT��w2,t8$&v3c�)oe���n�Y��UY�V͎3 x��s�K;u���d���n�����������ij�k�ta�*���,C��j|,�'�A70�o��R�em�x&���@H��.���+��h_�WH�]�-&���3�#.2��v`c�����D������q�j����5"�HB�C����<�d-��S�"�$9�� Xã���)�)8�_hg�xJ�[���"��ʍ���a�� x}���:�!>�U:�jՌ ��T�y�l}���:=*�}�a��{ά@��Ż���l�/q�D��1sqO��;��:a���l�&ﮞ�pf}͘�%T�ch&��v�)	�]��:*ɒ�5�3EiQ���]�8����V3�7���v�z�"�v�^��4�[������Y��˙o��Kڠ7
ibK;����!��|3I��pB�Ek^���44���J�d{���q�;�)�'K���s��pө��&�[&��]��P��@�����x�;�.r-Q_ÐեL$�h|z����Ư����'��W@1![s��Iز�nJ��#����(J���� �j
��!���������z��:{rE�9�_t�K�/u�~m�0�Q�N��B��1%�b��`N2\��ʅ^]�y���J�x����9O~EP�a�ъ 	���k��3%2�W_�u��""ڃ�+����8k���e:`'��-L�� /���:d���op�)�r���;V��Txӹ�?���h|Ш�������Q^��u+�ͳ`��EK�R��f*&@��Vr�{5a�[�'38*���/��!k
�ګ����%ek��9h+@�_��9֠������ܴk�&�w�%G3��7�M�z�|�*�d�	D{Ȱ��pK?D�yp0�� �W������_2���9@O�n�f���"��}����y L� �hݕ�TPQN��?+7sI�?�Nqu<� �ѝ��M�9{zj
��nlڃ��R�1Ɏ��`���"oЁ���4��n����O�.*�jL�>���6qlV�t��k�L�#h����qC�������xZ��P�O������G��jQ(I�2*�+�)W�Ĝ1e6=�OH������h\���І#�*P��7�&"/>O�;��n��Ճ�WVM���S$���1���Ρ\�+����G�';4!ޛX oe��m�`a�J5�6��ܷ˖�%J�`f���/ k"-��S D�� �t��K�ؕ�.�	��;���OЙ���Ԕ��j���A��l?"����.�r�⮧�f�(6i�L�:���J|���7�2�:�{�C�^�i�2���`��md��������z
�eo'�-û��#A�Ƞb��!��$Q0�ʄ�u '���(��!��VP�݈��8<��CA��[�[~Ů�%���V8��/��ճ�`I��	�8ֆ��n��4�h�}8y�u�M/r�an�9V5���c{���& P�Y,�(�4b/�z1��0���x���u٥��8\�h2S"M	�_�iOɹ���-��;� ;��&�X�F��|�^/;�}t#�G� ��z��+m-3��5�IO���]�v𹻖��-Ik���D��.�*3���fk�2�Ւ=��ѹ��U]��R�l�.�	Qv"��hv�/���!��cp��f�/�/}��Ӥ�� bMU;�@u�( �t85��k;�����>�-���s�X�܉>f�g��}F��( �c9�:�{����7���g!l� ��?�~(���k�1�̾J�y6��Ʌp��7�d%#|`UOW�힐Zγ���Uc�S�1�j���|5wXߓ�|����~���|_��eM�E.ܗVt_��=��Ȕ����{v��JC���9�wn}��'X��S#
�5:������4.����D�K�z�2�3Q-4�����kw,Rkl*��@�v3+�6��|�x���|S��;~�@�����K�r��H�5�B#Cڜ��K��#�6�������?�gY���r�_�D5YZbG]d ��w�3�A���c���dD�q��c�z����j.��e*Nt7g1����z7?�O�H~��z�:�l1)��0�K�Ե��0>�	��!�	'OJ�fq�k�Oӽ��ܴf���0���[!�(Y�NsP�B�����Q�x`����;osVPB�7��=
��ʪ�\��T�4snZ�971eu�b��n@������P(�d���j�7��h9���������y#QdշҦ�c2\���$.0�1�M���u��S�۔^f\h�p�8�&������Ӱ�v7��hiuPx\�wQqA�������A�f��]-ZpVy���4Qvx��7�9픍!��B.�̀�?5����kWƜ��ML��>E'�7`��A�fޖ[3ׁ��% Z�Fr��õk��S�u1��j��
�R+�B��6����lUl�pu�nzN��pl_��y�(Kş�|�_饦���"�G.�5'�m�vՍE�uW��B�����3����{�]�L��oޥda�� z�M|J�P��.�ų'�V%�í���7���K���(1h��D��͚�{�=���E�T;k��:(�La,<�1j	�j��d�;��őE��Z%5cƈ�xX�� ������������_\/"7C%[�b�;c�
���-ݵ�l<T���z��r��kE�O8��Q�r9�#��c��+�[|�hÓ��|�����������w8�Ӳ�3]���̠���!9E#S�G� C��Y��ڈ�n����o#���3g���1ڤ閬���N�ˋz�pi�V���d�)4}��k>��~��rpw��0�8}R��`O$AO��f��7?�>G\:���G��� >�q����_�Bd;��U�MHj�F��$�E©��`�]L�B)Me=�Ѻ�o�q#9���
&6b�I��W�i(���0m��\7����3��I�Y��
,s��1 ��%�$�eOQh��7�'���B��oU�<�~4��W������ۃ`7�qq�!�����nL�_��9��O���!���.˓��
Z�v�[��X�J�=#��^ћu��8�2�<nK/ъו���rY�=1��.Hd_�h�Dr��8A���QD×F诔�9p%���Ս�*.�,*	ʽuC�$�U�wɂk�>�}�C��y`g&�6Z��CEY��#�M`!����"OC�ғ}T�����Ql������c�i8��`Ɋ̢��̟�"�zx�v	{f�I�mn-��#�c�D��S>��g(�~XI��[RDi���Jڽ�d�uϹto�:��?˷��Hl{!4$"ɓgh
�M���9=~�&�[����O��°�-��%H@5V?<�������w-w3qӾW����ßw_ݖS:';Ϫ;��aU
g�D���#����ga�^j�,��ia�bY�� _�`�$ojI'�KQ$CT�����p�@e/���ǿ�\��;� Jϡ��v���@K�hMx�=�*s�ͅ����g�ӬU`c���G��d��{�I3j8 �13ڤa��;P����R�b��%�_S^eʛS����i�L�V��Do��;�����I�C�x�l��5{1��-����&�mԩ�c5�ͅZCv�V�*�+��_"`���>�8�߽��r�%Kݪ�w٧ׇ��	z�v�?ph�5��	�	l=����l��	#���=���l�Q���ؗ�M�[��D���������j����Qr�/)��z5�DH�`��$�0�-B�Ɛ��є�*��2����d�J]K�I *vw:u�΄��.�u�E�NY�4�<H��D	���<�e�n�����lv�i�TU��%�j`���cz�М�,�7�Y�PD���!�lO29�^@��`�p�I3b{��v[P#�`�&fBX�<�!r�{���$�u�c�~6k�@�6B(�|���JI�c�FR��݇P$m�k����2y�8���o������|]EE��;X�rR���`%�����9<J���K?��q;���o�H���F�K��.8EK���ə������-LǊ@�������
��C��e�QN�e�i�U ���.6���@!"siZca)�&������x2�Az�NbA�>��B�J���?��8�O��c�3��/´�UZ�d!�,�_�@�o&�?h�C��#B����)P�uġ�ILé����C�Mz�I!�ǅ�)j���=��k~z��0��r0H�gCRD�V!��c��XKC��<nq�$�x�3U�m�$��̋�'o-�h����K[����D)�1�Y�����"(��˃)�ZB�s�S��rȹB2����EZ�e�sۇr��N���&�jRRƕ�Q��Qۤ�?�]&�W�댿�C��|-W���J����D94$	݂�Yo}�u�=e7Ty0�7K�tӪ=���G&U�	I�g���B[���ʛ
���2�λ����q:԰�˳��9��-T���K'$\�A�ٲW*�_L� �Һ@W8HV����ƎT���#z�B���<W���V�\���c�~F����pZ���&�!ݾ�F[J�0�
[]{��ǎ���KY��Yoq� :�O{P{�j/7��*ET���2���NՔ���
W���$4�8�\�~n-0������ՙM�4Z��*���h��SIvot��F�GT
�Q�