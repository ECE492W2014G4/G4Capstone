��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P��v�"<ߞ��&'��k%P碶�R�ӣ�sĞ������FY&����-�T��G|[�|V�=�C�<��QM�#{��}Q��l�嫂�a�n1�	C��-u)�?|��7�j� Y�1�k�
 U�����ӤR��c�&�٫-�6��w-G����Uk����/�	�sg� �$����@����ym�1|�F���I���5�g�X��Sa�A�ڴ0%�)���g%~������ǂ^!*���|Qgz��%:\=�2:e_�Oh��(p	�9;DY���*)�ь҆��$��_��olWS�6,@��	���W5�E�xT�~���U>t�ř#��.·P�m�Yhr���6���{r��y���D� ӝ+�ȼ�
�!�ي��$xub��8)kʹhg�E�ֵ)����	�{�FϙƉ�-�W@�"���[׭C��Dl��}�S�Pl����2ʵs��%�LPq}Q15�+���U��S����}_��t�M��w���iR(xw��(��r���U>����cq�ͫ�~hBvW*S����0r��J>*����t���}!-S �}ކ����u���\�� ��'�2��`��jfh���~�$�:Ģ�2�p���C�\�7�#�$�nh� nX�U}ѓ�0�Y!tҲF5@H��.����pd{E ��E�
C�+�q(����>>���}1�n?�?��&��<n���	��g�"�(�@Zf�CI��E4�����t��xY�S�R�x<♽��4݄G�qOw/�#��7��y����3��K��aʘ�-L��b:��R�>�2]e(�g����ւI5kA<G��5ޅz+)1��Dwc̵��_+�l
�}�Y���3�6h��v[�y7��H<��N�l�CĎ��
�*%��7���_?�hq�i;I4��z&�.ZY���K���6�'��b�~��ע��s�5bd?�cF�a	l���Ȯ�wYoA��Ƿ�#�M1V�ۥ����;���(A��;4�q���s96zn�?=�I�ҦF*=��ųR���κ���rZ�3F�8�K�}�F_�P�3��da��a}�$x�X&�
z/2��`�G`Co&*�y�0���:]~l��t$F�y�d�A���t��j�xm��8F/XO7�g9�7KmF����z��_�M|�&Q���S�1�^����ȅ�#|�K���Tջ��2�v�+����핼)�.��}z������x6�b���
ˍ�����"�4Ɩ:.G����L�	���UNȃs;>���rS$+gej���M��� ��I�_P�p�
������%\@CP'�gT;{�H��qů?z� � ���1����^���a,.�Z�kR�׾}�����s���[�5F��]=��8*���0J�jb��qi"d���vkr���Є�bg�db���F�D�����Ƶ�TYפ�U2~��~Y����8ak�6dr�L�y�MS��J9�j�����h���d[G�{���	���Z?��{mSr��'��ʣ�Db*��J�&sP˰��ը�������!�t�)�v\�d�s'0RJ���p઼E"������?�O�݃_E����&3���<���/�,�m�4�b���H�l(@v��cW�ā��uR��gM��u*��h'pW:���ҿ��A�t���:���?)�n�����[�i�fW(�P��lO�48+iR �U%��rS[9t�m틖Sݽ);�>��1�>���_��{۶�M��#Vm�!tf����������Q/8/h�6��ʢ�Iؽ��	p�yakX�_T��-�"<�*}�-�ouM�}��ݽ�\q_��~t/�ph����,�$�q��G�j?*s�`1
��h���A�}��U��óh��v��.�5�%2��+lb�j�hj�h,�� �BG�0�f|P�Ra��s�$2*+r\`��+�l�Vk,��|�*�����h���kw��-�?��J�Y��t�ʷ`1�<��?\O�ypM6L��`B�cj���:>��2R��*d\�H;�i�ϝ�[����,}R�D���j�7%Ѷ�(@j�����|��I��APB�����n�E,���i���2��i!J����;���rE�ޡ+m ������U�$P�g���'4�.1�y�
2�w <�w��2�<��mh%Aԭ���2��o/#����m�BJ�#�X3���vyU�~�N�2j��V�辴Ҥ��S}�w�u��:���ijB#�Ԗ�8��60��rkCˢ%���?��&ʁw*�Ϻ�g�wl��ޮd�ݳu4�Z1D�$G�m(��/�Ɯ�!�WBn�?b4P��1 �M*���|������r���p�ҁ�o�O��k�?�I���O�>��m��	QpO�s�m��q��_ᶐ�; �N��{��'�
��ս��Q]�(��P��9�|fb�#��NG�q�4�xN��ү��th;�h/5eV	8���:���Y��b+3��󀯄��s�h�=�����U��2�\�s�'�8;ώ�'D�!�1�5K����4&{ߦ	\�0��tuiڞ7�Ct+�t�4m��EQ�5���*�l��T��vG�<l��'!�#�
57"�g��SF������;h��(xЖ�E�����A�2��Z7��݄�:Ј�9	x����8�$�~��Od�W�x%d�[+i&w�>#�'V���2���� 'lnaA^BĀ5��)��� �oL1�,lF �0��rӭ��8,����Me����Q�ԍF�`Ł��n�)��v��ؕ���	u^
&�����Tf"��ӍK�u�_��O)�5c.H�?	��>�w��ή�%kW�uXB}z�u�ץt/�������T�� �1I���6��S�\�0�(�&�(i���[t�2�o�"R�x��*iI���寵��i#�=j��m�͟L�7e�Ag%2��Eo��ʐp���66sv�ԳV�ɓ����u������p%������K�]6!_5jV��:Y$Vg�dtOpީ�'�k����9$��UN7�l�G�i-(ǈ����ry���-<ӎ��a�5��L����C� ��\��2%������!�Bp�u�;@�N*�,��+������aL���~��_t<���P��'��� �:y8��vݕx"�)�-@�	a��DZb��D�t�3������޼`�L6� 5�^���YW�J�p��+$�7>�x ��?���m�2�+)���X#�L|Q���-S�����@�i�w�$�=FÃ��H�!ջ��t|���S	T�uI,����pq��F���b̲EI�>*o�>��컿�	ET�*'�{�Y�p�ߑ�F��y����CL�p\�-\�7����j��*�P]�>x|�G+)m�n�0�f�\x�p���IiU�d�Mv�$_NШT�"߶���
�ޑoj/���=	�.�9ӂ����&�X�ϭ��<���$�<�n��-�c�_�)���IJ�"/K�2��R䡶Y��" �� ٙj����^~�K""K� ��7Os������Lo�Di�K�0y��$����^	ș��s�o�J��
��Hl_z[fc�0���)�{
�=���1}
��r�ω�I��E�L��~�5�5� �CQ~5�bP���Yw���$!	�0r=��f�T�.,�����F�6���hfR��	�S��Aʈ��	���$n���Q�L��� ɺV���2�r�bN��Z��Qt��	[)����2p���Ч�Y���n���w*�HOnT�$VO���}�.P�r�a�5�[ ��ڹ�lġV�J"��Tb;MOD�%�
V�/_7��b@-/<��:4{�O�'=V��+�V�ܚ�G�b�ja��N�Zn�X.D��Z�(q����c�����qͽ������|��5�~S� �V�A���=���Z4Ԑ��m<�k�-S;�֩V�5S~�K+}b�R�gÕsH�Z�㰚�q=���Q�B��5qa+6��
#�l)��VDs����Օ{�`�C4�s+��P�{+Nv	�4� �."��� )�j�[��z�#5�Q\�j��{�B˗["$��V��*˾��<�ͼI�_��<����b0��zMڷ�]&�+�8k�r�'0�	� ���a���>��c+3-��pURV�q��:�p� ����N��jX�0���{�a�����&���y���z�{���ZG���_��N˘
�PU(I����s6;�_GX��)oUF�=M[!�PY��K�4]��nG3r����#m�M���H�wFJ�s/�a6��8���}�;q֠�+}�;�K���s`S	$4�A}�J�J�F�,G���ȔG�.'g{�UNז�YAv�Q�ڗˆ���tAa�Be����h��,���K�z�PSBZP� ���^o����a�Ǜ3��c1I6�'1eޜp��̙2�
3瓼m����џ��Z�p���t�C�lh���t�K��J���/�EJ�D8�ܤ6�x���DP�֒�A^U�=��4�;c�����Uz��1i�}2u��~M"��T��@9�/���u)xƐP4��(>��?�0���4&Vue�Ǝ#B#.��o�U[ɗ*1.OwjL=����6|���<�
u�D�&���N�DO8����7`ɰ�����.?򪓠��C@rZf����(�/y�Cه��S\LBfG�ӏ&���!��ѕ=�,��X����2�"�Da�-B1�N��
�x�b{,=~���9���증�{U� �	�ᷯAA�_��a8<�7*+��|*'s�=�F4Fa(@�&�֞f�KFv�����e�HP��VQ"�.����N�%���B�Zҽ��O�����T�扐�v~6���D�D0�i2��Yb�yxp�'������# ���k��e:~�Cn-D2�M6Ma����=�ނI����#�웆T�����ǃ���nZ��Vw�rUj�.�@;
/w]j��j�߃�'�"=W��t�jCX���_��9I����Dzުo�	Wj.$�3�=�74.��8�*Y�ӓ����a�kF�$�l�_�(��P�o��6%�l���A�rk��Zr;JS����OF���V������ݠ�R�w�����O�����m�R�G0C�X�zմ����S�`�<��w�᥿�������]�}���3q�:]��l8I. 4�Wh_Di��i*#�p;:�����ߔ@���B<{ad�N[xPA�K�4��@��7"�i�'Gw}6�L�ZQ���&����7NX� �R�7�;��^˭g�ΕQ�%RR��~L������[��u�?��c0�8����g����K�q��i�����(zd��$n$Sǻ 5�F�	4�m��O��H�P,����Tv��4ss(��7ؓ�F��&z�گ�BŹ1��O����_3�,�	;���5�&�=�_���Tx�3��C��� �������Q2yo�8ւuJ�A�@��P�'?�IJ���n@^'K/M�r23�\@ytb�KŖ
uKZ�p�Ŵ�v�M�C�8�vep�}S�aaB,�Z��p��q	��'P���C��_���ѷ�t���^�+�K;��t*����+��ɓ��s#�Ԥ�)10���Vcݔ��%y�s��-Qe����N�]<YHB���	�T��
�F�k�4}	] �0Î��K=�Hl^��#L����Yɹ�4�}@}��D��T�׸�3i:�8�XH�r�R�N>��~k�RA�D!�MB��҉
���7gQ�8B�+��趺Z.������c=BM�66��#84����&_��o����O��G����Fө;D΁�|���#o��*��
��?��(.�:�Dl*[0� �2���=���
#�2�E��4vKjb��t�|��D\�6�7�wDi��3��q4��X��9n+z$h^ڙ��x��W�<�q���3�kljB3v@� >+�C�$������$�_SG	�{�`z�	).ppBb���	r��{n #nN�U�B�7li�
Z]��_������k����2d���&���C��S�c�y�GؙE>���w*$} [A�<�Cn�ذb�a�X����h�/lA���&:��Cq��@�����B�K�k5;��'K�=!gaT�d-E��F4�Wt��w�p	�N/��A�O��|S�(4URoi�-��70:���뤚�Lfbt���vq
���AM��;�z�����M�n$�M7�OC�����Z�N�E��'c�z�����-"��NNWl�� �b��w�k~��-��2\r�b� � �u�y-��dn�kv..'�E�Dnv�)���0��
�i��������=���m����^��MQ�$I���}�����67������ b��$�^`���� ߻Vx��,i�A�j��Α��u��+��!
�H��s&��Qv�8,M��b��K�KD��1C!2��%"FF����#U!C�%QH�2C{A6 s��㏴8���.�5�\(W�����a�䋗�����ӑ��,��}�SM0~gtD��pE ��e(6$��'�[Þ?`�|�$>�Lx�"�#:)�3��N��{4��a���@v��Q�EBBս.�,+�#��S�q;2��a;.���IY��L�>�zK1�7�᭵��M�7��iKv���9��ěF�L��=�dq���z׈���2���V��Q�rx�k��rZ���_X��dh���~�ϸ������X*��13ﻪ^U܀I����d���Z�+�Ӛ9�~mcz�_��و+��\����^�&�>�\��X��z�⨜�n��/��H;�,�3]��69	y�4�jp6dU
��kky�̷����������p�aQL�3^��x�cN�0>�ǓAǡ�o�����TЧ��"�J��s�!��@4"^ƙp���Ԇ�F����y��\��������Ǉ�Jy�J�MB�4ԅ<�.x�Ԃ�Q��괜)�Ɋ��a?#&����1\Њ�&�:�����p��z�M ��A�g�{����?�i��6�ͯi+���<nE0S:;ԃ
.1WTs����|E��.y��$�lB�SU�ڄ��� K�.5l/Ԫ؞�Ӭ=k��f����L���Zot��:�*�)R�Ų�n����Z4kv�2]S���:�ݖq��N�<�	U��`_�
��5z'�����h�#�?�B���kP0����!,G�����m��N?]ٟ� I!��_����:���ބy��Q��T����B�H��E?뚘�-\y~���aY�D��p>�IUm�q�(�
�ы5q��	��赆g8B�U���eE&��)&�8ލ-��x�rqF����ud�e:5/m�:�[��@��+:�ێh�a�;mXB�z��(\���,+LYD�ut�҃�/�RBQʼ��`�m�����g	8�U�a���.h��"n�ӧsw���7f�{j�If���N ����r�`�4r��n�Q7�k,R)�Nq؇�BⱳK	���|뢿×@]�[�z�9-�p����XzS������	��#;cdm���yk��?��K9�^�r�ij�Vlo�L~�t7^�b���nE�섪�YKwȭo�;�K���y��5˥���tܰt�R��������.��=��[��+�)����&	l���{%Hq��
ha�_�'�+)a���2^���R���9�r�#�$���~YL���I=dz*���� }Y`M;��j�u�+���sV{?�#u5T[���	���:����{$w2ƪ}�c�2>���b.=�D$Gކ�,�����*��g��*�cJ�e�}A����ɧ�~"�;X�2��6�%>����C�����,k��p�Ĩ��F�$�ю���-����dv*�`8F��#��tz@3˲:�禖�!�ܙA]��� ���|�n#؞cv
l���
W@�W�a`�eU��$	e�	<2A���������+�$K�,J�fM��b[�W��x���M���Y:Wk��v�Dݩy��ľ�셪F*�_Y'�	���ߓ��b�J��]�F�yc�^�H8&�`�Z[�n�&'T�(�͈��z���i]?� >ߒ��"�Ϭ'UH$�Wi�אb�8�Z�nQ�:6���t�����su���G!�p.��WH]ya�üQ� ǝ��>��Qwa6�jށ�O��H���:�^7~E���*jw-�5�ea���� *�w�K��h)�?MH��H4؎��Y~cY`N��  �D�^pj�^�Һ����N,�l���q	�ƍ`��
P�P��oC[�ػ�Y����`#���2<`C��'��]f+\����ݺ�S��=k��Ui֘���\�Rh�xY��%ik�
�px+�icb����������A[J9�����L�.��%9��!
^*�7��`e��uӔ��o���� 8��cՂ���G� t�����7�@J{�)����A6��P����o'�����2�ɳb�9�qE����!R)t�q�ƞ�i�w���������܈i�&0)~f���`#=�h��ƇЃQf�<|L�o��s�.P�e����� G�f	tu����S�ݚ^4��D f�R.�#�ʾ�PK�F����M��+���ƞ$=�bۘ̌�{��}2(�F�f�Vll-�m���5���7���8��z�ӕ+fVx��ư��g��H�[U �~�.m==���sx��0�_��ĺ��@��3<&r ���z�ѡ��ب�3,��sI3s�-�{����J��!�sZ۾\��	c͡�|�&���$���˰S፯�wv~3p҆nd�
qn��ج-�b��J�4�n"$]Ş�<20�Ʊo�ܽf���1��W�I�6B�G��ݩ�:Df뺄�)�v\Q���$Y�� �M�B�W��g����{�A�#%��K�_ ����VEՈ.��ɽ��T���'6���j��ہ*>ʌt�櫌����f"��@wOů`6�WA��R� R�q�3L)�t��#7��m�rE
�)�(z\��q̿7/��e��A5�Q"���@M�`����C�*J�(�v����01-Y������M��^�~��Ǻ(��Z�m@\oྜྷ��ٞ�Aőtz�!�2����C�W�䊭bNP���~P�(-^��~��p$����[�S�S�
:�I�'L�UD��®�*�/�"����M�I]��!]}3{��%h��X',�m�/�
[�`�K��X��g�*��Z�C��=�j
QX��ov�ˮD@4��%�d�k�PD��$_��Um�A\d��=�r�sdF�g����
����:h�oV�T�������Y*�nT�%�y:c��t1�w�$�� �.��ҟ�uq�	uރ��*�na�x�O�O��e<���(Ӆ�>��U܎��/��զp���14��t�r��B�(f�g���q�T1�/�W����@�
����3�`�&���v�1���d���yHXu`�r�r�cPY�}hg���dSX�l�}Ә��I�H���L2��L.'Ϲ�́�j�(���B�|@���m�Cΐ`7�۹�A�Q9q};L���TmNx��q�W���6-��#�E�x�>� {R*�Ä	�"�-�]�O��z��ӳ��>����=±�o|��H	�;��&)ئ��Έ,D�F�t��־(�1a�M
*����#.5[3\Y�y/�G��Z��n�l�?���6ҽ��䕦:I��"eb%Y�@��TGꗦ� ��ѽ`*�ZXh��`n|7�~�����2��+(`r�S!Uf�C�Vi:񡬣��a�=>7��ݓ�G=�|�ؐ��6V�Q���C�@��7 �Dh,����O���gfm|2�"'�
R;���1Ap���Kgf:�����x��'}�T����t)̈́��&+�JX	��t��G����x��i���G����~��Kh��-�df8H� !�>���w�Gg�j�7m�2�e�^m�{EqUl+Lg����/쐡���Qa����W���o'��k(���4�NHB�ӧ�?պ�gt�XR�˒��Oz�Κ-�&E&!6�=��0�p�n����9��n��S��JL��Q�~@�l���ũLLt(�?;M�`�ْ1��n%S�["���t�g(��.��)LN��!ic�j&y�)��r���I���9�v����X�!����ijU��3�ڿ��BC��B<��	�����%Ec�6c"*4�dC& ^EMȓ�y�׼�rG�JI��0^Y��"T��p���'��2"��Q5�Nl����Cџ��b��s�r�^Va�B�92t�/<��QD2K@j��	�`8�b��Pl��.�����r�Q��(���]\���]�v]�!�e����T��P,� qb����i�;m6^	�e�����4�.��IB��s|���ٷt�ً���V�O0�Η%���tPx��<�� e{���k�=i��s�d�v�&=/���"D��_^^�C�W��/��i�|����G��^���|�[���j�4º�Q���."��N��	
���Y.���I�!=�:��03!'�O�Vq�e����T�Ksgn�_�����A�OG7#�{ӓ�肪B���N3(�����kQ�@Z}���Gx��f��l6�J�HUWꌘt�3�4���>��@��[�tq��Pa:αׄ��� �B�IՔ'�9[jiٹnj]�3CԀ�1F��Hp��F����C�ý�a�s}r(Q�6d�,f�x>�� �hz�� /)�/[p��ف2��&鏈:*�b��ʴq�S�&�m'�
���e'I���TIݝ��̐C��Y�l�#�R�Aov��l�?'ɋ��Сzd�����l���zĬ�[��ƫ���H����� Rt�@�ѳ��m#<K�M��Ql�/��U���`���d4M��<���>�4��R9����ɲEQ�����x�!�Z�_�n�R�[���%��<G�����%c~Z��9��%1�~s�?I?&c%���/"颯W�H#`K��ߧl��7�B���qRq��Ȟ�V<�4_�*���`�z��֜iQ�����i�<Z&[<��E!���ٿR�q~���.�A�G�%c�pt���N��\d)�'�h�7],7i0�����z��Ѭbd))�;��&g8�履t�5<��"k�S~�l�S��q�����#�CjXb,5:��va5H�O>����|2�^<�X?�7�,f7zf(YU� f"@��Ѕt�X:ami�{J˨�HB?4>�HW�:/n��*w�U�0>p]�4#�L�3���}s㲻ZM����GVV]P�����<�RM~�䤙 �z.-]�/l���~dD�?[�0������'`��_Oi�����d��dB�áV��>����#��D^��F�-B��� �NY�"�&�͇�˯&���%<�8��>J���(:�r�������횁��X!�۬��U-�/��X�B`�����-������X�R����s�=CF	'���|�B�Ԑ��B�Ԝ�+o�