��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P��v�"<ߞ��&'��k%P碶�R�ӣ�sĞ������FY&-揍�2� $N�0)Q�Nr?@[�|�~��,����Z����u�){�.��r���zi�f
�|�,*������o�/�AE#�7�?�/��6��[��Բq��@x���f~`��ՙc� |�h �S�u�N�Rd����(?�Vw��k���i$���QG���w`@E߷��H�j���y8ύn�͢���o�s�����V�P��¯��' 1)Ĕs�@ �/���'D8j�_SSG}���u���P]S���T���-� h�/��ʩ_���_�T,�<�#�Cj%h�|!�HG\��3H:��%���K�����Q����D�,,����ߞ��~h�5Y�u݅%�/п�P����epؐ��L�����cr�Q�;��j�Ћ`?��fD�)�(���v�X8xruv�P5�զ�8F��L?���5AW��Je��I��[��-{j;�=�f�V/�9�2�MpK�8-3bTkW�p|Mh6I��Y�[�J��i�=v3�1���I��G���+�=�����yH�g��щ\V�۳�D������z�
�ȿ�d�F_6e_q��q�J{e�
�.�Ky�.�� ��V6��+���)V\:$�;��7v��j�5�OK�וj�BEO~ƫ��2d�	�砳4��e̩�(�PL�G���$DvƬ��&����5�L'DR7����\�n��l/Qaa�>cu��q,��..l���0J�0��i`z�l����21O^��/��W*�o�k�������1�"d�֢�׿�86O���Z}\�#�k�eOejU�����RL�0:�!Q	n�)l�[�;=�;K�:��ig��Qs���\n�H��p��]�M���F�b]U%�U���"_)[���a�Qs&�A���6�A?��qhDȁx� D������yƑb���t��y����~
��j$�����6�בzF��^z������j1�:,.E�����~�3��c���\�²n.��M���)�<y`0k(�]�P1�|�c���6٫*��{MoM���ԫ!�c�훍�������q�0c9�����c{����3��A��~T�Z�=a�?��6R�V��3��յ¹�%2]܎��\�.WN��`<U��>e�3F	�W�n�z�[�i�p����m��x�=x�kCe/sY�d��bh�O���i�1j�m02��67�紉]t����`�ĕ.}d���9BQjLN8��i�Ӊ��'|m �2�A$�#��0,3�׮H(�~�>�l��8W�>��d�ƖL2|��3ړ�� L[hk?���w��5Gsz���M�}��.�
*��gP���M{�&�H���C���� �<!@ �w<�	uT$^X#�BL=4w�=����Ԯ�U?KV������ ���[c2�`��"օ���I�v
ۚ�z�ݜ�p�({�B��6.y�I�nuK���N�� d�h	^a�e����3$� M������tx��c��<�(O��U3���uW��w���as��4"��9y=%�owa�}���o[�VU����(�&�z6G�h�{h[lo��+�=�3�7�W%[�'˭*\�T(��=<eǢf�R�rd���Y�Ut� `>Du�K�c�n6��W���X�%���*��U��h�܎����6��ѻ�:wP�:+����@0�`?����4T`��dѬ��eK���F��G��%��d6UU^��:���Y�*�`~_gq��Pl�p�Z%)��nR;/���{b8]1�܋�SF��~�@(���YaÉ/��RKD����"�]�b9�ӛh�_	3�'{�!Y�9>'V�� A�T���j�F8���/��QܦD]W-C��րiF�ˀ��LF^�� m�.R�H��К{��%��ŢQmZsq��3�{����H��}���SKG,���et�#�VF�7T%~k���n�sc0���B�9�
!�1��b�Z�N6�#���dPZLw5�����-� 7Z6�e�9�s��$k���u,��p���^�#��,�2]*��/�?�~
I�bv7������-��+G�kO��Pg�H�Q�ɥ��d�:�����yx���<�$����������#�s��M"0uP|ڷ�+(����rO��E��e8'�)j���Z�؏�{FT"z�����qU���������%p�oG��}Q�����E��	�*j�M����-4��8��<��[�hT(ݮ��#,����?ō�[xtm(�'0~���6�~�xj&�n����+������N ��#�6rڥ1���-��(���C�?4��緳�tS����īi���jo_��s�¶Д�{ �&cŶL� �0<
��QE[(<ݨ�2@��~��t�=�-A��˺w�����e$�6I�������jo.��YС���� ��j���	�!�NF�;��וO4�њ�kC(��kc*�9O�g:���n�j�_�0���`�M8��}���tu�M!Q���4��#�=QV�N�)�~��_o����8�D�N Fw�-�U���ǽ�@РxhǾR�fb��S��F6�N�(vI�!���F�1��ʳ��=no.����׫2���1�T��Pc=��N�)xC[��i���9�R�Q��9�f�2Y^��܇:�U&t!����JK����g~��H��)��߼M3�n���0RD37�_�Q]3��T��6ƞ��2��l�*~`�����$��[��I�6���2?@��Q��$`̟
�yh����Y�j�P�T��~�z��sa��^�Ejr#BewN������6����6L]�a��H�IqK.a*���$���^���T4���ݸ�����n�;S�X+Ώ��[�0|>7�]���{>ymǥ��]���py�[���>.����:��d3w�Ӵ���Z��5L�4�t�'ʑ� �:S:O䞨�r�
���,E�~��4�	\�NS��Xk��Q�iͨ/՘14��D�,�UKjj�l ~��hL+�-��ö��s���\-zOz�'��\���<ID��H)Vq���d�!C`1����n؀�b�A�g�	C.�qkc4�kQ��JQ�[��gJ�o�L�w���kVdWU��3�9>jK�����O�c�)�+�e� ���"ʬ��l��.�$�q�@��,�����B����6�7l&+2����y���C�`�^\�T�P�9:?�O$Vj��]������|Ȼ��4w��D��'������l�x��6�:���(�e%Y��<�y��u�8��LA�27?a��p�#�%�).��λ}���g���N�r�!��ZyD�u>Y��K���;���Mm�d@�±	2<��� ��ڹz��F#�;��<]z?MD_W⺎[�O䯪+&ӳlE�鿔���s�C}�CN,吝F,>��6C#Q:�㴯���l��/�m}����&�����A����	i5YKo2�Z���[��y��yr.{��9�%�h���R��'��&A�Xo�1�Lu�.~��&�R�!�^���szm��y_�Xu��?��y�/����w���O-`ؼ�vu+�(�T5٩�;���j×%� �3��B��O{gy�TV�.�f�tv�%U���v����1�� �[Q��/�D6�V��@�b4W� �*ꞤL���v�>��R>���h��|��z�0�1^=}�,��LQ��������%�8{W_Ц^LQd��u�Ä ��A��{�Vc.�Vj:u�a�&���q+��h�,�3|�@;�3�X��L�T`��UG)Hv��c�pc����vLU��<H�r�2P�踲e�t��[�PE�f4+N��C�v�iw3�$
�Ѧ͵�jWO<N�eH��&��H��!YG^֨3�c���1RHX߻�Z�fh|)7[�L��� ���+�_�U�_d��o��3��Iq����X�-��y�Z2Z��x���֯~�#".�(�BsO����;��޳��$\�������+<�;Z�j?da=�TDTLf��'����E�,�l>�d`EBƈ�d�d�ܱ�7o)�Mn|-+<&��>��#��n[�8�`�oZ���ÔP��w��D���y���R`�iݴw�d���i+X)�	C7J����&��\�/	8�Df!'�X����XYe@�O�Y�2Mq���{2vQ�I��nζC�	N�qQOf���F\�F�X�\��4�L�yl�l~o�P�g��8K�~Qcs���c�H�� M�4a=u����i�#�
����&/��0��+�N�f{l��tS@2�0]�*��5Y�]��@�k�b]3���墂��ک�n��w#��"K}ڻ����h
!��
��%�~�-�[,�!�=$�8�8m{�
�y�[��E���N��)b�ĕ�W#V]��14��E�{M}_s:�\�a-�NC2�&ơ��Yқ��DV����_~)�	|��;��c��KP's�{�J^Bێ)J�[�G��L��=��YFAx�_�|���H^��3^;�Q��E9�L6��X�zN�:��6o�!z��֝��<��$��X��_j<fx:�����Lķ�T�C�q���+5���1�,�ʾ>6 O�k�cΰV�CCT��i�=m=�����!����'0���ȫ�'%3�#KL}��v�{ GpQ��kb3%>!Sx��-�s"�a�U<9��Hj��@���]�lBt�\�H���b�V�Z[�x��#`|�kA�x����}�Ikb�Z3�6�������!-	�>6�d*�c�V�wzut���X�8��vJSj�d��@��n;��uyA� ��<���e{�XAs���J��=F��6�K�}������hspPl,���W�k��=<��ۚG6g`���ז�B��ౡr)���������yKː=R����>>wm��5��f������$=̟�
ϭ��}^v$�}&4,�*������fηf�w�k�f��v��]VAtt�CZ�eC1�v�8ya(L��c����� �$ծ�Iܢ��N�.��K��S���/�vO�ZE�I�\&R�Q��un��T�jij%�z%���.�x>�g���
����^�ű����P��8q�v@~��SJ-T�����-��y6�$Ҷ��b���3=��	V���@:4�C]��*S���RJ`M�b	ut�J�v-{��`,�O e<�8i�V. a0���xj�r��sKl$	�Ȇ�)dͤh�_���'���^g���j�����t�V����Q�t��#A��;�`)kB#�Ujf�D��t'p+���[S��)�T����ތi��P�!P��1MY�U���W@�J��ۿ��_�ϐq�;_­�dϚػ8� ֒l�������V�2~��~�:5?�ܓ4~��&�Ĕ+��5/X�}V}S�n�0���H==U���3�Fs��CuA'���MeS���Q�
�Z�]k�,7���}#Y�����5Z��;�2��FCȕ>��D6����j���8��{!3��{2�.�=v��ah�T�Y�qn���_q�BEE��K�2���af+�R�� ^�{�~��y@�.�l��3>	�9?Яׅ��Y����k��r˰�q�� ���"�g�"ϓNv�̉�֮�-�`�\c�VAylB���z���^=��1��Cr�S���'���%B�(���y���͹?��>N4��mxiAc5l��|�]RY��2x�I�k[�W��i���|ხ��e1[?�O��%����^Ŀw	+?�z	�du��/����=������e��#]��)��5S�D�l�!�ho�bjsF[m�ˢ*x�W���F/�$g��٩�b)�*���a��K�Pn��rG�W�o�.��� ���[�����
�\��2b����v�ז�7�c��K%lCd[Bӳ~զ�?	Œ�&����-�w�;젔�?.ϘRD�	��7���ӛ-�E�WqTZU��6��i��]��]�{P��������.�z��В��[Y8��X	c�$Q�E�e��m�r��%�V��>�z�t1~t�Ԩ}�?���h�M��0�w!�:��.f�;=f)7�c>F0N����#\���
����\.A��)�5����9��P&��w�I��Q�q�S�7_�䲒o��)�A԰>!.Ms&�t�`���MgLQf٤bKN	�,Mq�x��]��^�_n��!l��>H��"��7�O�gj�����){�ꪍ�YDz�{m��6������6_?���MG�g�i�bVH�����NZ8�?�Mi�r([�|c����\���i1�fi�#����o΢�ޟ��Ò�n�I�|�f����2Vy�[�P���I"�u�l��뭓ȏ��]�s�!\�T�z�ѓ��o\����eO.J$�|�"y%g��tUqp�P�K��Ȟ���[(3��{v��llg*��`d Ө���!��P�h����4��8O|�L|��q[��#��1\6��*ߒ���x`c�@�1�:P<E����L?����n�Z��)E�m��f�f��4X��2�v����{Wt���æ���.7�[
U�:p;�5��k`��.����~.�"��;��i�]Ij~���ˠ���ͥ��&��gYdI0th�oE� jn����/�N�!�#O�^<��z`��
qlC2x��(!�FI"���H-���{����E1�����'|����Q֩�RŽ���(F&iZ�	%�����<Eo���&����Wf")���5��/����w�"�#�d2_����ƚ���y*�re����'� ���e���@Qy6'ʋ-�D��[�z�𲓪L��ui<-�Јs�9���%6�,�"i����|��#�oa�Jy^��d��Ĭ�u
	;��@��-����4� �X�V�{�0��'yyX)q����f|pġ=my�����U��k�&Z9����B^y��]l���5-a��.(� �I�#(�����S�b�K�@=��V��"Y�>��(V��#ҫ���ݼ�>Q�s)V�y��{�Џ�0��C�Tm�ү��fd�mB�.��k�.P*�����.�.k~+t�R
ioe�6�~��F:z!-+��b�K�'�ry���-���A�ZGmC�۾��򗛿]H��I�aeqLǺڼ���È�z�ҳ��e:�s�AL�Z%�~��''��y���攣�$v�K��e�$$��'��^�md��\X�����M��vAV(�ix���=�=�k���!�"��E��$�Z��jS�:��ѻ1��U�D-��|�;�s#$?��p���`t5X�J�y͙)e�D���{UCx�ъ<1?�}�
P�j�]v��Y�`Z�Ę/6�+�q=����H��%��ƃ	(�{
VE�ik>2��»e��������X��v��oj�=K>���Q�*�olg�	����G7f�E�[�[$:��z1<�ܿ�����g�~���H���~QOS��[�s� ë6���7<���N4vNme�\/F��?���|#&)tu0<���|��S���`k�Hlng�\�CD"]G7n_n�!��0E�������$Sh��'��{������D��jd�;f�Z�&��[Ab�Z���G58c*�NV���D�Qy/��꒬�2u�V�m�t&j�?��^HyT5ٙ��[�cc���q��+,1�돢Dmi����F�:�3�?��2^��Ȼ�2��m�7��-����1�!�t�o�e5�bO ��)��f��3M~KN�y��$�@�1v�KQ��]�F�	���(�ǉ͏F!�a�)̛u��~�ms��CQ�x` �<�s��~m�&}����B!�;���I���c6S�ꄮ.�sD�ƛ�cY�6�=��&��a��,l��ݦd m��`�o�F�h'"���`��Qn�-vr���2a@�w��и�� �k\p<��U\O����w��* w?h��OY��f���4��Po��Ű{��a\3K�uE�'�;���m��7-��O~�VȚ��x���0~_u�{8��	m���;#�~	j�#�y >��'�4N-x�l��e)�^���B�H�C�		г'D�/S�"5L��[嫕%�|DJ��&�igi?�o�׷2vF�����	>G�`󷝕��B[I,��M{���f�����m� ��8����q<h#�ۏ{��Y5K!�l6�u��C�p��d�!Y��s�壏O1��r`9�5lE}1�E1���H���ш���6h+5mQ���#���&�pk�KS��C�8ȅ�O��3��y��4��%}���yk/�-6myYN���5����jur(Q�j�q.]��kZ%��z����sNզ������콨�[���O7�44�^��q;O�K�6��9����/I���&�mjRY�J�[��������/�O�ɝA����.E%��/^ط�LD+�أ���g���p8����_�(�T<��YFeJ�I[���[q�j]��P)�,�[Ѧ휮}���'������T�3<ʹ\7�b5�yD ��)���g (Qi�RB�S�����	v � \���9��,v��9��?N)��]OI*�����Ҕ�L�8>�~`���?�C��1�� l%_�t���M��0]<�������H����#�/N�4f4�������)����р�fF�-r�/
L�%�{A��d�_� >>P&>7X��`^/�>�;JG7d�mi�CU� �t��h�>�PL��-	�8PO_�j%�;��6w%�i����
�"�W%�yBŀ�,^D]��
<>~�7�@�9o-�<�$=Rb�g���v�����f��Qj����|�z`�G������E�j�6M2" ?��$⊚)��}u.��/�a�F,�Q�����q�j{+���ș��d�dq����k�n�,눃��X�����\����:P'Ūqɻ���n�\p$��J��o����}��c��namO��ܻ�^dZ��I�hb{��GJ���2M�ϕad�����tw��QhNE��Tf�a�QW�(7�gp��m���l��w�Q���p3���~�[�������BHҮ`(����[�CF�Eh�3%�*!d�wz��м6Sc�^�g�
*5d�6����F�"��d�A����a��朼���GU�*蘷�+¾>�b�p����R�ɤ������rB_־,D����2�:�9���Mɟe,�l�[�+�Z�S�����b+����0��͎���%`ѻ����ȸ�����]���������=Q\F���t�LCH)��L�K#+���^�����R��E@��R91�p���k�����[lW]���#=�-$]D,%���H{�(�����=g��w11�RL����H�c�CT�����9O���W�H��0|��X hR���I�YA!���v]:B��n9��a�Kp�C�=M���M�>�qHdЅ/�����Ȥg��B2lź��Q���g���!n��ɢ�KX��ZyD�q�6׹��CSc������av��x3�}�)��g�f_���9 ��Z�7:l�M�Ô%���͹�G�ߪ:�g.��&��=�&����\V���Aco�f���WPJm�Cp�ݣ޽a�?���d9�j�}�dDS��nN�2��� _f�ʆ�(S���b�P��� X�{T%��pQ���=�ޕ2��P��廙������@{k<�{�oI�k�D�D抢52I9v�N�a��V,��+�q����7�Yǖ�)sj0��V��U�Rj==�u����XNq�*�۠S&�o��K�ݧ�|��bq�M�<�l����v��=ď]��ö]�}PM�P���e��.��=^>����6K���=F����P7��?�MΤ�A��cR���{�b��X�1��zǧL�	��[tJ
ݕ������o�{)�E��uMF��%�c~�N���~q��	�*s��p���3��@k��Vj��������wB`[���S���\vC���N��d�g|(��	�I$(  �����������8%���va���U^�
�u++YR��	"���WE];��ܹ��,H
0@��W�^���W�R9�$�D>����U��F���Y��L�Kֿ�Zc�WwYZJvL*!ϕ���o�L�ջ#����X[OL�$�����l!�#(�[�r�k���f��?tOv���I��Q�h:u(u�V6�#�@��w�~����p�SjB���E]p�x4l��j�*yՒ��Pd���Y�ԏ�C�q4�1,�:�K��[cZ]�l/��s���9�1ZZ^��UGa���Jk:�̆(t/m��*�?X��w����9�7�`��`�iS�e@�K�)�N�Mpςj�|h�y�jW|ZŃH�-!�ڀ��`�R��E&J�IG }bƇRШ��@�0���J�n��c�)z�SKo^qB�.�pwvp|~�E3���LP0+���OKA*?Nu��'u�ȏ����3�)��K,D��R�ܢ�"��dM�j���;jf��K�!�gT�N��/Q�ע�_W�u�~����#u}��Td���,��(l�h����TҪ�kr�)`�G#��ŧe���,A��=�@x8l����k������+��q�O���G�>��O_����3�T	��@t����]�"��g9sIa��<� �^C�ޥd���V���Фq,/bk�]�C�2 3vM���� ��[��(O�LTG����m��DYb�v,^/X]�"Z��=�"�?a�Ż��P���[�"��ǻvs���doA��� ��aZl���n�� 4��]_#�������
���8�c- �8K]%��-\��UA��yc�v����#��N��E��i�o֖�곧��1")4=n.Q�`Y]0��V�0�M�dW ԇT)�Y�❛�%~�< )�h0X��XGu_ [c�Y�!_����`�p1cն@m�[,�M���9Q���`���>�A(�Fn���X5}1��ol#i����W��礂�$�#�@*$���A�cݠq ���2�n�R �K��u��1�U�#Uj$o/�E��e�({r�­�yވ[�ks����@a$l��`����_%A�J����H9-�O:*a��Â�~�VIk����*��|,V*���y�
�`�$`�x]����GQ�?����X7N'B��
�'���֌��[9��;��n�q�tD7R�	�()K2��xc>�C�>����F��x���T�:�8e�8��l��I\ǲ����^$C$f�����fa�����[0�qN�teV&۹�:'Vz����+1%��R�G3�:���o�h:����N��uH/`P>�UM�v�l�6k�s�j7c�{�f}�Z|�D�&ۗ�ؖ����,�9��2甞��48s�M`MP�t!CK��4G����<�.t���_D�ՕQ�=uٞ~�Vs��x���5~��`@O}Ę���|��{��U���'>\p�,h��l�l�zD> 6�e"ջ��ɥ��jm�0�T��ӹ�fS�q�����������ۉ��W���J �/z�~h�x�VO��f��@=J��`([�b�f�����90�S���m�ӏ��@��dP�*�M�Ĕ��Ub{P���h�F:nW�i�wY���d7�s��@?�%|�w,�iy��|�7�m7��KZX���4Hb,r�[=bۊ�$I`�-F���_����FH��t$4����y�UC(C�E�ů*4��/�0��l�-~J���B�����i9�M٬�ml�T�t�y�����;�D��v��N��3m�/t��OӴ�u��y�H���upo,�P���)יִH��H,p��b���� '.m
 9"����+�|8��9�[jK-5\I�/�i��5�PI�����呶�H���"�=�+F��a��[{�<�s�r��S��N�X'�;1g��|�Tf1�Ud�)E����u��q�mCq�����:f�x�k�vH���+�(v���s�^�$�!V�6Cg!^��f)����(��������dԴџwx�dh��BG�{-��uy`P�	ݙϠ^O<�-X���]�a(�]�ߪ��!2u����8�#ʱ�^�ν�rc$�w��֯��0&!�t��*z`D����}Q�!\v�o�WZ�������.z��
������,�%�:�4�o3��"�W�]QIq�e���v���,��/�D�O�e�~�M��y�Q�e��\9���n�*f�5������z���M�el�ם�7�g6�BM��\��&]��V*�A>A?4De��:
��9��,�_�|Y���[�����Ǝ�K
�l���5����Gm�c���9�+�R��;n���_���
������C�`�7�1�Gi��S�w�n�������z��N�{��ڑĥ#�����֒T��ED	s��q��P[͆z8	��!���|o�{�����K��/Z�����"+.��
��0�V�8'��^�tAi0=h{u�#Aj!��J�c�q��=g�~��Q+#>b6�<�h��-f C��_j�^Ox��A��롧Q{�jhߤu:��`��6���b	�5�8�.߰n>X�����F����F}�{ƶ
��!�(�<gz���}�p�� �"/��#\�f�����>5Q����Kr��i�S�^R���dlѭ���S�Ե�j^Au�� ]\�ρ��qd�(<�,P��K��>��-0��K���7e�tEw��Ң3�?�USE�����
9��#P�}x