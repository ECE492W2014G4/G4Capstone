��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>��`HX����5a8Sjf��4Oᐢ��\���s���(���T��p򱯋��}�w�i�|�typ)4�eV߁�����o9�␬+$����lY0��S�6�ڪ�<�]�Wų���2�:wh�GHFN���Ҩ�*CC�`�CJV���py P�{Z�����a� �w��������V���ѠH���C�Hp��K�l�)X
�<��#�����ð,�N�����ק�H�����H =���O���H�'N�� <�\"�dɟɯr���ORh��@�-�>Qү*�I,�h��9tE��-`�ɰ�ɐ��j�����0B�2�^������+a7�z��x8p}�S�G^�C�C����,XL�ݨfo��!k��%
�`�Iq=jh AF���ϩ��]M���k�����2���D@I�Az�������IO8���{��w��|�;F�<df)�|��s�ʯ�IP�F���Nzq$0h��M`L��b�$7�:b��&i��}H��cWw&���xD��#g�,kz,������q�[�|�� �H�;������Xe��LԹl��	>���Y�TD��v�@�ޟd���ω&��f�81����-/���_v�����T���l}+O����6Xٲ���~��@�PUb�[(��g�Fv�b+�ρ���Ӓ�r��Z�Sҿ�O��>Z�H ������KI�jna�����E����@�I�%DF������W$�(~��`�{"m���4�_�oF����2T0�zG��3�rv�������i>7��_uVQʇ�(�G|IaB�Z{���F�u��|?���{�*{��oǉ��C��B��7��G�@^�P��bRl�"l[�zW�B8/�`�����Bh�l�Qy�����9�y'(&]�A��t�Hp l;Mֱ%k�Fڴt�;�	Ӹ�dc-��Yu��GϠ�U]Tz�	0��7���2&�8��騍��R�H���l����᝵S�$0�q�w��)�g�W�QG*%���4܊�I8��nb7*��TC�:�_n��d�b���%��`)$�/oN���.d�d,���#@f�Z֭��'�ڂ�A���ZNV�������<M��������������@|q�� ݝ0�\��ԯ/��<��݅`��1�B���c��1I�0�+��`�K���/����#w�������/"�4�C=ѳp󈯫`�w�d��!H�%3/�/߈9�C�ap#*�l*=E_כ�tj3V>w=�:�"%>�P��>!����ƙi��H�z�%�W�>��<̈́&���b��:��[u��Y��E5(�3��F�J��,�up=��.@<�XN~0p�z0�N�vLK�W�@)��{/��.4K��Ax�jq��]4�C,զ�餔�(�zĤL�2)�`�h�������(��N�t�+��)���y!�'��������dW�.S���f����?	Cm�}j6��/�J�W)�~01��#bߐ-���M-���h]МL�����ZREW�˯�]����W� ]��_r���C����U="}G8��
�:��b�!���N��������4~3�]&�Dt��S�
�|~�?�����PΊ�3�j��0y���YB��L8-�\_������`��L���i����M���rT��?l��$q?�w��EU =��rg}�L�F��uFP��F�k&g׿*�����}��s�[�F�sW�>�@a�5{��	`�Q�5�=��c@A����#��Vې��0y`@��@�wk�l�eE}+�W4��j(4�,l ������+�Ί�As@�i�R+��J&�n ����O�\��y�`&�k�Xs�⣨��A�n��s�W�,���F�e��թ���3aYZ���$�T�.��a�7m]<��F�Nr���l�����E=�k��Vu��M�`H#fr���)�	��+�My#�t�j�y}��wG��Ȋ�S����|���Sѻ���Ʉ�OӢs��򙊰�J5�����	���������ulﺰ��˽��q������w�Z�A�;=�w�
�ď��`�{�z�e�wi�W=.��-�9�lyD��40�e��h#Қ�1�� �t=��C�����/�"�A�̽���_dU	�$�MZ�KFR�2��{tl�V���v�!o��
����`�������4	�!ko���s�����|�=�s4�c�0Z�[��|@C2��tj�1�a#!Lw�!ۑ
cѣ����"V�Ϛ�Qu���!<�5(q��Ei5$?W
b����mذ�fk��텡������#_l���N��8�i����= ������h�=�<����u����� �Ej�,,�^t��]%��M�9���s�(���Gû�#sz=p���l˰b$��&�ߓВ�L�����~J����0��,���FR
<#�Y�B��$���/Io��~@���/����<Tߦ�l�)�05L���&� �÷����������.�?�����ER�NL��ƛB����_P�q0�:S��_�Ga�ěx�bJ�:�JBQ[_�r��t5[�((����ehnޑ�~��f�)G�>���(^��?ֿnEP�"p~�!2�Mx�g��"�^^r(˻6ɓ7�� ��I��3��Xr�KnaAX�/��3�����-�6,F���ʸ_G�R�>�\��r&ִYyFsf2��i0H���D>���i÷Q�W�b�!<Ni Q�~H�@���޳���4�,��K�q?�������W���
s>OA�X�ʎ�GKJy�����0۽.�ZR�G�17;��W�}��ۃ��k|���(s�лӴ�5�O��r�z>j�=u��O���d�2��y9`��ȇ�j��o�������ƙk�C�+{�H{�@ړ�4#)?������9�4-q �1��B,��!�+���Nm���q�s>�ǔ͗b�#��G`�&��߹4�_=YBgI	Y9)��p�B�V�����N�x�~������1~m�O�Z�z�WmJϏR�sY�N�'Ӑ�Ӻ騉 ��/=�u]�Zހ��!��$w�U�#mPؗ�ܖ���!f�=B멡;^U���љ�9F�d�\5g�XR>���(�E^��:����r�;�q��6��RO99��ѓf�;5`݃��W���d;��Vf<Q�j�wt��А��|�I�ԉAtt9c��p�f�3�{%��:�l�����8���ڑÇ��$&lv�X�7ʍg︫���d�ݭO��[���ROI!Y��%���z�dܭ�v�> ����/�B�,��p�b�E�,��v�4�+GI��َ{�w��L��&*��42�.V�
y�6f��L��4/�*Ȫ�"�璛��K�ȡ!V�f�|^��}á)�ZEV������pZff��1N������k��/5گE�I�nؼ�be@�0�<�,s~N���������n��>#oo9ܶ#�=�&���$p}O�}���e����ыH�b_'�?���Ja�lBʱ��<�{ �jk~�օ�'�,�<�5�u���Z��o1��~Sr�@Lџa�p�A����I �[e;F�6y3?�)dK�Qh����'��l�@��=p��:�����MIz�H��C�yb�>d$ �`{����E><���
ғ�Ռ�ďXĚݶ.�+M^ʙ�7t��g'�X{���3C��N+��7f������.�%}�.z-uS�`�Y�r�c��|�:r'���)E� XG��7 *���<��Tkׄʟ�!d=�zh'\�b�R狠���o+q�U��f�{��7:LO:�}A��|D$���<AN��ݕ��"��N���\��/�B�TW�m���O�iI�Ng�׫#GxȌ��2�O\a�4_W�R'���	��=�u����� Et�2��U"A˗�9�H?�Yl74ĈV�>C���hN�w<�ΜX����;�Q�	�2q���.���5�)T[1
2m�oX���3>Fڸ��'���� �h�����a��E�M�����?���f�ڍݗӣ�c�z#f���rNժ-�.��ө�����y���J9��x���z]���Hu�?Fe|1�u2�H_x�+!��4���'�,��V������ʱ�����D_(W��)0�-eoC��K�2�
{v�a�zw�Nb�D���R�%z��z*_ �m�]�T.�V;��/�h��{�!�1�x��ޮ��_}M]��9"��X�H���cVQ�����cJ�\;P%O�7c�x�
^E�hЛ��BMNDJ�Mq\�w��F.c��{a)���ꃋ�S���~q�ϙ�޸iJ�L�����	>������c>v�$��2��	�I�Q,�e����'��\g�b)L�Y��cz�H�����P[�<���Qsؖ`p(�N ��PT���&:7���*J1����p1n�����Ue���f���&@ry�ۛ�"̀�[z3�i��
%��͆?�r>+V�5���&6wD?�� ���� W  $�@��D��h���N�û_Q�ɢ����a[)�����ُ�-Z��"US�pR.�V�cz�,�����~�,�h�W8��o]ꧧ;KYY`#�}�
x���x��i�`1�3X�J�M���fVߧE)L})�Nْ��D�#5���b����o;RȒX�|"e<��A0$���x�*���:=Ê�YT��l�P-��ӊ�^��o�c�kq���j��7BH1�!��?+��C�8%0�������"�"i�m�A2�0��c7R皎�7�5��_W��æ,	����>�F��8v���-�{`�@txCq��Waa����$c$�O�w���C�T���<oFF�_q}?>C�d�3E F���cb�̫��1�\����	X���[	���f��|
%�<�0�nY�g	n��f��fR�p��DR���=�MȬ�[�rm?�%�Ԭ�R�	���'�;�(/�vF*�f�����*ՖC���c�o3�!��y�X�P���]�N��֮�l�j�d`���L�c�0�kJ�K4Y��fԇ|����G=}�M��4�l��#M}@���ꛑH��Z�)$c�} vvuV���(�Aآm�1���1�e���G9�SR��X��̥
�t�D!�k�Ƅ:c;���x�Np/Mn'��X4��<H����Ь��I˂j��LAP�����~��*fWg�8Zv������V��+�)u��s��}p_�E��1��w�����W;����G(�4U	�5R���7�ک��L3|�2g��p�f���56��Hbfj��uj� ]䔵��Cw�k�6'��F��zٞFJ���N�
����YZ�"�^�$� ��`4�I>�~�N�Y{@�VB����叵OB����.W�Я��*�,^W�������X�Xt��\�������׃s��.j�L�B�!O�"*��~S�����3F�!���^��g�H��-��.L!bC熿���76ٯƯ�q�������/@�xi�q�N����`8wZ��2j6�bh��u@R��������(4�UU��7�	Ɠ �1)s����NS�b+����ٰ��v�{N��|@|
��]�33��H:Y�B���A|-����lq��s��0��v��_C:���~$q�S��i��;��t����M�V���r���s�� ���e��o��G�x|!�b���.����:�P�)���4*��������qà�ODg>Y5��j+�����0&��M o_眞�(4�׏T��,�7Q&󷍢w�϶����og�l~�]��6��SAH�o�pB��fx��Ҩ�n%��1wں��h����X/D��V~Hp>�>�ӿLщa9�8`z���^ן��<&&\�r��F���O�p����jE���N���[J��C�0�����].&x��0��D���MD�5{����TQT��ߦA^yQS@��J�q�Fl����
F��KXG��1�H��@��,���K�P 4n�e����!�⺎6�Bw�O�y���,$�{���Z�;���>u�E�|��?MKTpB��d�wvtq���TG�H.�5��ɖvE�p�������� U�%�(Zo����KY�o���͸:�s����t�qlo��i�d�я�����d�u��t����O2�������p��+��o�(	��@��mNl龍ڗm1���ړ,��6�:k,b)۳�Q�{iNO"l�<YiM1w��1,����E����j�2��W�q&�<!A�ߝs���?�d��VtTs?�e��V�j�H��2�'&�������Ie�����lu	+r��s�E�� ��π&Ҥ�'hf[����0���H���Iw_-�	ZRWݳv=�����L&�a�]q�s(����3�D�a�=�<���n��"��;��<�<�˟x18�3 ��%w�Y,o��l�8�d�"�f�u(�4V�Dic�Gп��1b��1>4W�����D��ٮ��y��ۉ��!߇>� <{W�VM����J�ݟy�p��̚5de�����Ӎ�x�i0_��Rq�\���@V'v.>�Z@z�0�ߊ|�"њd@`v����kd�IJ꯳���AQ�93\X;��a���}�?���n���߮����j/1eaW"�b]Ơݝ��	���`)-�<���hKMƌ`̍5����L�]�u�u뚁]�� 7����o��^�������",mR	�Z`� ��i���š�� �����ř����'}����R+�B���;FhJ��J���7������MŢ�&�pDW=�!a0�^�*ꑅ�ӹ�9Jp�*Y���fY����������kz��~�]@c!_���_!�'�h��y�L�6�8�r\���[��Jn��9��=���g�[�򊈧�0kM��3���-q]��eȆ��p���#�pj��U޺qb��ɍ�ZN����^Q@����T�J�Qگ��u����������rĤ�)Ǧ��y]m�t�Xxp*������3�p��ӊ2�=��W���y���-�+?lIfb�|�����<#��4� 1�/�[��Ի�!9�sM �!V�D�K�Ȧb�ɻ\�����R0�8;��*�C��܊��0��i��o�C\9��B���pm��Sa���	'L��:����Q���+��"0�wjL����%`� ]�˞��}d Al��Gs/�V�b'h.�N�����e�~G�ݾ'��%!�H�{|��}s�-Lzq��h���i�0Dr@�h�U�1����~�BK��S��Ӕa�,��nĎ.��$o��#��c���)>��ݎ�$�G�������X�l�$�@l��P/J��ܯ�p�]�4r�,|�M87g��E��5�щ��M��Ќ�,}��{*ѳb2��sNL�6�����c�X��ܖ�	!��}^;��YyY&|���3Y߫G{��ɨ��	��߀g�����/;��߯���[Vo�_��cХ��aʃQ-�Y,�%�>;6F�?z��]z�F�ފ�;��"��%��	12�3N�<�K�zwN	�����w↮�b��o�(�6�y��^�tZ��Z;dr2��ikf�t�±t2h��,J~�&8U֓ �C��k�^)m#4�i/#͆l���W�X�6!c�_�&M��r�g�98�!���9�j������v�b֪��)��xw�^�T\j�\�=�wP-Pg���}�����wVp��D��U���y����
��K�H|��66.J�p��ն�gp�s�����}�5&F��@&���y/�mxZ����h�NfD_��!3���	�!�M��5�	u��Ɇ�#xJ���/_��>�������_�l��fWH������juW�z/m]�&��5�j�ɗ��h�4L=��|��bµ���1ܗ�B�ҤUV�$�Od΂�H���b�dFO��(�>*Z�9��@��i�C��v���k��Pd�"�����BG��:��f�Y�;*�c⡷���jz[�����_S��N�Y�_�i�ƭ܄I���7���w؍��(�$��pS�N����1�`��3���%d�ƪI�r�q�4��' 4�-��VPcǸf��Kg�P3�C�$���^kV�TM��g?l�LX/�h� �C�P�Ò��:��i����q��}K�9T'��7Ӓ+,հ������O��6뛗���U�k�!
LI�����7P{t��ҷ�ą����F.M(a��Ҥ"wo�)��a���?�Rt xnj���h}G
��3��ڿ 3��N�Q�C�w�0���_��=Z"@�*Yc�W#3�-��2m��'�Fګ�V�X�O��;z�d�M2�	0Ƀ��q�?ش[J��2�ۜ�W]&1�R@$�"�g(������D�8�ܹ�W��� �����0���Ȃ�~��
EeȤ�.�|��z�kie/Q�E��A�p�����{����'U�z$��m`6�:���#*3��V M3��EV�I~_R@싚z��7-�٨n?{L�,����鳬w�!�
p��6�Hd*�i�FHtާzA����-�*\�KCB_���P}�ѹ���ł*
J#�A=�	:�S��DXoX�K�����4��D�v%���IF�g ��V3w{Q0��la.%�*���s�򾂫y���������OHEF�#I���|�^k���	:��\Ih��N���s�RC_�Uۢ�r(�Q����nA[�c9��< ��n�aS��5����
xcC�X���rkT�Pc��\j��L
̵���C�K�F��>�����;����<�S7+Aa������9��N �\s��Z�2�5AG�)���:k��MWmEz��y�^�8���U�
��)t�.*C�R�h,�����ʖ�k��&�Ȫ�G��ׁ��ZqQЅ�i��f}�+vmj*���:뼏�#Z/�r�M���7+�T�O�¦rXB�U,,��^���!_��)���6^�}X$��x](���W�e>�F�F�=Vr	`҂\�K�?gj����|<��/��z˜[�܆�z(]��KN���>��kL�J�l�G!�7<;m�;�������*�r.ZR��=��u��2��CqC|A�GѫڭO�?b�n�5�H�d�K �k�����.����ئ4��	�+M��)[
{�<Mc7e��|���^�[+��cTH	� =>�m�HA.�?�N��8�Ji	�tG�S�7�6�q�l�gDy�Js�)�<�2�d5��[�yy�,Ù!�B�r�/`a�F�X�502���+U��,b��D���P@#�END"�����吙�Y2W@�ڽ��nk�l=9���w`��x�~�pQ�`���
���U�K�ܬ�<��u�cs�.'�a���2��8�r�8��l�EK$i+� �{�S��V$��O?/ݹ�P�T�w�$�F��t���e=��G�9!e��G�*��n+ �����s�<d�F�"�� �Y�szX��%�)�k��F���Q �J�ul�X��E5�����d20���}q$�������L�����K+����7J�����j���)`�4�4[tf�S�a�-	u-����� �0�.�W�]�5&Y��H�
�;ew��n3	�q����1{q�z0ͯ��u[��%�lɧQ�f���w;i�όs+ht0n&L��\<Ճ�2W�R�YȜ�*�������aAg������C����g
��E�%�{=�Mm��ؼ��.�FE�ˮ��-2$y�p�P��ti1�6����FM�4)A�Sv׮�냲"��X���D{,�J�k�Z�C�����'���-MK��x�n-",/}<�����ؤ��1��q64BVd��}����`o9�ê�+�W�����dO)�p�&t����H'���O��V��x�Q�؇K��.�m�l�Ɗ:��omeM�.@���g���<{AB����Q%�CAO<F�MM�4��,������� ;� k�����I���ȯ��p-�o�n*���}�J�-���h�L�Y��ZF�	!�ٓD�Xv8�bY�T卶Bu�/��~���*�N2s��6���4��鎭���n+����mᅜ��:qs�5��=r�n�[���Of�w���hۛE!�dM $�!�e+�!�Vg&�L��B���$a�s�-�J����P���kd'��=!ϛ0�I�%PH}آS�${Pw�ݍڥ uv�<��l��'bF^-�p�6��QL�AFjc�PrLT�D���鏽��+��8�]���-�o~��.�Þ)��t4EM;�;� r8ݿ?8���b�h5�'��e��<��+HԿO��aѓ_V���s��W���� ��<�~�i&�w1Wv~W�#��T�U%��,�y-d��o�7��Q�HC��ã���ıg*4C��,�Bղis���!ڷ?߯�3�F�{��:��/B���� ��DW@Q��"'�4\p��z�x?jൿM�P8u���
�ģT��L��x��R�^P����"\��]�|�p����s�Eï�M���Y�Kz�moxg�L(��V�W�h�~_�4��>��r
*��-ai
���=��0�����1|�qՄ31T����Um���BmrZo򞼪lB�=H��ر�a��NZBHµ���tp!�c;�?�8s���oT�(�2�	2ɝ���fLQ���O�Ⱦl��2���^��5q<٧���v�}���γR������8��h-�"ऴ�^PBis�c�\�@� �?R��E`�3�(����5��(t
��E�<�Q����Z����o� �r��|,�_r�Ƣz�H��+���ǀIU}AG���{��^�/�V��ݵ�m��k��G<��T��21J�~F��}�7�|q�~����+����5��#�.1�'{p�,��u���{�a3H%m�n"�)C���#�Kq(���3����%\46�$��/Z~a�d��zl���Tΰ��M���<%�gô�~�|�(��qҟ��ִC6��r�|��D����ed<YJV�9�kvbe�ۉ��.GԢ|���v�a8�������;u���T|{-
��,7�g��D�
��^"@;�c�)��s��e%X	�OQգ&_.�C��w'G1c��-j����Cib(�(�2#H*�A�*��T���!/�}b���NV�eH�z��I�i���|��M��d��
���Y�6{�P\|���J���9@xq1,J�+�l(�j�J���Ǭt���?��'1��&�<�f�����FT;j��&��0bw�/ۿF�4$=A#(�	KV�7�%�����#SI>�@���lC�;��qm����v
��z�g�ǔ+�X.��3�Q�-T}�ƒךoe���:���Mɰ@<���wP��k�R������#Wl����J	����a�S���~��|[�d�KFw��+��qa��i;��r�fP$`�06Pu��݊B[����5kH�-ђ�yB4��L ܄�ׇ)*	�"��ϩ	"�Rݼ�>'d4b5���"2HN����̩�:}�I����AsDBR�g���OK[��s|uz��r�JS��:��
OiQK��o+���"\֓A̚f5	�7E��S��d�ӄ����	 ����.���=�/�{��z3`�q� nP�V��_�J��h����Zb<�"��_��A�<� h�]�Gjp��8C���<D%��cPu��2�`q%�@CT��t����փ���E��!�p��X���̃��=�k9��p�m��>�����[[}�-�'�tPxj.�H�����˪
 &T�P�L#��Rt_��1s�m8��p�h�)uPR"Ӣ�e�`�_�y
#���߅1��2d�(�31D�;�����9;� ��""�}��YU=���U�Ej��cpS<��v_�{ma��M�m���0� ���<@�+��ZD`G�-�T�͡��-gJ����U�q�����\�^�.s���f�7N�nO&�A��1q�^���O�"�E��O���IHK�-=ʓۢG�ӈ��}N�;�;��v*_�sU��0%+�9-,�I0�����xC�֔����E�t�i��	�}���: �@�)��m����qa��0�)c�V)��\E6���!o�ϼ���Yn�$��w��-S������Z��T1��]�����;'D�����ǘ�u���#_mVS4���h���Tp~T8ʟ>�1�uzzݥ\�&+��E��#I~�(�ǲ#��o�-�^؍=Yse�ȟm����J�#��s8�US`�{�Q("��J)���^�M��3�Zo��!c���t�<�~���(*�31H6l���M��kE��R�#��U8%�P�Ȝ*%R���a)،�!�^�l~͊�;s��3q�{�X��lԖ�ӅJ��a�b'jK��g·V�H7���X��N!���}4�[�m��ޛ��T�O)��2e�Ԁ����/��86[;�6�Cɏ�n��(���SMr,���,��?ճ��T��GM0�ĉ��G����wj/hfw.�?1��^
ö��S%�陳k�������@71tԯY�Z[���Dv�.�fy�	��&�;�,�S#�0�<���� k�E W���c��F�gR�?:Kp�ۅN�p�_H�����)d��\%��]x��L߁�1[Bp($�y�
�O@�f�[=�����ѠN30�,B'��]�$�<D��2�>-�bȎ�W���[���øT�����_?/��L�e!��0 �հ$�@,l����L6�&�C5�Ѓ��[{f�75^�$N-������up�a��1�U�%t�������z���}RAR�s`��_^&� ��h1����N��|�Ҵ͚���ĽWx��I��w�'A[�>�M)��e���ߗP��mrR�����0��kWh��I@�k�1�w���9!B\)61/�M1��}WѸ��@����mO&���уX�J�.���I.O���(�WK^�>�^Q
�G�q��;͉Ӿw�ȼ�Ҽ��|h<X;�W�8&���5�X���N��E�d!�G�A���Z)X�N3����SH�q�`������Q��W_$߸{[ �ǯ�;��0��^��k.0�㛩�Z]�aP�c�ֹ�QTܘl�3*{$wo��^On�^�a6�DzuQ�
���>�[�e2���\��X��{�T�4؉�۟4��#M{��`Wչ	����*��n�P����
j_��yǤ��X5��K	���M���o-�V���u�3O;��F҃Ϗ�fu�����VO��^C�"�l��.si.e6�f���4O\; ���2�d����f�&;��4�cR���у��P�<(�2�� �GjA���d�Ŝ�c����纨��]ߑy ���I��Ym]I2R�O�9������U�[�@$F2e�����U��@2��@�����fj���M��V9�V��Q�Os�X��ͮ	�)��p/�x{+`M#vO.�`�U4vv5��:�)�����%�z�S�G��9OWa���#D�p�[��m�kf�)���_L���[X_S^��NL	�8kI��;r��[N�>Y�j��{=E��o�S�j��P}�\`z*��L���P�,Z��K�є��<���&Oc��
[^;����}�1"#,	#�#te������}��q|L��"{���O6\Aqs��>m�82�a7�P)#u1��<Z��C��e��/1���Yi9��L����w��]O}���5�M������DwGWC0ל��X���-Hv��c�\?+݉����Ո��C���*�`��49���Ӡ�nBb�.Kv�ħD���\U����j�M�YS�� �sm�p+kq�Fr�6��H�"~{�a�����0C�+�R~��!f�\�5�%�%�%]W�P�[�p���������J�Kw��8�Lb�c6��:�p�����	�����UZ?�V~a_�V�T�P;6m`����Ҽ0�~�ܠ��\�M�b��@�����{.�⭬i.����ۺ$7׳�!Xɀ�����(���y�<jE��D�}x=~�LO�ɛ��]��T���$���=����J5����F;{W�yZ%E����м.�{�H�E(/��G�]��99�%�Y�Zh?!|����|��:�%7���o}��C@��<��RFI��C�t�rB�_��n�6��Yc�(n��QRƟ6l�[�m�/@=��/o�վ5bz	^�U)�� ���]���\,���<�GWt�D������XkrުZ�f�`lNW�W�i#�u��iH��.Dv0�ĄŎ<m�r&�ׇF�Zc@jى�����ő��)�g�&"  GV�@��W�)C@&a�$>��c^�|�;k�F#>k���זֻ��^""R5�+�`+��<����鸩;��-��@��;R�o��tw�1��na^���EN���@�A��LA`�*�k �CJ����u�kD�8�)-�������q/G�l��%\9b\ך?�����e�r����z���K'T��C�����-�P�:���

�+���a���^LlAj^��s/l\'�]���EUd�8/ү�=� ��F@ث۟�-���W�V������Q�EE��#�#y��̍ �-?�(����~O�F�2�;�{�8��p�XJX�Q C4��T�6��kG>^x�aӬ���IT��Vg�F��H]���#~� ��,��4$ (j����4��J�g��� љ�7����ݗ1�CB������V�V��M���������ʬ�T.�:�ND�^�?������^&�ɺX;eԪ%���q�p����^.E��S���gqz���ah+kv�m}]L���Ӆ"M���x�A\�cކ8���f��(N�K���DD0h�T~�16Z�f���)/��9FO�k�Q��ls���ʎ��B/6�]��XP�Ȱq���P���k�b|;��I<m��;�/��i���:��� L]T�9�'����F�~�7�5P��j�6TIv~
خ�T+��!����30/��sq�
�t����Ƅ3F:>���u���������J'��w+�>H_4�i���Ѷ)���d�!P&�Wn���w~��w�(��ڦ�ԷP�`����'sk�mܠ� �8��&��9��&� �(3�.8�lM{C�oB�_����<qpL���Mq'I^pFFѓ?����C�t�Z@<�n��h�N;�c����Q���6�p��4z��Δ����W���4�a�	E�j �yQW�f~?���0��At�>��p>#��0[( :�6�Ԁ��ԃ7��<Ec���Zt�Q�4�Ĝ������ai�B���!���s�Ɵ��ǹI�|�Vf�@�g�۵T.�~ŗ>���׼�����o����o�@g��q���R"ɿgQ��|��3�e�%OO�.["���]@E5�G1���#T}�*��{�lZ�8md�!48+h�@�t�Ю����Kd!r���jA����R$!��=��A���q���ʮ�uj<Y>����h�΅p�4�o@�W�Ov3�� C��A�{f��k�ֲ�M� �e3]��9�����.z(Q{׸h\����ѓ��,%B��}�$�|:O�F����_�!#Q�~�&-;z`��Pj��� 1e�'8��-Ɍ1�:�����n}m�Y�r��` ��.g�^��f-3�wf��$�0t��~���,"���Kg���9S���/�϶{�}��|����p/L:�jV~���U~F5���r����TcМ��H56 ���1�s�3vVT�>�ǽ=�������Y����z0�[b\�O-o�;�9��*�����Rc�Y�љ�r��R�-�NW	�P�I?k"���)z+<���-(,�2 L�b������{�qn�k��<�򆍪ݩ^���
ꪜAB`PL�"C6�6g��Lg�����l�U��8YvSd0i�S]�Ei��f��/��v[�h��)��9�?_���d�����x��(���Ln�ҽ�m?HH�n�^��|�Y��T�e8�V�>[5����Gh��+�`8˥q�[ң�@�y70���6ax�{ ��7U����Rj)+�j�j}ݐu�3��<w�x,:��?��}K�j�'���D^�x�N�!NJ��Qr���6�g�BiN#]�h���؇���Ji��֙幞�AD2J�_M�;�O��_O���6!���/[����^=	c���pi�)U-X���-]���_��(ϱc��j�lb[�������o�_fXU��`�\���'�C �7��s�32{�%�l����J0Z{zQ�-��q1bƎ��=�M�%�'�ې]5T:���
�G�"�
�&�+�/�1?a��[
���C�U({3B㤀Q:�@{P�7g˗\&��6q�Y�o�'\�������d�th�Z�o�O�-~}	#�lʲ���u7�){ZΧ�wwΌ1�伺6a
��Nk�j��u��k�������-���ыe�ں|GC?d�±���t���v��t��v�-N}��T\�Xm�{�`�q��p�k:p��� .�*�I�T<��z�q���JS"����$���p���o�4�N���P���s�x+�����bN�S7&�����R G���r����p��JR�)�:'�3��fy[�Tz�z9�
�ޫu�y�	�(�}��,��RI�&���]�=�
�߲���L*������N�8R��6��V��,s<�>�1Ddg������,�DO���~���s�����+�C�Vp�?�]m��\�~����`��L�X�� .��{�1�d0��5��F����I��n�b.5�l��L���6t;�+Ѕ��=�'���A�]D�W/�؎��C�}w���U���ͫr[�P�Q�WE话-����<�Z�a�S�9���TN=96A�7g�ᨀ`��"C)�V_����2[��ҭ���g���FjS�įGE�P�b�h���ư��8��Y��9��Ǯ�:EF/�yR̟�A�c���p7]
�u�+铐j�eǣ|��!��J�