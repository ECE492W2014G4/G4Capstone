��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|̪��q[�d����0��>�����@�Q�b\~�-�X3i��ī�D�M����|��Qyc�
4�HJ+⿕����=x=�;��_N��;�Z�g��0�1�Wl}���a�K1ǘP6�R�&a1qgVZUJ���ON�Rv�շ���z��}9���W��dњ��:�B\���_2u���ɧ�J��8M�{/aߒ)x��1�"�qC�6칹L��tG� ��0�٤Nu�Q��$77���~�vA�&�q�[ghܥ�γ��vV���j!gZԤ�����w�#u���OF���6�i9�.�������#������&����P�}y�&�H�3y���Vm����_~».8G2Վ�6��2��'����Y��O��g�t|Q-���9���.��c�bgn�94p��%q0{>4�V{%b�>rKɄ��M-�Ǉ�gz���j)�c���YE�U�#�.�����)���;|ɚeܘym�3�}�E�G��0H���ڎy���`�]i�A�vj�(P^wx�,���ٴ��H%���r<�l0E�����"��p��[i���s/x|�s/�������:D�7�d�m�7Q#��q�v_񌙭l��	�6�YgR�"�MX����=��L���¸���wI� 'k��ۆ�w�cZ����^8]螗TЎ��߀���ۗ��(6�v�9�7��FQ��`(�L�C�貄[��cܩ��ۿЮ����(��0x�����zU%?�����!:?/+#я2	��	 `&
��A/��=>uýH�I����:�[��d+�GM�<��^�*���-�6M�N���Ra.�.�v\�)?%�%��Y����d�AQ�����Կy��Viy�u� },��>����UJ�O5�a�k��J�0��+�W�?�޲o���Cp�����6A�D��e�L�2?S��mR_'V�����d�8�Yf�q�:�F��;�ơ�ở�ؘR$2����i�[�q�`��� |,EJUB)�M��u�{�WlMM ���鎃��R���<�@�M�:�῝9�\+u�Tw #zw�<�O���'�(�iX�U�# ��uwC���O��_ZM�]�~J�>�Nz1�#��K���(�&�V����,�@��ߑp�er�gUr����ȩh���d@��m�C�5�]�%,���e���!sU�bd׾He#x�Q���05QY�pW}�2�����i4ݰ�K�"��Ǔ�ݗ)�,OW�� E�ra���3ڵ��4Z����j�q��LE�ٴmTC�.�5���p	�b��*ר��$dV�&*��+�y!ߒ[��e7���k��E"�}^
Z�7��;�ӫZQ����j��J��@P�׍��b ��D4���O�j/�\�M��Ï��F&���{94�� O�.�74K��m���z/~�bۄ�v��׳Mi�<����.QK�z�}xe����!%�zvH����;�3g�'�t%�� �6�*C4C�a>�7�w@S�ے��-��g�����M1G���`g���_<��,�+^E�>���8Xu58 ������q���.J������������5����_�<�fp�?��ۀ,�8&2� N��M�`�/��n#�ߊ�}��[|#�bJ�� �bq��)܉�8N�@���	�)���� �:���P�}�|p�ة���`09�*m���x���/�\��
��v�ғ?n@x�;
MZNH{�l��B�ث	�������l�|�4���;����ռ�Aˤ!�iw���W
�	���
B�Re�h%V�]���m,�8��$�_�CX+V�쪞g�|�*������-�5���1R�J���2�3���P�C����@�]:;zN(���籇D�x�q��x��?��?�Q�G�ƨ�n�}l5#�8�]ǯ��\�F�n��`��i���c����0xz��I!��p�v��5)_�<��fwêb�.�Cu&]LAf?��j)�L�U���.;���
�_Áلm�-�V�Ә�z�L��NKTRqT�A���A�;�
����p:[:�,3��s?D���wq�L^=�$���
�g��<����W���P�<��s��JS�/�X�YF�/��Ø�d�- ��'#Չ��p�yr�@���\�8�=pk)'�]˝O;��V���q���ϖRHe�f��E�� 9���8)��qm�ޒ0�<���a���,T=��RH1����s5���s!�Hd�x O��|�����`�骺uwMx�m1��
5ڞ�2i�'/Q9�F�o^��2�iHD� (��#�w/H���JG�?�{cCh	�%a��fe�Ly���P���8UC+���1݌8�$�=�3�(��`�\�������4��vr����iߵ��z�e�0�_i�>��#|�ˋ����:�+�z@i�\�e��q����lU���:�0��Sd��؆<�_�[7랝�z�L���� ���X1����t&>/6-e�A��5��^oӳA����+�H9B�Alב~���_�eĒ5p����p�4[�WÂ��T*�Fu0�6���F���6�e���-!x9��QD��fn�!D+4K��ɂ�bӸTA�"���Ef���Y@�-��p; '�r�h	��
2 �> V������C�3��@s9%E9qA�����O�I--��.��o`ō�*�����:ZP�����|�:���B��=����xdGѮ�åf}��y����71UuAW
К�w2�������.�?Ut f탩�A���n�m�_�xמb�%�2��>��E�g�Nz4ֈ�r~$�*�k>���v���f��Ųc�/�+-�SkS�U&r		���KG��7�ctt\�a��ܮ=���BO�
�~���Zv��BE|u�cИh��4³�n�P޲���S߬:�q���[�f�N2I��V��{R�����|�N�Y�h��⺏�B�Yr-����	�2����&a4g^[3���`��qǐ���6W��r���UH�;��_���#�Ѩe= �,�Xt�&q�gs�˲<X��\>~�h�����{4�᭒_�ʕ����p'��
<-p��d��������i���m���xpY!����4m
��--4v�DU)��,�m7l��T�3G0���>D+�Brh��D�p�H�y
�s���Q/]Q���K�$�d����'V1Ϡ��S�p�/��<[����{$TU��">>���	���q��;g5�׏�j37G
(�� +�,� ��m��U���X�s먋�i�'Iи�+�Z|-d��#"1v׬����L=��� U>g�XЏ2���*vP<ZB٠%k}���ȟ8c��;�����Hu�҅�U�uf��n7 (�L�̉�J
!\s�3��R��m�'xQ���ό<�������t˒$���i����Pw�&#�%ee�����~s��ݨ6�?�ε���s3S�g�F�Z���(c��V�36؊��{|9u�l\���Җ��F�<D�@�>`V��g��K���d�rn���>������8.�7D%D�{�*����S�'�0'3���6��;��{����e8�Ej����]-��r���0D����3?��Y���B�	�p/���"�aP��P�BK���}u饩�Ǻ�����Gr�\0��:�~�i�bl+��/_X��P�&�BO|/MY��Po��@��ñ���x�S��,��������Q��J7�H���D#K?;C��ޭԹZ�����)�-2��!��I��`_��*�-x�àh?���'��Z]�Xew[��_��I|���o�Ԇ���� ���5A�	��G`�L�(�r�na��	p�Y�+٬P�SWHcn|��Hmp���8�a-�:��;؇�S0�숀s=��j�zp���,rԔ9�3a�1aG�\e�4J3��j/ܯM`��0p��t_�n�(��(���pF��H��h����@�m���1�·�b��-�Xo?�ʱ��(
�Pݯ�h����0���S�Q7%��l�Jf����a����96V�WQ�E���E6�#d��xF}�B�Y��z��o�,�x�V�:��=��8J���<e�ճ&w�Á��37�)�ŭ�^滑g5�e��gUGZ3�����r�:c��FNp��x,�G^��7��Cg���xF ���P�_\��վ�Ԙ� 6�^RIO�Ù�-�뜓�&}��P$O��� 4#�f�ӑ���AL�Lƣsf��6�P�״i&~����$������R�a�?"P�����F1����]k�A7�*���7�i_��f��H�>��)�y���C���3�ZlW ո	"��{@v�:�U�Z��q����, �>Y���j��p���a�9E�=�͝!HۂJ^f!C�����Z�*q���4*q�r���p$Uݘ1Xʤ�*q%y-��>���r!H�e`R�a�w�>����P��kSv���'v���L����AJ��1-s �W#h ϿG	:��yHkԫQ��l1=�_�՗�����]s��d���t���v�n�r�6ԇ�6��D@�=U|�YN)���ω�9�x�C�O�S��w��)�V��d�����Nā��W3P���JE�*'��fv̬�#1��k����u�Q�{��$N$J�*���
��Y$T��0p�!.�rݴ<����x'�J	n`��(.��L�I\'f ���!�/���a�:���<@��7��=��z�|F��(~�i��'���?e�����&�0�i��N�tx*r^{���F\���w�q ��s1�T��N\E��n:�<����8]���;���K_�]�&��:�&���]�Qc6��KG،k��#OkDb*j���"�ٽ*�*�}�T�{:�c)�6ʪ8���pIJV���A)O�=6�c�;�����-	��R��|��������Qc`#.ۛ�<F�6�"�g�)%����%�>�W��Q�OR?��F��YK��a�*�c3b�n��NQ��oW�x*�Y(Dċ�mdcR�,}O����A�����@�)��j�qr/�1g�4���5�b�\��3�Z����C�(G$7�"�_���H�����㄂�*��o���ԋ�t��?�&�t٭'��"��9Ӭ��
d�PT����QH��O�O��v��,U !���O��>�@� ��d���x`�h2��~@�EI�