��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|n�\&�����[hc�>Z3�S4���"KP�$��h�I���@�O��m�SP��Y`Sڲ�G�����'}�f�n��Jf{�k/I_8�~5b�(����q�OyC]���w&���{���t�Tג��wr��[٠_Z�m�Q�p*K��A�A��� Y��������(h�!��~���H9J�u�\)_Hw����V�d��+?�Rm{A�9=u��7b�]j�0{K�ɷ��c�|12��
�1LT\lZ�F)�N¸_)���LBs��]$3����5q?�",�oeM)P�"�gO���Do�Y�{k��;|M��F|�����'̆��<��Y�3e��)� 2�F
_;?fLp'���[[ɖ̣�����������T�J��QOӿ��kj��_�	������ �h��_q�t�[woa�$��x����-ў�$�>���l4�"��Da�q�ݠ���`IT�yG�b9��[u�i@���R���l�h���Oۛ��G^e3�L�:��ѕ��Ao:�,�g������[�{�o�*ܩ{��K����r�_ �P�\@�G�<X�Z�����fn;��C��T*9��scK�ÁJ)Ur���c���x�H��6(��V�=�ڞE�&l8z��QTr��	�g0�k���D�׏�Xc��zzģWR뿨��
�K�ȿ�̝�T,�B��r_$�C,�F�4rN7���H�\uR�c��
Zm�Y~�.��Ţ����K���ɱs���O���z+��	^@��L��:}!GM�x*PW	� W�/�c����
�4�~������B�NƁY~O/6N���X��,�$r\Pp��z���<z��!l�QGj�K���k�E�/�5��/��Tӧ�R�{�O R��
N�C�yk��k���Cg�Y�KM�35�h_ӳ%�H���Ԫ���0w8�&iV�?�n���`��I1����#��j�'$��d^O7���(���m&�W�<�|�E������Sx��c�广#��ӷNL�ld��ʩ��B 	%��&�ws��橺V�^��vc��m���o��1����"�nEN��T�K@�7�F8�%�r^�NT�_�GWD?�,H�O>�b�k�U�C뤙N�
���u��;��GW9�	3�T�(���tQ�R�/ ��&�����J��	�G�U���g:ka�"6Q�+�g�V���1O��19m��}�����Ǩ"�{1x��G�'�}�����z��&����`}Yǃ�.��L���{�Ϛ>{3qP\G��ʗ�ۋ�S�����Ѕ�xP�6���/�TK�gK�y}wDi5�"_1g��c�V��Y�I�� \���&�F;��-���7y��������B�A�;B��Њi^[F�C��:�cpç�����#����՝`U3��VY���d�l�Ӌ��'m��B̍4�����C���`�����-o�+�ja�_l���"���o7�-�7Rp���L�l]9� ��M<���K�7������)o!y��z�_�Yy���!�4L�I�Z�˽N�$����N�%˞σ�ϓ9AW��_K(�w��؛�=�O?�;�q��i ���Mi�z �m24�!C�Re���X�e_,��F����<I��2�.Y��t�3M^ݷCO����&�_�*ja����Ǭ"j�N@��*��g��۵�����#�TZ�.��W}QI� _ڋ0�$��tq������tq#/���%�:�.��P�XJ<C]'�#+;��nww�D�ޥޝ��_x?s����B�T��Yҥ�/}X�cgCw0=U�������4â ��*�$w�߮�K�����Q�Q4?��ǡ�d �Ƨ^�.����ȇK��k�&?�Ο��\CS�!�VNp�w]l���
�-� �Yd�逾E���^���4�"�"��h���ʪ ��Ut�M����`�L�d���,_<h���{�ݐ�6�õ�6�i诙�dw�R�q�'s?�)���_�5���Q�˻���`��&g9�Ĕ�gj�t�d>���{A~������S�'"杦�����y�K�2�ʻu ��֠��˲�?�1j)n�Ӝ㖦ժ�>˄���x�l��v��.�l.��^�����G�|�G��w~���i�Г���VA�UZ9JˏU��7I���KI2�H5�Ly�ae�X�FB�[-�0$F�G˒��g6�7t��5��s)0sj{_�N����xH��^��?�P�@�%��)�4S�����A��TXL��[�`
���Q �z�$�O;
��:�����w��|JU��a��+1��\g�i������V�F|!�\L���.�¸���v�e���*G�H�<;S���p7&^��x�;o�ђY-<���Ե�[���eR�J�R���T�G�ضT�)���6}��l�4e��f����d\~K�-|
<��'���%	v��*���8��>d���u�{����|p`�ϣ4 ���0 �I��F�P�'Т��mDSX8	��p�C��%=WH<ڼ������?�����h��r��gK���>|.�C�j�Npwr����$�6�`-'X߱�AY+�e7N[�0r���p0H�F�U�@�/���'� ^\��|B֡�m6	�t[�]�=�5?:!��j���(��� �c��)�-;2��3�۩X:�l��c��Tj(�����D �s6��t�X�6������ZÁ�|׃�;����s�4�������2�(�K�vD2�S�-j�F����`ĩ��3��b���ˡ���Weq��/�(��&x];�a��ۭ%��f��'_�ZǱ��wİ0���y��_Eu�{���!��uV�aK����u�֋������L,H�u�]A�����iTF�1{�E��KJk�N�j�cڵ��M B��4=�<�#�Q.�ޱbj/n�_M�{���"�K�Ø���L�&^eN���n�l5��y��e"
�F����`vxā�X������I�E%4m�C#��t�?�0��J�o�� ��aB/O9 1��D�ĝ�ؓ�a�P���hй��/U��	)��>;�FSKgj$�ua\w:$��w��!ZY��ĳ�X�I�Mk��8������-|�gD<�P֍Ҝ�C�h�)A�hQ�2߾}�)�f\Y���Ҭ�y�L6A �t�`�B�)��j9���=1|��y@w�n�v{�f�����}g1�6�mx䓈bϱ
C;FvuTS�M�c:PH��/	��`t`��M'�����B�4�o����}�(U��y�/[�cr|?l�5ʿ̏����n��Lw�}ٵE`����G.�̧S�E��+c|6/*n�_+�S��K�=J�:C���[��zy��v�V�{��UP}>z%Ԁ�,��9��+zc�p�=r�6�	PcO��棃�&�̋��@�+����b1��
d�dq��e���1�B�>�EwcCo��:F�\��`���~������~L���fu/;����?�
�,dހK8��	X�@P)�"�Uw:����oj�b�ʨ�Ga�w �I� X��\�\�h�Ln�	78�|��9c����v2,z�~0Bl���%�k���r�pkl��������f%1��$���c��]����#.��Ξ�z"����D�?甀X<@��J�	����>����<g����;���-KyVΙ�iH�kg�T�]������:�^�tsS9$-�^n�#0�M!����Ӎ�Uk�Q�H��$�)P^�T%�XM�>�*���/b��pjo�PׁؑC�\�:q �:*�a� 9�cP4�`�V��2w��
��S��.�.������\I[��1��� r<����j�� 5l�V)�;�ϐ�-/h�%�;ڣ���K �iӀ�ˇ��揵)����dk��F��7�����7&�y{��V���dڀ�&�[���A�M{6� �(�T<�'���l�<�-�I�]�b��<�X�ߘnU�u���U�������X�~M6�%v?��ޝ�{��劋ԕ�8B�����ܬ��R�'���0}����>Jpb�8M
A��q.d_�z
�D���$5PH��*ͬAs*~FHbW;��*Ir�2�pK���L���p�Ѽ�;��iP��W�w��f��LU�$v��VJ⋔�G&�a���|u8\�K
hBY'�0xjt��ڡP0�$ �"�
� �$�ˤ� 7O��0,�ȣѕ���E� ��~�%c���.,���E���+g��O�b�\�n�ϙTO�zwC��#���aE��)-݅ƌ�������H?�_�/��@MK�Ka�A�/QVء�F?��꼏4x�cY&��"�{��y@
��nbA�nF����U�:�(+p��m�|�r�K���Ř�Wc���f��m|6�����p�r�$C�c�4�5���L֎4��,�f�$�\��P�b��<��b}�Ũ��q���B��9�+�n!�迤hYU��J$f�B	�<�	�����뾾����"�{#? XR_,O�% 6n(�<�����&�3sp�R��W"�x/V�b�v�)�����G�HI�T��th���[9�������h��S{ջ���'�R@Jוߟl�5���䟷)��crK)i�)J�HE�̳C8��-��
����+�Ӗ�����|���E�9y��b���T�6%�=���9'��OhFr������B踕?�:���ݐd�1�?�1�Y͍���nR(\i���ZG���]��:I�J^�s�e��I�{C���� ����E��2��u}]|�^��We!5����ˮ�D �Q�h���a�"a���V>n4U;T�15Hrn!R���G2�O(@ߕ�9�2���.�� ��$�Xk/Z��� &���Ldj�J�k�Z8��R���1"OW�(��U��ؒ��?6L�.�o���籦q;��'qw�V������gF����
,� ش�0%���+|0�M�&�Mvrp���!5���n#��b�p^���_���s>ֹp��[�b/�hذ�Ic��B��-�=���ۛ�e�(+j��;�>V�p����3��y{ �=��ء-zqWH��.�����!H��A����b��qVyJl�۩�l�F)̋�.1��q��SZm��֧ߘ�e�������������� �RT3�
�Qi2dav���Db�� yQ�~�'�fJ�s�-������R�
�=-by+O'��\3��qlr�M{�;�ɴ����:}�����Y�6Y��M���˕��B{���������H�H��t,�,as��1]9 �C�h�!���~;��ze����%#I|��o-�hAL�>o�=�G�y%�ͮ_:�-T��]:t�B�4�O-��(N�ɤ@D�<����=�q�܎�\L]t,���7I{��w��4�i�����Ϳj7^����p�X�e�E�j2�Y��hQl���ÿ����O��҈��xH�H����w�ŷ��gxX5�u�j�x��j.`��]� ��;nv�%VR���� �<���p	Ztgv� ��l�F9!�0���#I;��|���_�*��=�v����-�o�XstR*���-0�{ ��B�O� �Prk�u |3�,���7g�c"yׂ,
�>�]�lz�FQQN�.�ـ��a/��-�
c0�hɶa�fE�R����F�D�
��&-����Aax�?�O�rV	��� 18c	�o�a� ��y�8����?�F[��-}��R"�i@�i$�R��n�E��Nlq�e)(��!9Sۨ�\*�)G�@@��Fq����B_�Ql��2��������Ċ�c�Vo�MjQ��ǅ�7huEG�[��j�j�^�"��I͡U��}fSU,u
E0U���?%$8�����}k&@d7���{d浪2!�:v.b��W9z�\��ӹ||MQ�$��7q�0�l��B��l��> ��i�>9$ q�	�k/gO������	�UAm�V_����R�Q������<��I�B��U֓�?\��w\v�QLt���u�� �%��IJX�F������NA����Xb�
� pIƏݦ�/��%�Ǯ�*�]�O�[HU}����6�^��H��O�]��*���B� �H�b֦�Cٛz��mH���P�7do���:c6�	��h ��ֽٙ��3��)]?���N�O���(��W�j�����;���n�;f"�/����
Uv4�:��wE�l�s�S�����%��w�6t�F,2l�>W�]�.�]�:���zvS����6��+HoL��>�%_��ΗŸ�lxl����,�Z�6`%�0i���QĦK�N 9�����/vr�ԏg&>����$�5W�D���
�774E`�$N�$c�q�HI�?��԰��i1�f3� |��R'�[R�[�����}>�3��� M[���r� ��m��wK*���$r)&V�����}����A��p
�8�ФD6��OY�L��h�W����M�ߩG�����vv��{�CK:�*��i)Kˠ�<>L{���׳a(�t���s2$Նbs��evn=vkh��r� �S
�`56�������g8z}���N_��6���Ⱥ�I�ǯ%i¥�@���hL%�&�wM
)�+����@��SB��>ߒ*Z�z2v���:s`�TiW�0Ƴ�e�AM�_"҈(ϓ>_��w�G�8
F���%��sч,�ûܟ�Y��"�i���=��s�K@�9���l��f4I}~K ����Gtw�o��q�/� �7��X8�&�}LU:�%HIӬ��h7���Z�H�0O��#Q�R�r��>y�}�H���S��� `ce��T�7����U�b�$� B����ڷ8#gwi}xEz�6��5J8�w��G}��~ݦN��?@*��yљ-�ѹYt�O�����(�aN7�!$C�,�k�+�_�01#�B�Q�i[-u�Ʋ熮�X�(ؙV�D����)�����I��K�;+�]ʯ���1���h�#Jo2�?=��O+p7��/�d��Q����ڻ��F��l�[�:�܍"��>�5�ge	u�3��;��cAC�{F@����j��?��2s���q���{
��؏�V2&-���Z��dg �yж���bH_��	�mD�_�l���Hj�����Q\��>��I\�FE�fkaז�yNํ��r:��'w\�=p0م����jT��L孝�S��g�څHB7�C{��Y f�� yk���8����ߎNw�����lmb�
�����Czq����(�]�LD+��ߵpU�|�(H2��ŹU?1�����5؍��b�E��{(���Ձ8٪g��B�j���A4�x~��m�$\�~Q�N�Z"k��)-��:P���S��K�6��Jr4�	%�k����n鯱������E�v��&fm�ܺ���]q��I�.G>!ae�^�F�s(۔����������
:�������)�����.c�G��J>��]C��6�w�I���h�A��^�j���U�mU����Tn�\���ܺ	�f�ݩ{mu�ϸˬgd��CٹJ"@qF�C��;��

�K�2�X�f��,�52ݗnڑ�|����n��F��}od^S�+�ݳݨ� ��=�F�X��>�N X�1޶9�Q�;��Gf�i3)jP���Q���RPN{S����h�\S�呇�SEw��HR��n�(Y�Ќ��t�����ʊf�z?6������v����chvX�v����Dñ���$���op����[�/�߲�H���q��9�sx��p���?�ġ����i�A\���8uL�m�|2�7�#�C��_Va���\R*�cEd8d.��q~㱥U����&�~~��LW,�6�ߦ�Mq#��6�x��Jup������J~%^GLp��"ώ���|���̡��nҢ$;4��B���6�3<�$��f�Nw�@p���~e���~tO���h-� @Z�#�>ۅP�B+�GOvbR&=�Kt�+����<!>�loJJH�1��|&��TŨR�E���~��*�|<s "�@ޑ�٠)4H���j<���NwI�#G�j�?�g��'���jL�,��`�sQ6��s����(�
�N��پF�--��`V'{����Dp�͟]i	i铑�GWLa�/��⼌����������[��L�H*:�?��� P2du�=?�&k��w�P�{|+[�$�.������|!���;�m|����I����v�<�`�������SKh��	�k���-�!S��9�L��Ɥ4�t�b��B\G�a��J�f�m&C�GG���@��t��]d[-H���y5��)'#j�SSk��Hi�41��v��]�V�^�6Ē���̍Ǯ�V_Ia�ΨF�?g��fiz�cc ��
�sxFF��ݽja��M]����/N9�m���4:���P���Pq,o��`�C{Uti�t��-��k�	������@��Pr�ܟP]�Z�Y�,a�&�A�U�b�ʊs�Fu���pݝ��^��[%=�fV��%t����X�a  �.����^Z�Q�Կ�ö1h��`���뛝����$ybO�m"�D��Vvd)������Vg�����	�p��H�E��ѭ�T0Qs��	v>���:qy"f�}OcQ�t;�,܅Mo���	F�����G�K�g���z��O����FXs��/3H��r\$��)U��1(�W`���a��c �ؑ�s�gǸ��=C��z�:rS��C-��1R�,-?IJ�R���c���#cC�"��Na��tb��nKs���X�K�Xi�'�h�d���BÄ�NB<r�����#�U��<��x���a+�~�q$9
���#�>=Z$Y?��兖�bd��5̨�ԣzj:{�!��k~D@DH�����\�U�K��H��@aȘ��#����R0T�Q�/�/��(�cTR$���i �����D'm������3Q�.�ʛ���$?�?��x.��D�}�?q	MA. ��`��S�.	���q���ڐ�̜�_T`Y�XJ햬|�xW1�7P����کC1hP~�� p�v�W�`w���FD�/��S?F��?e�ǭ��kר;V
8��K���`�c?MMSؚ�:|���Y@���"�ׇ�k�T�����~t0̏�*�TX�X��e&=��m"�B������Ù�x^��q�A� ������.g�Q�7 �����}Q䌐	�v6�Rl[��w�:���"P�6�����2G�pj���l�w�2I��$��5�5��gYP/�J�l���\��M|<bN�����K�"0��˒0zc�S��N'V.R�*�R��v��g]�ECw�%{�Ρ$=i#>��,����bܤ�����v@�cD��g��R�sl�۽eX%
)c�U�
��N]���ٛ3m4��%} �1�-��7��I���Eo����v)iG���p
3��lc5�Ha;�=At��b����/�A-�J�Qe��4 �,���6��4C�3�� �����B��w"��a@_�����Gm�ЏvʁLA�VW8��Tʅo摖���r�Ӛs�
�
��2�~�十{�-��븣@4�9N�f@_}�%�E�d��%v���ހ;ޅ�y��bJ �k{ɫk>�Z4��e��ݙavb��iO�z�&��*���w3����"ؐ��&DE��!Ɂ�;�1�R��ǘ�;e�����֪�,K�=f�M���B�z8�K�ۀ���!f�ʭb���<��X ��6��b��.+-�+$}V�ƻ�cK^ː����Ux��L�Ӏ���=UKcG�4v�r!]T5�c��觧��-ncl����]�[E�g�~ws�@�yB�iQ�d�6 _�G��o��h5����o�Y����[LL�k�'hr�
�"3�Ձ�ΟG`?]�1�%~� �:H4N�������D���4�.[�%d�6Y��¨O�x��?�����xq"���b6S���ń�O5�]60�Ȓ�
�)"+ĵ����L��u�wU�n�7D�a^��i�h�y��L4���~����3b��j3����i�S^�������,f��'P)�Qu��c��У�z>���*�^tcjaWX7s8[nǓ�j[^���~e�Ao�Rj�!��'�����*����/��G�I�����ܶ��S��|'Kt�X���+�.�`�nҭ�*J���i�s��GzB.$�E����l>Q���<���4�:*�)�52Ɯz����	@B�
�y7��#��P.��/w�S�-e�J�'4�J�r�x5�7��N�����1�(���F����Wtdwā��.��\~�"u8�p2��Y�c��L�1,���3\�~�P?5Ej:��@�V�M�h$m�P��Q�+^A��nh�� ;�:��2�����aʇ��>���?�I?@�>?m��/A"�?}��ՁDt�-In�̋��<���S�X��]����Z���P�	t�6�̉\jX�4iۼ.�	~�> hX~͏���K�%��Ѝ�M�Y2��`)T6�ܭ�Oݖ%_f#�����}��{?=�N��3�`�5�>ow�+^1̸���l!Y���F9�3qʥc}.D�H��8��T�t�/��ؾ'u�^0��$����3y����@?�I<	�;c ��U"�P9̠�#���`w
�����.�ǩ�x�j-�W"j��/��)� $�k�_�C�(=�/d�h��Ʋ�T~�G��o�g4B��:����&��w۩����匡�Z�Lz����d,�����.$Y��*ד|9�Q�D�e�e&���v� ?���o˅��S1!��
N_�S�q�vI���lW	V�Q �d�Vu�T��A��& A.Yy�/�Y �Q��;	m�E�A��M��d5��,q�n�Ҭ�ｎ��]!�!��aB�Ѻ���7V�M&b��ΉN�S�o���/���͑��`�}|`*���5 ��]� �8C]s����~�&���m���V5̋�����%���`�X�������+Z�!M�ٯ2,���Ѽ�E�u���z��T���öq=�pUy���R��e>.�ÙI�3VG�@�ğ������Z�����o�/$62�-����ڍ�A��1a��b�P��mkV��s������~�y#o�G޴�m�����DҎ|�����;N�Bs���z �'���mnp]�d<G>pe�H���13�9~�����Q!F��A=?v�q�5���<������
lg^�����T�ef8;�<�s�>t3b�p�F��G���Z��(˶���-De��2z)��}�wHj�f�l7E�|��_ע������F;\M?E�D������#�~�jc�C����Z@�����t)�*
4��#���x7JđyR/�9�8����s� ���~|2��p�}H��3
�JwOUI�7P��i�3�9�q@�#��eJ�.�:�aH��$�3󙥂dd�\��	�i�~I����OU����m�Mq�J��TT�!��{��\��lq��EG6#��V`4�[�E��j�l��B�+	_�~�#Z�(V�<ݵ2|�ʞ��%)��=�2���1�6��:���o���%E�c:�+*��`�C�vU�5�:^?弰��Ί=�4.�c<f��J��"�b�>p-�"5�YK�4l@3��`��Q����,ݑ�̮����C ��4E8�\���)����c������lQ���|t^x��]J.]���}(�4����d
-���������.�v君^YPH������Sh7FÔ�KP<Ƭ^4�#�� �7�l�Di{��Ǭ��TV���6�%�2Қ⣕ ���v�d����!	�%�ԧIT�
�b�"dP.���.�`�D{�	��<w<�\�֗e�q��aH��E��a~T�=���(��{��g\��Y���좪O�-
�ic�q��F�����}���["&Ib��"�����z��'�/�T>���O;�������rZ�K��L�Ĵ I�QgC���2��VӇ���(�,�$����Q�`�ɡ��v���ߑߵ��rK����<!�7{ �����*c�8'�����]���ȡ��a��-*U���&��`g���8ްK!�׬t�@�ɮR�>s������t\��t��ݩ�fYf�"+��|ϓP[�$��&;0�5w5��B&l<vS��c��6/���:qbJ£�x���@��dӁ��l�t��+��0B�VKŭI�[ ��&����!>s�w��3���b"�C�*�>�:)1�`��qL����/�5�>�x��S���F�WH޿V�I���v�М
p$Ӭ$^|���`�Wκ\à�ӥ�E�-;�aH��Ux�g��X~����?D�<����$Ǌ�^�$W$qձ�����z�y�=����$�����!JF�P��2����9P�謣�o�s�)1��TpW9dY�8��d��i�\�}<'.ETh�����6���:�����3�C|����Ui5"MeaǏ��d��������T�n{�}�!Y8�p��i�ӼR3� 0�ӫ��]�;
�L����?���y��/LL�XV�E1�Ԑ��/�e�d$$5����U4_�O���W)Ѯ�<�����@CA1Q�4D�dd#��$���-��U�Ȧ�S��;Y�<���R� �Y��%a���䁤�P'���F|<���G�
��c��((:��8�N7m�2,���Βj���G���2��٤�_!�2c\�߽e߸D�"�-ٽ -J�cB��s7�u��&D[��:���v��g���d�{�������޺a���o�"���%&�}YR�d�9#��"hΜ�
�y�]��\	��4&r�K}�'�;�JN=��e~l�T�}������U�3����u���ڹi�i���u� >y�Qt�J�UΠ%nvd:o���OO�dl�˷�K,��\]�`g���i�P_	V�V��̄���l �X�*��'�#�+�0Y2O�:�64a�vg=,"��}�{��V�5I_�@�����ޠ/ӐU��!s:\��P��.�g��V�����͉f�����f������ȩ�<�rF� m��٢x�6�A�l7;y�!���MGA������7X(�T�l����= ���o>a�f�{��(����]G��C�͆�B[i�$bG�Q�l��#��Cb���w;��'A�h{�aQ�<!�ޗ���^'6�����l�}�'�E���Z��|Cd]�M䢖a��k�oR�#Wos�b5;s�����9:g��06����!J�`0��䃫U��Nϴ�?t�PQH�T��^�JW��#�T���������IgS�H	�� ||��Z�I]�+�2�����َJ Yr��N����1�e�^�H�/�C����H���.���-��D��-�`�u&����^�q/�{:b>�M<0�<����x��[GInf9�M��.����0B�0䛼9��u8u��$���>�keڶ�&�^4c�sw����=��W�e�$V�3�Y��T�u!#�� ��S�S(DभϱkI��1�zR	��)%t�N�]����nv~+�b�䯎[��*�o�p�v%�>�u� �~F�#���`n8��(� ��'�1*U���n~Λ>�i�vJ{Sj��QjW�^5�; n��[��4�=y�t�N���a"G��kBfU�6Z`��Z��?����O=y�[&�M�����5;���04*v�C�T�񗟒h=�.�o\ɸ3G�[���e�t��(bk5[�p�x�^1���<�e�V���/jV�9��k|��.��o�����"h��Х�R)@��_�F�Ï)�S����BI�`�Xxyb�H�����qtw4���6 /��w�RH�s+ڣ��1�h��t����H���Fb��+3��)z��@��90��1��UR���o�`]��َ�eAZ���'��h�̲�(���O�
��U~/@��y��k�.�zN=�z���8W�j?OTiZ��:@6C���ĻN�t&�sa\ܜ�w/�s�HAa�ܸ6(R�����Y�g�%��u8"�,��L�Bl��<�rab#���+`���ly��,L���^�(�zuu�H�����Qkb,[�$����l�+co� 0- "P��uZ�w�0i�{�s�N��a����	�鑖�Co�"�!���;��c.`�hPS���<���<Gɲ,/M��c_����zmr,Ok���M��[�j�~���"��Wp1 J���$5���D|V��rL�*),�I����K�ߚ����gj&�ܩ'B�	�<}����o��y�BK����X���1zח�9H}�r�p���E��M\�)mٚ{�[LW����}, ��^)�����` ׊	X;i
��V�n���@V�� 5��y���]a�_Ѿ>U���i��K�B��/���t��i���΢��'Eݤx��{�+�pp B%-���dq'�
��P|z�-(yzXNȗ�����Ñ���%���?;Tu�X�u�c��7�*)���g�l�ē��ͿR/�s�?B�Bv�=5ӧ��g�$�~�!{����f4)Qy}����$?%y��\r��Q� F�4[l$&zA��.pc�� �b+aST���h���D�����z�פE�C8�Q#�ma&&U'��Ҋ[??:��}g�{OW;����~�	}���u	+c������꺐��ɔGE;Jy�-���""-��Ю!v>vt�	�����݁��9H`@�#a|C̦�`3�@�94��j85Z�93�Z�j+�����M	�s��x�f�}�{��oȷ}�݄�ҁs���E{g�_���1�/巴��T&N�I� �`�ߕSB�ܗA�u^�0B������l����Cbqm�
y�