��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P��v�"<ߞ��&'��k%P碶�R�ӣ�sĞ������FY&�7������pDe�@�@�ػr���#�xsD?��lv%���+�wp���b��u�U䈍h�Z���=�Q��	�Wk}��ĵCL�N���t���&�/nlg����!n)���J��e��P����GQk��lea(Ժ{xS@�euM�҇���;0Kؿ/�㡥x��@��Cb��)�'��8} 5/� ��`��ț�����bu�8��|�^V���",=>�|�5C^�MX��s�q$?OE��Oul��-M�$������wT(��V`�")�Zǩ��'�[���3#S��W��&#	���yB8��F�>�]���\���ɿ`�����ju�n��Ya��<5Vi��;��gS�.�.�Cu�OSi!p2Pڢrܦ�]�]US�Q�OK�qu�cG�r��x��ޏm[�\���rx����mL��]̢8�B3�\��oY
����`�Ƥ���o�	>����?wA;h���}E��Oi�,��e�}��bB��"�O��m�s:��3S�;�v���pv��!�d��;��Ú�jrv��ӵ\�!w}�+�1~ �!?,!�exr�;�xn\��6$>�x~":'��=�� ��pX���h'G�2�d�>�(�UY�hx�L.� A�N�b�!����	BޒG�C�����T3Ѳ+�*#���r�������3�c����ߑ�_�#��Ҡ�O��#H;�#jCZ'��0�qQn-�h-k\O88�i;h�>!Q�����y��D��`�-��CR���3=z3��;�%�s�$I�Fo7�|'��a��ܡa�s ��[*��X�"���I�kE@G,Z���O__O�L]�M�Z���`��6ytfe�/���D7r~�:�z�E�.w�@%��(�Q��i|�������-c@��9k�綃��ގ�����L޿���j�E$0L'��� ��]]���SUDs��4�IBX'l�1P�?�1>�����2���0}��";f��dm���W�zu��7����t��OK�@2�EȽ�#=Hz�(8�z�X%Z����8��+<����RV�+�2��3���|�2���G;�U?>�j��n>���M3U���٠���eL�s�Z�M�;p
���Բ�[xB'�k�9��l�q��
�)�r��O�p\X�>Hf]���h<S�S�4n ��6 � �֕�׿H:�3��7���I�V�	IƜ�Sm.�q�" 1u"g�~�*��~� HBe�6�4Sk����W�ܼ6*C�,*�I6�͐P��L1.�s���Ù�݉W}�Q�cT�[�~bF�l�k����n������d��`�6h��D��4g�!��1����Q|�"`��9�h�ȹ� v��Q��!,�?�Z�n!\��mM.�׌2������F�������=��L�bh�b�g�ag��gaXxo�іN���
��f�I��xzc���s`B����<��1N��pӯh�/
*W���r0���4J�����XYr��QQl���ء�\�0��N�<u(5��Qp��-Dq�"e~���R�����h��FHMm�m�'���'>^>�RY>̿~H�v4^~��pU�}���S�ʬ��"�>��R|!F��0���ySϴ̏�H������x!ʆ6.���p�|�%ϼ٫_)���O�g�r��)�+m�Q���Č�B�~0��m�ׁ=B�`��*$k��X~-�v�O��87O$���$IBP���F�,�.l�`��k�kڝ_K.2��M���n93�sB�љF�'l�d��K�i�s>��i�PA��FϘ+�:���� ����e��(����<$7�*���yN��8�J�V�rCk�THx0����R�0� �ը͍1^��C�7u����Y(�i�g�D$�+cY���2I����0n	��X��P*D���acc@���g���O}?9 YB�ZF�'�W��Z#&��ܪ��z�z��	,Ӗ��bR�mu:vF��J�?jp2��1Z�'ŵ����/]�9d	�N�W;��r�w�{9"����{\DN�a�r��ڊf��a+�CR�${V�nb8��̫��7F릱�@���m��qN�XT�|�a�I�3j�=c��ņ�r���+(��L���������!= �w�o���k�_KÜr�&�UCL75S��˂�M
�'�ʵ#M��"�R��	�E�گ5�q��NK2���8�|����'l�	T<)�1ا�`iq��U���E9��9�a��T�9�-G�I�/yZ���lI86��]��D6嵻�S���	f%�酡%Z8D�oɵo��XFC�;�-�|���En���j��7k��ї�c2<��EH�t��a�v��=$�}ezܒU�0�Ƣ&b/W˲���"s�$#�AG��s�O[BEz�N�r����z3�t���3��P�3DV�h����ulw�K1Q�X7�;�W)"N�a
���*jL���|ȾAd���!�6���AO�uV�I�-�"D��	����jf���SM�C���ٵ�5 vt_��Mjs�6�?x��f��b���+��o��K�9��/�.����	H��|��[��o/pn��l���2`�����D����Y/`�� ������h�[#�@��"E�p�l��g)e������/E�8%��g�>cRf��t^�
w�y�[k�c��Nok(W����Tlo�:C����jz7|�i�v��6�=,J�؛^PV�4�����{tv�Q��J��9��B%?�:<�ss�,�ӪT�ۛ����0���$\�[V��u�3�
aPU�=^&(#�d����#�ܠ�M��U�J��~����J�v1��j����1iA�K5)�#	�I� B�-ƼP.���Z�!X�n���]1�� �4�cf�Ť2{�w��0�gsJ!~�^~�{�r��.���)�=i�M���N����|���Mݡ�CG�Bs�F�a�VOZm�DK�o�5�l��Ōy���<h��Pj��!�����#S��<�1I�7֬w����j�6\�:���$�EBǼY.�9O� ~ �"���T��^%F}�ߩq�WN(a��)�	xcr���1i������s�'��
�]g