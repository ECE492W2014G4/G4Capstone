��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P��v�"<ߞ��&'��k%P碶�R�ӣ�sĞ������FY&/���3�5��0���Bd�7Ѳ� ��h(����O�)���Ƨgɴ�I��PtK׈*k2g��W�Q��������?���sP�}[Za;O8M��H�X�%Rf>k�(ٟ*���#kBAa� �б�4Ӷ[���7i
!��'7� a��Z�_�OG-k��<�a���ܸ;���y7@ԏ��ԃ�����l�����z�f�ŀU�Y�Ժ��g����Fq�ɞr�yW�0:���o�w�4��on|#�0�]b��J��2RH�:‾��v'i������E�H��]�Q��zH�'^=��[��4&lEk�h���Q����&���q=�0�~J�Q����=uS3�4Jksp���{�Z<Z.v��	�9'�00�<=��I�EjMYE�	���$�����ᅓ@�����A�f:�l�����n�iMFL�B��ׂ@C�Y��ͅG�& ���i��ک`����UJB�e�p��ļ �������ݪ��^3�wDK�C���(zY'��O�U�W=��* �W���af�B���cQޏ\[��E&b�O%����1�gkE �,�M^���a�3��G����'���r�H_Έ�P��~QEGI3&<��$�ϗ{����(�0���vׁL��x�/t���H�谊��K�̉����Mv��m�lu%�[~!D��w�znǿ<;��nk�g7{5w��O��u�a7|)Ù�����2���j�c��	?�BQ>��B*�q}�P~�`�0�Y_����X%����Qۓ���I��?�*3ϋ�N�Y#jJ#��]J׷���Q�J!CD���0`�}�0�ҡ����	Q~n-��+��V:$�r�>	i����YQ�ح�/:.��6Na3�\��u	��֏��ic�؞��3uу(��Z�/�_L�!��s��|b�~~ȶwo����
��9�4(b��wb�槦��~L�|���W��WOA�?�I���<����C�3�B�zͻ����i�_��2X��|��G~*����V����C6�G�%�Ğą����:,����	�9V�F�2��GH��#�'2d�Xa���p�����\����X��(�Y�������Rw���=���w~��!��:�1^S���nSy�mc4%��Q��A�v�>�e;�k��X)+���"/�1��q�����+U��K\W|�ަ�t�:{yɏG���X���`��U��Z]�c��|�)������F�\_ ��p��V���Ei��H6q�Z�y�@�����̐Z2�B�Mm����T1�m/�ļ�o���9N�ƈ�@�18+���AS9՘��,
GlTz�T����/=�;.�13�9��V.�ģ�����nc]�e���c#�e�_��	�]<�� ���9���:iכ/�r3g#�2
�e+�v���I��%7���,@'	R��[�H��M�1�p"�Г$��梩�r��`��y�T�i懲��<��v�o(��m�ҙ(� �Y捓% cֱ�`ߕc`Lœ��:�܆t��<��[ �� b���L92�=�&�lַk|���Fp�*�8H9�[%�_��ΪP��j��ڮ.�['u�y�W`..$�������[���+z	�
����c���ü�F8�Y��H��]VM8L��y{jf���2��~+���g��������e�4��9��	�_WA=Dp�u�+(���0�⎔W�<R�[�:W�_w�+�28%Ol���,���_�c�!�gf��f�P8$�&�����Kݩ�`uC���.2���R ��~'V����)�cv�=��1D�H���56�ߌ�NZ&�r$��4{��@�)�{��<����GKѨ����m3�jr�|��?�֮F3E���6vX/��;��$�}m�rU�^�adsk�?��(��V�l��"l��y僰c�8�G3Zd"ȃ�e��=@e���#Q��p�}?m{��Z����a�O<^2>�	Sv ���*K�mi�ZK���ѳ�~�M��:& y�ƻ�����r1n6�,n���X8'���T������]�� �����w��$ן2� �I�9��ҿ�+	�Z/*U����M3����{��s��3 "���ԋ���$�sj`�1��.7��������VdO��3QK t��18 ����7�>%R�]x4�>b��y㡐;��d�D���~|#�����?�7���7eѬ$�n950-���r2������yДz�A�U66��[2��y�=���i�|M��^7gF���f��+�,g�Kt�J,"�&�W2��}a�N���+5՚�>J�S���e��B�!$x:up�h`�+��*�(O0+:�p�ap�Q���2/��[��@Oze7*v9�m�o����;�'Z���M�l���W)&��E���E^���9�oץ�.̫dd�Tsz�+���8,KJ��Q�Q�9�eRW�+�:frN�����L���24,�o�a&���=���?G��D���$o���I��rzU%e욡Ir�]Iq�ިz�c���u�
�Ud6܋���\�W���7�����u�a��5�|�\���3�G�NF�_�R����Tb=�$f����gI�G���miA���NJ_R�U�%x���rXn[Z��=����4���I�	i}¡͌cK}`5�;��A�����o���m
%�DQ�����O��n�[L���Ic��)�dT�,�r/�C���𯃒F��X�@�h��~��&��5}��>��o��Gj1ߒ&MoPa���p��i,M�D�:�-�L����S��:{C�R�t�{W������(��4�9�vuXpkJ�ʮ�қ�g�xԹ� x����a~wb<=�6�8�|��."��8�l��$���Bc�@�=�dw���%�:�1���&��ҝz�S�*��׺����[K&7�%۔�k��Q)Oz���F#ʪ���H�<�2ͥ!�@�*q�z�'ݹ�+�U�P�w�
�T@�+��>S���	��h`I�+�!7#��H=�P�d���4TF�;'�Ź�<1�=��K�[�`��K����$�NX *�����$l����L-���@�3�9soƜ�Z����b7?�Y�rD�䮕<=�C�]��H�������4��ӇkhY����7Wo�����g��r�b7�n��{a���[h=X@\�U����N����t&D|
�v]��t������T��ֽ=8�s�nTՃS*�-\��{V@վ�boˁ��� 0C��
8�Q`}̾KT>�å���+�k�A�}��oM���[��5�v�l���~IMP!-����r&�֮� d[A�� !uoAW� �7�j��1�%��w�jm(L;r�D��u;4�3�U�P��"�ߥs [�4�Q��v2�(�~S��
�Q���h5l��{F5?��iB�A�>�B�
$�EP�*�UQʾ�e�w�d�[�h���!n1?���Xn��p��	��a9���F��>ś��i�pa�K$S�I��5yY��в�u�<��0����f�rG�ĻD�����k0�x+�d߀S½|ُ�z/�K�fbm�;��*��%����^��h�"��H���:cg�\9�+�'�4�xdG��'�@�z�t��� ۭ6�}*kp�����[�)l�5$Y�-�Z���ܯ�����j+����%�|>{��?�L@�u-�~a��};���>�ϟ��H��f�ݚ�?L?�����ZBUiU����f?E�T:%�(�Ҽ��-ҹyB��W��1f���&�|��{�ɂ��vǅY>|�����H��sb B����!�>/��H^9?�m'����'�'u�&+��Îo��]��̰f9M�F���u/|	<�qC�T��'��1���������X>v �>�����N@�^��1fx�G�r{��rl�xP]�kS�[��q?\������#�g�s�~�!:�4~���˦����c0vXa�O
�����x��A�$i�+JYz��U�F��u4:���y����(��[˄x�<�y�yټj	�ҋ���
1Q���q�W�h�� ͇l]�9✥Qbag{@�˄lq/��W�r�b7� ��M�eA�g���W@��H 4B����Cͽ�|��d|Wy7�E�v�I���K[�]g�_oOp���b�;qj��{6��p50���&���?]�[l�Me��ª�u��17���7��+X9F��6��X�����#��Q跳z���,�/�U��$�_�=��k��jL�U��M=D��si�Ɯ4���z^�ۯ����/=8���_�M�G��Ƞ��/e�d����)�`�Ԣ��&p�H]�7�����v�xt�N�H ��d�o����)7TO���-[�p��E�eα�A�"�g�1�u~-���ZYYy��Y,�� �2fՋM�(ۢ��@x���� �~W�����Z�h{'�M2KH���J��_��]����1� H�i�����Z�z]�Y��BNJ�.�j��^Fv�����T�o�Ű3�,.�(�eݬ�O�rZ�P>��U�V��١c$o͓ې���М�VP^b\�>�P(��Y�Ng+�د�����\ز�D�PW��Mr���0�d
��0ʣ>J�A�z*:����u���૽��323�<�*���~���QY�����ٛ�sjQ�LPT~ϫ+�axIA��c�u���'LNZW���l$	~�U��5E/�#Όݧ�F\�zZ`;�tnфY�@�`�&��ũ��x��/������-���v'P��U�`ɏ�L��t�2���8�s���9U�����K�K_�h�\A�\���y\�B�l��3y�rK�: �/���.�����e�T�U������f,�o��C�a#������.�+H�?��}�m�
>Z���4%֚�[@�6|I4��9��L�Q:�ԥ~t����GB  (	d�.�%o�*b�塗TS#���=dZ�wQ����a�~��J�e�&
c�6�]�`+�p!j�(�N�8s��H�*��=U���])��D�l}Xfƴ�����z�l�� �q�\�~�������n�A�[}*Ju8�n�dL��R��ԗ��1�A�ַx8�Нs!o���`��H��@����×�Rڒ�J�������7u"�;�{��~hQ������Sr��G�Y��^�q�&�M^W�[�>(��� ��)Lvͷ�x�O���>iӛ��tI�;�ĨR��HF�SX�>J��S�6�{�Gr�i�����l�L_��j���&���A���:2;��tB�?�������T^��V�G�|�#6���vm�S���z��FG�"�	�pi�ʲL%0�O�>�0{�k2�d8�d���t��	G
�����֯� ɽ�����	rr��C��[#Yx���������Jl�w�X���|��������߱�Y6��-<��9��_�~�X`�X�sdK>3@��!~6b��Ԫĥ����  �^����*{��j��[���8�}}�� x7�h�ÿ�w<<�/��=���a)��C���R� d�x+�GD�uʃ�ם8X߻�i��
f���T!n���k�Ѳ���]���
����e;�� �>�V�##w1���7�=eK�*l���k�H�%.��/�/�ً�W�1�c�^ҕ�*c�8*}̋�����⾺�f�Z�A|��5GG;oEi��J����X&h�Z�|,�4L��0u����$�9PV�}�Y�T�i�9�����A6��3/��lMѺDU��o0�#�Y{����n��K�@�C��� I*���f� ��ù/���G]�6����k��4�� �C��#�Be J�A㷼���D���_������AM�#�KR_�p���G:��n`Nd�5x�A��oBw#��ӡ�P���%�1�f�`��� Kl*�qUk/]0u��Z\a+=��y���(��b��7��B�5�I�ffB$��cT	�g�!�Y�a�����+����ҋN1}�a�����v�(�	,��̄`;��WjJG;|��k�ʙWT!��P�?P�)���p�e��Ih	�w���2��_���(��^H�T]�(vr�p'ExWh�[��'��C�����1��XW�,��lx��j%w�@��u�N �]uN��t�k��b�[�k6��wGW�B��ӂ[i�:g5Y��y碊q��v4��!b�x��#o�/��$\��y��F*�*�H�*N�%��^̏�YrZ/��CL�6�fܪ%o��5���o���[*��:�	_r^�=@���/���V���j�S�����3�Hq�4=(��f`r(T�'w=lR�g�?�>��x�
�ʊ���nt�9n�F�tg]F����'Q�� jL�Fqs�<���	���҇KE�Ի���&�3���7�����9����z�\�a_Z{���s
���u=�|�'ˋ}<pN݄��9�O*���!�h>q��X�y�jeLy#����JU�Y'F���Yl���5�ĭ�<5}n�ǉ�'m5 ��?Lk��4�E]�w�?����v0�N�i�r����w�d��{���|�~y��\�毨�u�������^L3�qj�j���^��LS"~���JƘ:IAo�5�%��	�7J�ZDu����Ūk �ZA�x��_nMWp?ZB��T�;]"��q�e�'pfү���"6 �|���6��a�J�)���r�CG�5�_��Qm���G0�p7�b��\Ӵ�^m3}�Z����'�x��l�V9�8լ��Q����ȦUm��A}�[��=�=Me���� �sf�'kx�N)[o�y>ܽ����c<�lRh�NXi2R�J
?�.Ԇ�;!ס��_"�뱑�7(k�����Γnߝ��[��3�o��)!� �V��	�59����y��f/�pq����;��F��;�ي���bE^w��A������]��s��[�E���ڹ�0���Ea`(�=�/t<��j��% �5�}U�3���y���_ˡE1��v���^����k�?h��2����5�b��υ
�etC,=�SB�\�S�݁��6S1_�7���ʰ��^c͵0�ą$�� �	LY3����$�w���FAy bj��0��ǽ�G�7YΙ��b&f�a��@�[�+�F�V�,Y����ɰ��:+J�`�k�m��)�Z���#y�jWE�z]�׷�~�0��V�A�5(��:���O�l���-i��c֎�\�k���:_Ĕ3a L|-��W5>[�g��+�o\:�	J��i��s�{	3	lx�c}�G_��}�*~���q۱��_��)�LLT�uE�Q�����C�t� �� w�S��R�J��ZO��I��x;
d��^��+�D4�cj�R8q��.b��-F��&�p|N���m4B׎�'<�I��?ssK}�|˙���Ȗ�dI0SswF�k��6)
��7W�'�]�{�)Ab�%�e3B������|��������xɹǥ_�F��<����(%�q��J��❺�e��hCWzZn�}�c�9ҟU�$_?8z�6P٧5��hѿ^��Ǎ�1�p���x5��z0TI�[3Q챎���g���s��N�)	�$a�󒌘��K���4��]���O4����4q-=�=�]g��J�'g��O.���7Rs��
����2�Pk�Kn�����~�b�c-D���D�ͼ#o;�˝��G=z��/o*I��۹qm�!�%C�Ӛ�t���M��88�돝
oo�~-	{\ #S��[
Uܸ��o<]-D����6�����M�Q����$u�_�j�5L�^V�>��TR��"	��-#p�NH���ul,&�}8,F�w�a�_�֮%yz��Y9I��T�GL���\�h~�^]�a s�����k�^Fd��}������}�j���(�<Z�$�U��G�x��Zl� +:�^~5��q*jz��q� QD�����7���! �C�Son* s��"�?KRҨ���7-U��l� ��D��x�PdjsFĿ��_�5��l���B�Æ��i���`��Zj�
��I�$��"`&���� $�g'r޳N�$�cN��)�J��Q���i��з*	���|�x�v��~�#礗�y-p�fW{E"���6O\���M(��-q��\�q���JL67褬��'.$[�73�P����u���un���cN샽z�E8տ��&`��Qт�j�L�C���6>"����.�u�Vʒ� /?�
��ܽ`{��&�ʲM_sd�H"2̖=�<�!E��қ	�G�+�s;"=xL�a9;�.�X^qh����.���`����c�����'ˌ�q��4��J������Z~ٱ�bm��]Э|�b�a��B�*�)饾���y����$		]T$A4�
��z����V�(à}��M���ZC}>�]�[�޾��T�-�h_�
� ��ބ�	���>[��43L����MpR���I�F�9~�p��N1KxO'�*2�/�RU㷧)^a}�1e;\��Э�
���+nپ�.�f��x)U��)2�ڎ����IN�N!=���x(�0��R2��o������ l�=uwN��؉s�� ZT��j���֢�d�J��o�U�-����=n1�2�/*KD��($Dq\L���f��v��U_�6�=d�J�����͝������S�a5l>J��J��X�-"ɳ�'6���ei/��j*l������;��#p1��͡�;#!�l:$�Թ��h)^�F$���Ԏ��^.x�&�Cux�����ʲ��6i�]!Ռ>Ы�|_��СK<j�u|��%�L����%�7��k����<;(՗�� w�a�jY}�" �����g}�&Uj{Z��U{T�8�V��a�C^F��H��P=FɽSE)��lj���t�0��i�a�竔�x+= �H��	v�5W&�YM�?���A��C��Sd��+%A(�̨� �/�g�\��� ��Tpw�ZA-��y������s-*���,����K��z�r#HO�<��5�O������8/�X��!d��A�m��$D�bX+U,7��\1��*�ܲvI8=&�l�2|ݍA(e��
�sѧ�ݱ�x`�KwOaf��Ow��vd��o���A'>,�|_ܬd���!�gˠa&���r���u������o�!z�f��Ψ l<��f�fZZ�p!Q.� �iA���d�- ~#�My������������<>��WL	Ƈ�&����/�v����`�^����]�Z��1}.H|[b*Dm�A6��X`�/��������-�={f��D��ǎ����lL˻V�.�ae@�?���!z��!��d^���$�AP�__W+��*�O���E��[�r]���vﱝ^RdXN?o��2{�K���ݾ8���?��$��$��u�WZN5KQ
��k��7Y_�����s�T��q��;���N�e��nK����Ɓђ��l��U�JO�)��O�dByY�E1�7䩱B��ԟ��=^���{�5�?6�^�u�&V;�$�^�������9you��M�գ~��7��bk�>p}��� ���|�:��#/V�� {�X��īSң�,HL�?�&Ta�7Ľ� �.��h7��Ɠ�:�p�^ĞS���b5"�chep���GY,d�9C���b8f��l5l&�[d�%���yɍ�/q�w0)����0	�ZTƘ�D�����F�c_���xj�ٰ�����x���r��`M��POe��J �.��_.]�@�p4����,n��F��c)��QQc�E治5%� ?�ڰ+Eݗ�|���r��ͩ����^r��\�����qGEy^z��x�޽]D�[�U��@z�i����-~n�lk-���g��rH�ZQc�`�4Ey+�|YE�)Iʘx�(�6��Zd�1��f��i��M^��S�5�Èo^9ֱ�Ðq\[���:Y�`��!J!����]e�9�aw�M�R�-�t��2�V���{��Ƌ��Y(�N�/WN��q��d�G���y �4�&��`ZOQ�q�r]�~�%K��{���v�D`���6�����jA���m�B�o�>��d�V.��)���!���d@����@�B��n<MH0;t���Z������ܽ��L�n��N�4B�ND�o�!:oQ`e1�Gy ���W@�)�,<nBF�o��g4��6q�h��+c8*����/ұ��»�b�~��Bx��	�sLRo�M":Ш�������h�a�;7�u��q��5B"W�%L:;��`1�#�o=����M�7r)��B͔Wu��=�9�ʶ�R��`(�"C����.���K?��zSgX)�f!u�n���� n�DOL���Ik˓�F!��]+����7�G�P�L
޼�4C�����r�Xr��pZ|-X~�����#u�:F&j�ӗ-ж����M=�-�ģH�^��̷����wE�h�;p`����Wf����]=+�37���G4��ҫ��26?��B�)���MOA��x0�Z���;RP��qY�Xأ�\��ږ5���A���[�=?����ػ��jJ�����-��5-�ɏ�t�*w�����q��q��i���w:�Dn��k�I8�����q��/_u�v�4���7��wr�51�:����gby"I��	��[�*��f�q��̦RO��n�r=�nL����bA_>��E�d�ǋL�Xb�m���'��_�A@�ERkn��v�>��pb�-'+��܂�؂�D��!�6�S�V2�p1P�c�r��"��TA�-�p��~x���xl�$��;��G�e!,���7����0	�.x��F���uC<��𕶐GsO�욁��v825t�@��=A�������6�^�e&#��r ~'`8M��Q&�ɏ��/r:�T~���L��[�����fs�☏b�jm�P%y�5��&��� �ᮍIyZe	\ԗY=j)lB0���xO�~�9��]���`B������+F������іc��嗺SS��͹��p�!�i����m��_���.�n�d�<d�u�#t��x�"�rmdC�%������F.\�9��!��a��Ҽ�jJYZ>��2���_m,;,H�"��k��g��E�i�����i9Cם�^�#w��=K���Y�GlV��J_�x�_?w�}�RF�B�Q� �-��p����nɟ�i{>��
.�#��� M�b	ĉ��N�X�Y2!+D�1Tdl[��e�d}7^:[�$�0d2���+�Q�.;xx�zT�L4�a7��?��4#��D�bm��]��y�U]s��1��A���M�����Z�FF)¢�Ȍ��2R�'�CT��^-׍�#�w��U9�@�9!Q���P�l���d������H�����rq+��@?��7hVZU�y T�/.G��QY��������;*5���#��ůp�'���"����� �6V�����t[�S�3�n�G���(&� ٠9nc�ůY����;�.;�8��ȌE����<��PPզ^<c�cz�q�纅g N��Ҍ�L����d�ֳ��A�����"��Z�rp'�4��?XP�c�w� q�˛�ό��Ԅ�T�0F�PF�jB���R���:�U�)��ז���k�`���#�HEKl-��/cZoVu�3+t��D"�De\ȸ$�� �I+���'��;b�jh9�jvE�%�W��hoN��F;�s��H�t��ԶB�q��>q��-�2���r���9�\��Y�����͍�*�\��"!Tw��X�5�F�6�����J�+S"�ǨX*��k�]̰�Ka��t2mG����~�`���:>M޿�{�WR��6T�[ݓ�;��R�A�`�=�~���M8�%��:ա4��Й;h�7WT;�z�K;�FT����SY�^X�9��9NLG��-0��8�3΂��-1'�[qK�7x-��bJ��>a�S��um�2��s�^?�U�gL=��6�����e�ݨ��-��8ύǌ�)���3�5/Y��TE�7�'�a��ߎ�%����3��n��59����X�];f�:��*�/����'�μ�J�\c�a�,2/��뺁2`���[a*\�bh�F&���G� ڥ�-�����!����C5K����p0�7o��^n�7Qw����W��yt$6�H��4WK�zMO���e�ś����?��)�ӛdI��vf�]J��f��i-v�W�D����Ҕ%��f�@�j:v�]M4+���y~�l��u'�ǚv_'MC�Y��R��EEj\��g�xn�B�Qc���C� h$����j������S�f������S4!J��aY�(��X0��e\߬y�03;f�'t�kv�o�2k�����2��
`����`�+��p�Ӊ���)Rq'zt;��{�Rl�.�gw��_�x����_i�>�Rb),�_<�!�>��/��F��Ӑ�F=���v+�Cr�$�G�����N���e!�X�P?!坊��[�B� m�4�:EhcLn��f+��>/G�O��zخ����=�m������ԃ��^��UY_Y��Z�յk�T��'3��Ԟ#��j�РX�tH�v�-��y�ņ2����<�s���z�<�BoJhN���9����nv�L>�S��H���Ԇ�d �:�jf��N�~'ђL ؑ�eh}?���HsY���#;���ѭ)8=��^ ���ʑ��Fޕ�¸�K�WU�GI�Up���n�������O ��nZ��Z�W���$�ip�B
��6g�z=�mLVg�HG���M�0'�r(�u+
x:�ٸ�C���3�R��P��~�SP���d�W��w��H޲68[҂F~��@�֮ +�א1̞rg������Lx��<]&I��r���&3x�f�03���y+M�e�=�"�e�h�^B����iN������}q{L����4&��N���3��h�� 3A����i���2S��V�+(b������$h���\a>�. X�� ��/k9�8#!M3�\�D��� x���p2'4�!!"�V����毳 ��x�ENqz��S/l����c;*R���9��ͥ*�x��{��T�I7�,��K���(3��(�t8c�汍�gH�EM1ڨ+5$8%)��7@Ǳ�K�.�>��<���2�d�!Y��/�'���D���=�>xș����������X�K��*�: 3����&V�&��:vX��}~�0��Y2x~��Kw�Q1�M1�����uТB�tO��{��%%�dqx��SM�펑|�R��Es�tm^r ?zh��<�O�N�&]���ِ����ߵ:�e�~Cd�C��Ś0�&-�]��u��|�|�\���F5V1+�uR�J#��Ji�J�}+s
ZT�'��1¤�=���b/�g �(^���Rk[͢����U��&�*�\�N��B?՗�wl>�w��	�`7)F����5�u$ml*Pe�r	@����1�pa��FNZ1�ɱ��$� �t��],�q�ut��	/O����#Z�'��;�������(�Y�
�aQ������t�5�L_����D���aļ(:�s��TfJ�чa��f�o~-HzK]�����Xh5��d#�0�8(-�ʻq��â�|�Q�O�� �nW�`ʢ^� ڣl]]�=�5�YA������m��v���:�!���3��B<9���ҡ�(�
�[ �5����ۘ{̴�d���9fY#��������2]0fݼ��'?��<ȫf"p�qK,��O��Etbc&�#:X���K�-�)O��۔�ɀ~�{_�6�R��w��S\2�d��<���q&�$p?ݐa�>����d �@�zH�Gh�Jn�RN2)�Q6�~])��A�V�	G�ZX�h�;x,,�S܎�T��-�-Đz:�oozh<G�f��V�?��fi�ks���`Ź5Y�.�I����[aW�j3�Ë/fƖU�鉷D�,u�K+0�3�T�ָ�|��\�v:��y㟗G�zsaĻp��5hv��p������_�e���@S�ͫL�ՑċQU��`
4X^$���-�p|�szze����G��$C�=�>I�W�d��V�lcek�H�%Z3ثb����e0�c��m�Ҹ������$�E�v?�Y�P�r�������M[h͂o�i�a��m:���;�r�o�Hܙ�:��0KLa��˞����dX� A^��S��'��u��h63�h:w�������G�4A�R�N�<%Sk�AU&ZT_͚��E����-E�&����zw����Ngw��~��X:������^��efo�¸|)�]�&�>��Ue��?Bh�}꿝���#�^	��0�`b���zD�?$ų0}-��ﱪ�����%lr�"9��)oG���S�W�X`��g�>��z�,�@Y��"&E������"�z�b`��DY,�=1����1}�����N�L{�{i���<D���c�jo��\t���`a�8h㢇�+���P��^o�jɩ�u�l���N���5Jy���Ԋ��_P��plE]�7j�ðr_�%8+�0��W���F��rŃ��}�-�+���)��n�(Z������#��qf+�s�m�-aSA�@����\��K���(�2���8�� ����^9T1���PMq�p�ea�<�þ���a�.�{��<�{��5�@�U����i�������}�9Nc�_�-tO4�.Uq^��RMJ�	g�I���?�����(�:�������2�e)űS ���kwI��L���%$�#̽�t7%���_G��3�� �u���;]���S�͕�10��mO�k�'W�v����g�ʦfm����6�:#7ĺ�*oVzgm���C��MՄEt'��k��߅cZ�hT%B��\KD��g���L�?�7r0?�gRxS��Sq��	���9�o�r��Vs�H*�]�I��T�!�t����'Oz�k��X'yUm'Gts��=;t�Z�������|�Kۘ���͂kp!Q� �������r^��.�Lm�		Z�mV�%�$D$&𚔅|VE�_���ҸY?���6{G��C6�*�� ����S����Sx=����C����b旯S��&:�w(�0"��5�X�)���7>OŸd��
�p��zo/}���/��f��ߩ>�C�������9����QX]<A�)12�莙_�٤&0"�j���A,�di�?G�Qm򭿱�Zw��e#�y�ߡ���B�<U�[ū���~Y{������>	OH>��4����# `P]0�ԎA�S�;��R�K�a`5O֫�0t۪q+�g*�0��ki�< ��?��`�+OZT����4g�uEc	�����(f��*w�Z��:F���d��4�\a��	�։'IB�쟪G���B#O�N�{������o�.��{���e�}ow���Ԁ��'��nK�QC�"�[=)X�+�{�z%p-<l�OE����UYVx�u�·mb��}����V����Ng��ȴFy�K~����A���ÍDjS���3��CfJm��آ4�#▵{�Fv�d �s�d�ƫ]Lm��rқ8�G���Җ,�D5��/� ���@	>>%� ;C�6�7]g�]k6!�!���{;g,�����A$��V출=qy���@a�����X�|��6]�ۋX#�G-Y��(���#L�VEwL72^��T�G?5�asIņ;l㷚I/�<���:3~���\�;�R�iU������R�!��J�|��4�9�M=bEe'��˵+���P����F�K7�}���<��mhQ[ꗹ�*_&�8})".�A@��iD��|@4�+��g���,UkA����z���9���ryG�����3��k_�s69޲�ŲK�5n<!<�t]�M{�C:���a4�,[��))��W����@Ԃ������H�V�R����&Z���/3�RbO�@��� �qptD"U���G��\']ٙ��S���.���GK�Y�o�JL��t�VVΒn�d���h�]�x$� F��kI3��z̑�:� �ICy�V=�t�%^�K��s�]�Y����}Vt�p�O�?��A0��gf�M	ה����⧬���H.7�>��;]I:����S��a�.&Jy7hl���U�Jei��>=�����F�7
hn�Kԃ�UE��յS�J�[�EF�3��(F"`�
���4X؁Y�,_�Iq+;�t�XX|m��c"�"����\����	mՖ;bG˴sX�.x�xF�7o�w�q�DdYa`��:q�;�؅J1\�%��ng���$�ĭf�^���g8��v����O<�c2��[�eg�tB��-<��%<��iȅ�w�uU��h�Q<f�� �YFl����1�$�=����T�}�N󀶐:���&rѪK�?3]����I�a$n��{rE?�ٳz_? ���A�K��F:��=�E~i������>^Si"�8��.�Xk|�ୡ���M��o?��.��	����L]!H���I�Ȃ��)��ƣu��Z|� ޛ]�4 �N�P�:��/w�~
����X������Iw��ҁ��W8�%�t�MZr�]}����_��&P��w��{	��s�'ȗc�!G��$�oYi���S䯕�mq���M����V���h��,���E7*�,[|h�.H�K�ln��������1å-���Y�0�ɿ�L�Us��Q����*���g;����nF+a?��:���o������)2�h}�C;K�4����Ψ�����0
S� �j����I� �YAp)Hu��>�V��e��=���<����X��t�u��ce�3���c/���=��C)�/0���
����^,o�vFA�m��f�@����	����ZȤ+@D�aսz����F��Iz>�t��@}�]�q�(�M�SmA��F�8��a�`��DZ�#����G�b��Z�5�baa����d�����츪d���*�438��]��f�4hMuf��-6�lz�*�_�3����)�׺�"��}j��$��Yp2�.��(�:n�~�e��	}��b �)?�	�=��[���.��<)䦠�Z|^��q. 9�\M&���W�z�x4l����`���=%��#v�Ǝ,ǵc-�[ 4M�G�f&�z`����"5?��F���:��d�l�����k�m�Q�;2�-��؀����vS�{�o�H� %D�a:2�x���-�Π��Y{�$8�f֔��4{f2�ˍ�K7f���'��)�e��Kd[�2�F �o��O%��������&7g���� ��i{�]���;��7�f�Ԇ�-b��3Z\0D�x���H�=W�޴��Wq�<7�nW����B��Y�2��ɺ����aC}hF���N��(�ξ�`��C'u?����Ig
�l����;�G���8p��4�L�2^��Fܜ�*<cY�<�Lv1:���h���,ⷃ�|;6}��X����-�cx���Q݃�M��R�T�!iz�l�q%f.�DP�-�}Wũ�������Qx��6븟4�s�{�~�q:ܴ���xѣ�b�p=�;���c"2�.��n.Θd���C�͉A5C)�Rg<��T�,�8`��l�D| 

4�~���x[P��n��̎k�<�0̶\���/	��|�ţ�/��/�u)·d�����;�->��>�P�!G(����jN�Ǟ}i�~K�1�6g��e9C܀00b�@����b�P�P�bՠy�gR�>� ��Z6.������V�(N
Q]z,f�s"��	K8!��|���~�*U�Ul�4^�۽04�X<ZB4Ku�"�[�#�yOo��M0�;�컮>c�1+DnX)s�g�3.�^kxP��V���W�eJ�i�� nW|�w q���S���i��m
���?��-��y9$x��B�u�V�ǐ�Xj�K�}�B*�> ̻z���+8e2B�w�3:����ԑ3<\-�"��qzz(Ik3Dҳ����R{����Si�Y7��֩ӷ����~��V�Թ���!8�~zK$r{-�;�m/�|Ca����>G����)��s�m�d㖼��1�&������0�F�̈�Wt0�+3��Y�vc��Ն! \f8��^�2j��
��4z*�*ꖯ�"��I�ԫ�R����i��"a>e>�� �5�?�ќG4���3�YɚW�I�xX���;?�3�3��ht�B��?f���e��M��(F`V�z��.L�S`*cq[���dZ����K�������ru�I3�n��#�|��� ���:�i�×�:vz�p�{zLȂď�E�t�'	6S�����8x鷤�}���mPH}��l���BO�4 SF��:fC���{V�N�o�1�TZ����=��Q"7�E�J%�1 ���z�����c���u:0$�H��h�d�_���l�ɑҨ"�`����^�ct�au�n��j��`��sf��������U�LKfAca�=��<K�<;�q�u�þ�=U�*'E<}i�R���^o��g3��i�0¡o%�?�O���2����2����cV�Ҭ�^+�?���=�;�Ԏ����r�D�a ş�͔.����!�W���qs�`���H�i��Cb}e��,�E����j�H�ϼ�Y­Ҁ<�,G����y�?�gO���.L��SKd
>��Ah�RX~f8�s��
���a���|'n��]F��Y�wŰ�u����"G��C+�a��O;��z�a2
���K�Fw�C�S���=�O��{�XB�wnGl}�������;�J_#�*;�m��R����]\�ȦvLb+,F������8S�0�)	8�|�$���{������h�`=�2�/˱���t�"�񓻭�wEy��ta/_H��mPH��[f�?IY:qr��0��2i�Y18����j�bQ'`Z�0��?T�涐��~-�4�lB��gT�=R؜ۢ�RG�&�ey&T�wC<PWN"�33�7OH�Ɲ����	m��K]�L%'][��䗖T�%=q!׊�~���3<�!@=<���҆�Yd��'j��R�ecx?Deң[A���y���	Q����D�^P�xO ��`,��\r�������]�rh��Dm��)�Њ��=4�[	֚@�I�)\�/�z1_=��4���8���Tώ�gxap}$�eBUtݚi��3����z��?)�uY���+f3��P)N�KN�,+�5�kD��%k��� Sw�� w����k�`G��d����b�(�1�UƟ
*�XnҀ�� ��%�U��I@�1bx���p�	��������2(0��H>)N����wtpr7�5���sZҌDK8$�+�)k�z���]����U>L.����'ZN��V�]�����k�_&�Q`k�~�:x�7�hgz�_���5��o�5�d2�t#3�V�'�>%lD˦%�Ն���y(�kc�{.�oٜ
W�u�9� h����|r�a7��f5TO�N>�M��FM݀P2*��@��	�v��<��K�&�z����|����:*#يw�wL��5���\t�PQ\?��t�|�F�C��=�5��f[~Q���}?�A��:�Ԣ����Ǥ�����EJ��v�%4~�����r*6fa���ղj��]�D��H>���VgF.�_�{ӻE��[�,_B8^�Q1)�ϊ���!#QFs�b�L�}�L*%���*��!�5�5N M;#�i�(n�8�׼zm��~�e��5<�ңu�<�ʻ�@z:�tە��F��vw���E:v	�{v����C��bwbMkI� �j��+��u���٭���%�n�9����忷q���]%PW ���(��D�(l"�0%��jP�v��=t��K7��bx�DϘ���b���#��>.��W�����?�@;�(]P{��=Զ�N$�\���%����������"�X�KQ6���֥�*3�`�5!9�B���:����F(����aH�{H�1-��nE�^*hi']�j��T%M�&;�pދ����r����mD	��W���<�q��F0k���U�TL�͎�>�V{�Þ���`���Uq���6Ε�=����,"���_���h����VȢ��Dݮ3�P۶��) �~B_��h���<}���h�5���G&�QB�uw9˛N�5�X{���-�)��LS�D���#*+ق>�J�o�k����6\�qgm_��'�A�sm�*��	�l={������V6���@t�{��R�x�*�ߝ��n��=pM������S;�D����B�t��3Q�A������g����������_y�Z��#mt���.�Mp\!��&�̰���hs�;̐m�	u��m}b*ZIljR2v3jufhc�n�@�_>�%�俧��~zP���w������J]�VkN���B��A�J|��aP�<�qTJ?���R^��d2�;����n�����Qp��?V%<���p�PUIp.��2�T�ѭRXk}@�;���:��r�`q�m���e�0!m\���u6���4i�tGp��TE����r,���>���(:��u��ah*��a��K������+�����2�����h�1�m
�!����!o���]L|�!�íE6���a���s�t'���r��R=����b^��7;_�s|�MB#]���c3��օ�Ha����v!�i㰮K+p�8����7,�O�Ȅ=Q:���]��� ��H� x#��n���-�b��!\���V| >�\�c��qQ�6�$��o�^�����4�Asמ�X@�q�0��>>k��td�~v�BϺ>u�b�j�d�~)xBd���������M�$r_��f��C$�0����leZ���>6����(�䁈��q���5�=��ɣ�Y�Z��h�=1��d���G�e��І��!9�'���Iv>P+^�J�ye���P�,p�,(�h����A��F��	���Zp���u9m��Q���n-�^S�Oo���oR�ҟ{���D�$M�� q̜�}�7�§.��S�ޡt��׹����[G�v-V���Nُ� ߵ�!��_?h�i�����/I�ad=2$����1��d�e>Յ�ܚl�暝 4�^�R:����`]Ζfw0X�T�~�8�>c-�'����t
�g;w�$�Ɯ��ͦ<{�*��DQӱ�^���Sz9�R!5O
[��2'Rw�l����؞�
���T�fϤ�b�8Ę25(��P�꺈,����R��h���1H��sge5]k�,qA�R$�TI@F�l.�=�L=ƨ�@ә�
��L�T݁4Y���w� P33?��a����Ի����5�y��>�J�
8���T�x��4ΪV��@<F��Ʈo����X�f��lz�Jd��9�m���. +l.�i��2����U<C���)4՛�d;���,�ݴ�r��3G�2��2)�(��ª�`u���{_YKPg��E�[�.`�ioCl+���"���|<�" ��w
�1��*=�����3U��2��)���"w��gn
�M�4���,�	1�$�d����P�8�-i��^ˆ� �������0�<����Y���~S>�
���9�;U0���Q�{	��N���c=��S��
�A���^��+�eyP���t�G���'�J0�j&baL��0�:. re+W�uZ!��/'�~��M��|ܨ�99�5sz��7���`mr�Q\�6�'��*?,t�I^�E܏���]��v�1�K�gհR=x��g9��K}��#�Z8�\��'Y:e�P.������cd�����Y�f"̞��djDFѤeg���#��pBr��{X�#UA��|A���}^/��)0�i֨����+%�)ߏ���"�Q���
��Dc(�D�!Il�ؓ�K�)zc��s�n�+�XCh��^��P�%s�����a��a��ؽb�-�+�z}y�^m�g���~+KM}���'��0"��m�n����WˌN8��N~i�4ّ9���w����(meX�`�<��F��?� ���~�0�#�*�ʹkۭ�l7��@{��\B��<d5?�s�j�zm_�nl� �m��1�q��M���"�������-E
�����{<m/)�6����$��C��S�XR���xi���i)���������*?��N�ƭ��X���M�7�$��?��B~m/s���AL[V�-�Z�eQ|��i�'eC��kmB����h�J����:�t���������/�
��SD���<��o��B%�XZlS6I�2����̲�h�,�E*�9@��fe��M�08�
�߽'<ȌP_�U�x��ԕl�]�0��Ty�ѧM�rIm��+`-jB�л}�~#���X#J�j�ͭAuW��t��O������"��6�a�ם�4_��,����r�B���(�H��'���K�?qO��}��a��S �ءEG��\��Į��>)A~��
���$/`���M��z��-��&ļ٧�ʨ�ֿ�rT�3]˲9�Q�����ջ�Ց��2����I&\����Q�~!��H��<Vp������^�,@�4T�!�]�������+z�x�#J�g1t���h��}���<F�Vx��E`]ғ�7��s���8�����������	����7�*��}�t�e���gX��X\ R׼�}��C�����( H�ڙԐP�������6E�M�*��O�]���Sǈ�鎴������UEp�_�b���cO(��8/�����\7�-:>�	W�m�[vnS��5�^�YX;x���e"	f|��bCj݈��4+��c���%ހ�����������vq���VҖ�'�j�[��� o�`!����Xڿ�B����5R'+ֹ��� ���sۘ�/�O��"�E��lJ/&D�08��2#��DRł���(+o�CT6��R�·g����8����l��Gcux*^��s'lkxy�P�˙��#�)i�@5� R�p�P�%�Y>y����cO��U͆��"��T2����qլK�#!s���U?c���<<���t��a� H�h�o9��_��4�א/dM#�}���<b�`����hO��[��ѕd�6J�
��{ �>�� ��:�*m͐O��#%��}��L�nC�œ�၏
C�t�S!.RB���W�2= 7r����T�E�k��yA���ZB ����{�����0ֲ���:���>{��}7�]�'Y�Г��
-M�K=Ľu��\���T��-����W�|g��P�C�zE\t���8^�h�?��֮~
� P	�po٫b�&�mTx�sM�����R��*�\��� ӷ�j{<�d��	�t&Q��@��֧Z���K�����kQ�w�k�E�V5æ=��:C�[�A��7����^�ivW.3����Q}*�M�8����p�
`Ŧ0���h!;�D����Gtrc�bm+j4��XIu�䃉ϳ�u ��0V?�Y�ز.�f<oP�����+�v@���4xc�	ǅt����/�!�z�3�s�rx�V��2f�	p�i	�de���m�j�b�6��ܲ����1܆�v���������s��
�|�y凂?��WIqBSu��{|��u0���f*��y8`�����b�#��XG[p-�h��Bޡ��7L�̬z�f�#�د6��]�m�>=4�N�GE��?����?��v�u�'>���`�)J�X8��F���B|ؾ�����*T�<v�A�0tm�� ��.���3�Γ�ײ��j���A�S�M��L����jS�k^�q��`�&*fX�5r��oi�\��t�+�nS"��YG ���E��X�	��Tj�I-�8��M�
��t�H��ғ���3�9��k*��"x����_B�:�v��~0��y��������i�������^U�ܖK=bai�-Ɛ�i�Q�6T��l'���B���¸gX���s�5 ���*
�tM�W�)�z�;������I:k}9�PiKE�m�J+/���b�`P�N>���Wl-rÂ�刧�]�����@|l�s>�m�͓����PD�i-8�L�� l�3i��>�g�҃]3��UDҿ;���R�g�ض�+F��D44��!4�+����b�iYs`�2áp��s �w��$�8Xo$�:a�8�F>���q��R�x��~&�,��n=�9g���/M^;�|�4k~������C?:�n���T���nW��\���,_���=��Y渔SX�$%}�
�wD>{S�0Y���JV2��97��*5�858d{?�m=�g������u��Og���6�<��dW����E�����1���q�0� Ơ ��Gy�4��>��&����ů�B����N{ 
c����.�~X��~J�oE�g��e�o�G��7ul�2BP�K\3�F�q�h*�7��]�K�omĄ��9rȁF	zI�:2���Q,�,��.��v���SfH�js���9��؛ [���KM��X���;`�b��
���CDn%�<l�zV�����s��Z��#2{]).����2��M���c"=,󂧛<Nqf�E���~E<.�c�� {+AĢ|&b�+B␳KYt�dsh`�?h��!�Gó�2�+��d'<��֑�骚Ư��bt��2�D���f�b�xK���� ���8w8X=ER���Nuk��7�!u��3^)�H��r�`3Gl(�X��U�"��W;ۣ���tP�����4�\O����w�L��|�OYSFm����
���{��j��~z�.Sr�{Pcc��]�w���Ƹ"�=Ψ4e�wr���F�O����`�1��KǯX�����u`���+��bE��ϐgGn���	��0�4�pƆځ��"���X-�4�5�,N�#���f1r���^6�P�����$���r����@+;�<��ɑ^Le�o�i�D(U��(K���i`��������4��>o�i�č�c�Yj��w�o��(_M+��>B9qDh{09�Tl��T���w�{Q?��kJA��K�/lo���a��i�`�Z������[+���^��M�`gX�D��pӿVL�E2(~5��TMޕ9 ��14�N,٦H���&1�$6��q�R�@YrY&LM��	Y�Sz�0~��xV�����	���o���|�Vıgk�[�_B����a�m玁�h�N��=����=����2
��O��oh��̓�!�%�%��6�G�ő�U9|��f8�=ޤx-Կ���G��pw���I|�~K&p�1��+"�c&��4=9��:pV�����d�>���F)f��������7SH���R;Y�)d=� {���D��|��/���i:o�(�w�Z��xg+X�xI�k��dŸ�w�vV8�T4��Rn�A��wVV�2��4�D��mҕ��~�޽��z�;��3맃��y��.���@���A��Λ�9,���Q)~3��
1���c�]u��Od:,�;� [<b���g�[~��a0hth�NQ�,�I"�G�e/1��N_���@�l�J�?�6�nM+TA�x����t�y�k5��f�˶�@�ꗇ�1Wf9��
s�Rٱ�SRw>�#k��ԾV�uH7\j�|�;��˝KR4O���#z)�L�V���M�)���|t\e�����+zn��M�ۉ��ݽ.��|��( O��2RԤ5g�������i�j�ljt�A�s�Ș��q ����C��y>U�i_8aQe�]��[~V���s�Zx7����SX��%�S�m�L�J�X��4i�mul�u��)".2��U����U�t��^�O������-�X����Pr�{X��d��Y@^��2��q(�mh��`H��3
�ܹ?�nڊ�'�	�-������Q����O����i��ev�-���f�'fpe�Na���[̺H4���.Q|��c,:c�!�Y���e��-�[���J�`��įj�qU�Z���;i�,T+�A��
K&�J(ƨ��7FQ�R��t&kS+g�"bu�O������m�Ӓ��	�l9�~܀���0�)�")����g[�d�һ|�F'ޞ�i��NĖ�mٯW��,⚌pAdN��ܒ6��S��(?[�u��H`���A�噭��{T�h")�B9k���/��$�6��vz�:E6Mo�5Xu���b����~ְt���^
k(L�|���Ye<\$M���8ȟg32��*(u����y�L �';��ڍ*'�=$p�P�6�]5��F��Z�اQ��0�P֥y�a�_#���m?�����M��E2͔0NԦ\��J�&]A_��\iV���.��U�=X���%�^�W�Q���x&����d���o��/M2ۼ��;B���!��L>q�G�s��9F�{�=Xd�.�������N��5�b�=.9-���U����2���_�j�M�v�b�5N��؀{V���[���ſ3���D�D]���!R��¹>���T�^f�wn��M���SI�W�H��޾w��Z-��bk,9WR��U�?Z"���{H�n�X�K�4@�ݏ��8J}�����&e�l搤�?Qnz�ą~{��CEL`{~*�Be�M�B{#���Cl����i{f,�C�gڤ� R����������	W&xvB�E��2��r�-�yA�����w8�[R�{���޻���B�mNG�c���4Ɍ�ai�`�l9��X�e��H�S"�1�����2>^��dt)Ȫ�29=��ti�0허�Y���؞�"�d�(��
㋩���]f�0��@��d�%}I�5�q,��"I�Ɲ�}`̛�9���; p����-	�q�~��yY�2#IC˽�d��sasQ�ק�L�*��v�Wá�Bp�[��~i�e�v�,f�t�#�*�gx�^;rt��[��@�r�E�b��۞骜�*ͧ�1T�~��[,U�F���>�+�vz�Fk8jQt�}?��pn��@i�b��й�|�$|B:Y�������"nFV���9��j��u��ݿaC{u�'��X%�E��w�.�&�T��Kt���:Ck��,�$ȹ߿�icB?|�ث����iY�0��V\W-�E�\���/NH���ǫ̕xp�v�@^g߫��T �Z^�惼�v���
�eŎ'��lCy̋�� ���k_@�Ɖ�D�.7h�c����.�y��"_<��2`����s*7_�>��`�a�P�-�9���	��(M
�n=O����6�~ªs<"Z�ܨ�L�P�)́����6��d���TP�Jk�aЦ,9k��.�B���g�'P�l����	n��~�/b��ǹH�Y�̀k���z~�d��*X���j�OצSi�5��aw� tzSƂ�H���{G��gB�zE�7�Pj��Й|l�%4�HgP������f'dU�����ק'��M(��2?~�"��}@(u?$|&���IÂ���k�`�iR���vG<1����S�Ƽ�ջF������߻��Qrk��,�d�ͷ1	�P�b@ ��Y�܌m�8v,��IH�nˀr&�����̓�L��q�#��mm;���U&� �&�&Y:�:N6��M�b��Z��d��4D����<(]��(��M�O�o����-����("�Z �F�	�(K"��:�[*q���Bx�\��X���!f��)g0�|}~�����u��֠�J�2-��O?񇽡��h>}��Ix�T�a�Ƚ�%eƛJ\n	�|Շ���GXv�Q�G��X�
��I3�:����̮�����en
� T�zz����/�6ݾ�
�(ra�dGL���]*:>4xz)Y�N��y`p��r[��}�]��~J�OiH�T�pRb�`p�!|K<�)h��Xz2x/E7��X۔Hg�l���M��;<���?7< ¤�;J.9	#�Hh��(\�����id&|�k�?\�K_>_��/�U�;��Q�}��5H�ڰ{�C?�mӐk�N��{TCX��J�"�kF��{�U��Zgo����G���`���[���C.�p�a�Y�pv�;������,���F�2�r��!>x�3����L���"�1l���2�j�]*�7� \^�0�F��NM�-)�j%(_� 	�8'��}��-{KՀ�2�H�"Pʨ�f��c6�+��މ
]���%x��B�?����-���Ϡ(���`h�����)rju�xc����@v�u(߹�E}u�{�Y�5��T�(���|���s�vB���x9���90֏u���0�2K��R5����q�%+�����3�⏔v)pR�$����g5��cƀ�lC6���HϺ���� �`��a�*H�g�$q9�v譺���Կ
5o��i.�����"yȯD~HD�����z�t�u���/daǨ-�NL�	v�͝ŝ?6�'��e����g�XNkv����jտ�eC �,6�]XE�!U�Lp,��wI9�Y�<���^n.����4/f`�b�D��I�?+�[K�VL��ɿp�:���{�#轠W������Ϛ^S$Ay�1��h�#>:��W�J���Uq�T#�%�pW�e@��CV��7oY���i|��g��D��b�ɏc1�̳��US�W\g�2�]�z��-F���3�+p ��L����R��	I�A;����5�
��Fc����,�{����C�Ӆ��xQT�ai�Qv{p"�P�g8�;��U[��ݤ�!ehk:�?�%�"�M�?����?����jJ��?k���z.P���Kę�c04��&�=3`�~Qז5�[͍�˔���͝�۞�@��:�T������f=N�n���k��s�2�~7�Ӄ#H{�* ,ɂ����M��R�T���ģ%�0��ˬ$Y���@Z"5n����_���%��� ��p�2��>{���6ͧj�WG	=I|m'ZI1[ܦ�OJ}��̮	i�_���1����a��g2��A�=�{R������#�����8I7L&J!�.s�k�N�g��<��}ǻj�H��Ҿ]���\��Y?!g�M�0A1��jp���}d�ܔru
�E���_��3y��:�r��h6���St�o��H�+��jVG��K$�t>ɩ	�G��6��	Җ�5q��������(��n�!D楼E���7�����+�~�>�ʎ�ͻ������=k�u�h����b���<oSn/��p]�U�Ν/��FR\p]�[~Iz��阋�ҕR��A63�/�D��1��)�d-���1�����GLJ��R2��y^���Ǡ2*�Z��P����D���up!�����j2�,[��p�`TÄ���r�=4t�����J�7��oF�A���p;(�����P��Z�R�;�$.B�km��%��E�HU�)f�g�$�V��D0���ZՉO�_X�ޥ�hEP�F��D1�g�(�yͷ1��oǮ�Ώ7�T{a�:�N;st���k� VODX#���nG�_z�x+oC��0P\6-��IM[1����һ�\tf�|R�ǥ[�ȃɵ*�,�5���*qF�q��Aw���`ܸ���6�Ro�H��������L6����?��g�SB�g�-��};{���i���1�0�����/����`��sp�Ed�V���e�3�]�k@�r�G�Y[�����A�=r�-cۛ���uز;�x'�/�_�k�U��j/�������	�t���1A��'�kem��Ix��@��n�敺.�M1��u���d�d�n�q��*��p����p7�ŭ�>U��_��y�ɲeOf�SH�FI��Ĕ���86J �����1I�T��Ӄ��Iy ��|�7�n�5����Q�py�-��$~���tQ�n��.��{X��/ 	�B��P���D{SF�Ҵ�xVBGv^`�3C!\���q�^)�Й���<���\/�xwêz!o����t c~+�Dc��iJ3�ػ5��#�x��7Y�������3&�l������,�����X=C���k�r�Ļs���z��`P @�&��ԑ���1������]#S!ϲ���/�2``G0��գQ�3徛��E��ml���C�y,N�1�q?�`��[2�L�:�#C��``:z3��Zܡ� |t�M:�F���%<z|�Ekx��91H+Z�s��s���G7��uJ7@ab@��1Yfd��r�/�q��E��{:hˡ��y��S������4'���Dtc���Z�$~w%[�	��0�*4Z���^�_'�jm 8�-B�Xm��E�'Sf���ۭ�� .O���5�b��"�N�F�I[��������	��B�q�{��_����g��m��dXϮ�8����l��d�̻uSk-��u�yN��7!xBt����|/������'+~��bܢ����m>�Z����x��B�?�@�k.p�{>}ZI��B��B�"�g%7=,<�'�4U:�?�6r+���P+?��Mw�H�����H��Ӧ���*�Φ�L��IM3V_ C��b�S���N&/\�pc�T_A6)Y�A�6���.ck!c�"|��}��j������O?�����%��M����eF��aQm}�h��6`$���N�T���\�G�]�	6�y�l�/~��]x�^�(�:��?V��ω�0���R�R�)_L���98?x�R�s�[�N6��dȯ^�Xփv���Wf�Mc��Rt�h���/�EնTz��+2�p�.�%�K�2O+z�%V���	#T����5[Ωc# {#
֡��� Te��@��Z��I�\K8 z6#:'۴3���'/8*�q�P��Q�uk�(��+�E�<�6ȫ;B8����i P�iRb+��
����n��g J�C�Q�AM׷���=�I�LYQ2�UI7h���
�u-���C|?��ܬk�9�p��#��K�!J�|w�,iI3��+�/D�q�*��܍��_=:�s%�S;�AO�4�b�#�W��_�/`���v��}���5ZSMJ��Ϗ��p,����My�P�/�:���KZ�5~���AA������!wA���Q����:Ow�[0�����*�|��Z/��+�b{xǧs�O�p�sV����a�����jq�$J�[k�-��RX+�n��=j���YEZ��������.��֮�B6R��_��|�:��sђaB lg|آ�fjE��h��s�/|˸v��y@���\�0���Bf�.H�������;�p=Ld���^�%�v���
���&�,$�tB<	J_@1�+�>:*#hh��陘ۃ��B���%a^��x����#k�6��.L��k�M�����B!L� ��+�|���Pn/{Ŀ0A@W0k�݋��F*�}*�1jEN�ϰ' h����Ś�)�\2r�d��)YC���S��[�FD_��_(��NT�n�d�F���T��o �RA�U|����Ol�AA���|�o�.�Sim f�K<���E�ÿ���jT��
՛Iݑd�u�	W ��si�����C���ќ��^z�3`�ﱿ~�a��8�Z�G�E�G��FI�t���t��H���N}��|��ә�aP�|Q�m�)�`��r=����:4������Dm/�z
1�mj��F���k���h�=�E%^��tD�r�	H\��D�ݑ��������^7u(�O�O���#�el�y��Ή�u���)���=Rv�} �J�ꮉ��K*�Ȃ)���Ā�ZF���I�B������ʶ��[��L� #U���F�	^�]풛cؿ�h�Ё���Ѓ����̐(xr�F�s�BA�p,�`M�V��TG!�$��Ŗ-�d���'SV��`S� ��ң���~���b��&�+�"kN�y+���Hk$>�IN���Y��Ffkʅ���{v��1��`��,sG�F��O�:)�6R���:�Gp͍��	fj���U�e���%�by��R���X@�!��W(\yZ%��(F^��(Ǘ\}9�=�ޜ7�_e'yn�҂*�eF�ؓ����վ�E��1MZo�՛Hc��_*;�xR!��bm�N�/?�����R>	6N���yy�#m�T�<� ̒�����9�+k��yeG��+Ts�H��I�\Ц��B�N�6�����z������cĺX�t����1�E�G^W�ED/n55c�q��@�؃<�^�'S������/p��9v� ��b�O4���Fl6ay���i|EM̪��X�wT���,�#�����:�3��<�`�1���M�%�j��#�nX_>�hS�.��:���\'u��|�{�R.����w{�����<}�pR1䀇�mV���2����\o��K�&�!�33a\�njY�DWG�m����.���~j��~�6���m^M��dٝ!��(e�8���@���Z/�Z��Zy��ĵB�loLKC��� �n=E��tQe�`�C�6�ۈp �v�(� 4�%�q�����Z;�HF�7<�+�߶f��/j�Ɗ�����7|w� �׀�,����P�@�3y�k�,�w�eF����Ȃ׶ V���@�(K@���w�mY�9'�����_:C2�u[	��2�`�-R�G�tK��H��[��$wT�h��y����=�뷷6]%1���f�Vk.��S��L�/�/����̵ٓ���
�R�	�1�G��u����b�����%���ʃ�o���S�:��Ǹ�ku�q�.veW�w�(.+e���xؽzq��lY���H���s���&�.M@~פ۪	Dq�æX ��mBR����F)_D��l��@�7
ң�ӗ@8{S�Ѧ@`�>�*�pjk8�L��i���Y�� _��0όju��!��d�27�\���r��uq��r6�iG�1�'.�%�j]��.�h:X"�Y�Ur�P��r�^�醍�P��IcX�Z����N�O��7+�f�7�<:D�i&���5����*��{�� nh���]�̶379W�_7N�f�a�I9�1l�1i��a�d�VfG�Y�q��0r��y���l�� U�̙���M#H6d	�۸�w��x��������>�K WUE' d/{���d��;�R�|�U�}��2�2���n��
�E���A	u�2��,9�e��,��x��z��4kjb�;������s>�h�YUό��p	�ж��y�)l�y�8ͪǆ���`�!��xwM�x��Wj/?�:�$O������Zv;F�%}�N8��Q�r���{��> 7���`��5��q{.��b%9Z���sԠ�#��JퟏB]^^p~�Z8�&k�f�e�G�C0����v��A:E״�~��է�8�?-��!����DWr��r}�4K�4��{�R �cW�/0�i�*g�F^t���9�Z )]�@:ύ�wm //UT�N�r�����~	s���{��������_���u#�(͕��w��������e�E��i:M�����w!y�髛��4��j�)�^̲l��.������]65x�:M��/6BuaBɵcyo�#X�Bb�� ��.}�q�|��<��RC�c�1�M�����眻֨,�A�Gx���j�������.̧U���\	�6e�< ���L��NW ���7kd���i�*$]R\@T�W)�h������%E�,������s��2W>�\�p��ΉT�^�$P�d�DVY΁J��-�[��v��`�Q8�
�WdRP�� paKZ&��rM�?��~���Z�,P�������^�k�N�����F ^'�B eio)>/�佦�}�մ�!WH�+�ܱ��up(<�2���[V��<<�&RI�qW�����J���1I��Y���WJ�j?ծ���1����d����}wޱ/U�(��`�
ḽ8A���Y�����rHo^bၯ��s.~�x��֫�Wn���U:�:���*݌8�y|FHl�X��5�LsDNb*���aN�i��h�-�~
�݆�Flq@8ʗTF�!�?8'��S�2OdA��<��+���M��Ēٶgq�����$���h�Q�PF(;_���l��aE��	�|�����бV�X��b�b��o� ���G�]�?�I��t��wIxfIu������w>������`{�r�]h��cd����"���N�?�2�7�ŝ\~��F2��?�k_�s[lW��ЫU����Nh#���yv	W�[��ڟU�y�����;K ������ɝw[0�Z��aݶ�9�U������Z�y~��$U�7��@�N�d�qX�d�gtL��@�e_�ft�	CO�!M��y��?lva����fU��C��^{�&ԦmA�_\�Z]�)/D�N(i��i����r��aL�!�3>I'*-��E��q.Z(&�W��v��6Ka�'���F�T\����`)�<?�O�[�Pf׭��Hr����n%y���	ҪYR�Mֻ�,!m�����r�욒@;�h�E��^��n����Bo<=��p�c��lR�1�Jjf�8��İ��iR{-�����iL�x��0��8s�g��B�1U�~�O[�6��@,�|F*��ׂ\��fCWo?rs%���(2a�G��E�4)�>�i�UB�� ����n�,]�s{6 �hO�j`�Tp�=����I�#R��Z���LT���9��*�y��(�Ȃ���嗏�4F.�ӻӲ� AE�	��*:�
�P�GH|{�)�k�M׆����L�|�%:̫�%�DO�^Fi�ڈ��&S�'�W�H� �i�?�-��,����%�7���+t���)?g���F=\�[豅9�o�aU����ako�nҚ��j�}��W5pr�ޖ�%�:�~�d��<�{�\V����O1��T k%�$ߧW�8����2�X�� �����ɪq���=P�|�?��b	��?_-�h��XJ.T(o��ͩ	�ƃw'A���[����/�<�{�3���kaq ����H�-�5=�P���ﻰ�4"�8����Y�ł���+��m
��]�Ϣ1���M�@�]�Y#�5m�)Q�F\��R�AX�&zvބ��9��m;-P z�ZPF���IXF֎�+�-M]*ඊH��v
����_�^��y�g*@s���w�y�07��[
�`J&Y�ef&đo�w$;� Q��(w2���2���ŧ ť��X}��b�)S����U��r����|+��P�$^�a���1g1�F�Y�0~�ͥFv��	ᵋH�SV��N�O\����,V{^�ﴄ&�)v���I!�t��+	~��=����󏓚��a����)	|��4���C#0Uc�r_�wU*�իKХ�<28
9A���ZQ�

�Y���W�q�A�L� ���f>�S�����3�m)� ,Q�l���¶�4���}�U�8��R硛�����Ҳ�-�+�+~j��h���!���,i�}�g���ݘ#:��-ɟ�k�,��~��t8o	xycY�^�e7���s8I)=h��m��ɱWe����P�a!�CG�z�@����̦����el�Q˸��p��犿vO�ť-�$/�������N䨐��=�Ƭ���e.�W��m�3���;�`	�z�)~/��{lem��w�A�䧦-)� �̈�o�sD\B��Fl�̓�x.��NH��F�� e=��+z>�ٌH�!-d�2��7��H�.���"Iutp�WHFسW���=�Sx�6���]*��[c�Q�vV���n+�9I����]�E�Hkm��l<`���O�4����3
��`(]�b�/�;��->A�7��bOǜ��e�5�}��Aw��X(��%+��4��8��M�T�!�%]�����V��p�r�w�5�Ɉ�{R��k�'�����"�-k�� a<�����d���e�q|��y�-D��]��}��S�Ya�~E���:N�]7�b���w
w�ǀp�!2�*�I$���_�挆��?Ed`�Gh�;g��t��f�$�����ɓ�3�O4R�������B?��։"B��z����[�abX^S���.�=2Se��K�h�|��bYz]uEnG��f��Ԋ���W�2��P�4�|4�6	���G��D�`FR�ց��kI��AF�F��>�_�t�9�2��8�ԑ���0�>o-� @E^�"�Vb}T���U���և��#5n���oT�L��)G��k=E!��٫�;�4`�y���!�� V�Q\���N�����7����O�����?�F�8��\`���G��vu�p��y�n�K�w;[@��� ����Ql���i����zuag`�cC�9�����#ʲ��Ҥu���, �a��k����j��ɬ���u�8����'F?�ﻶ��dN�M���9 �-@��Zy�y���̠N�B�Z}#�I
�!l�1/�a��� �}���5��b�!c��Z���)�Ay��)�PlDn��U{�2'tG.�p�mz���ix,!��`�W��XxW��Y
�t,��jbh�V��1@8�v���O�j����dy�h��4ZB�z}�k�X��I�y�Z���5��V0;\�+�[�d��	��6:7t3����1D�|g4I�o��AO�2P��b�A {�7nre#w���K��_
ջ(ً9��Fod�G$j�W-�y�t��P�2���"��˪N7�>#H������WԞf�X�P⥦C��Śu�;�#���I�LP��sτ��a�1 �����*-+�E�xnDC]�U6V�]�N9p���h��e�:|�h=#�qٹ�V+�J����ڏD������$U�h,k,'|��&��G_Ǒ�$���d�E<��t��<�oE_NWp�ug���D�=�A���ᩞ�i���K���b<w�[��|Su�sHE�9�K�1�暈�Z�ߗպn8��Wd�"fRiQiF���U8�R�SʕNR���~�������b}��6oop����]Q��y�[�G�*=�1B�Ŭ:���Ѿ�%��`&�)t�),�s����=��,y5�f'���������s��\�J���NV{j����o<@g�fVԃڋL�s�R���^�^�j@���7V��0�qa�>;^W˛ǋI����W�f�=��#��Jܪn�s�����A�6���T�p�~��}��.�������ymU��я�uă�j#!��sAP|O�&[����L�O�I���Cf�iɘ��ǅ�9�R@E�veJp���g)R�9�UQ,R�G<�=�n8�
��Z�.�i>�q�ۖ�"iX��ü�j;47t6b 0y�'�6�"1���8y e�Y�<C3���(D@��[�^����Û�PA��>�k&��j�3f(�E�-4O�ڰ��dF�S��E��}��u�H��.��8Mzj,>�z��Ϛe�;*�*^��{���.c�]���	f u�b�H�
��������.��Ê�|�*eJ�x�}Im�L�+��-�.nyW��p��*��_�q-��o��%�����g�;\�1]�<�bW�y�x��|�}���a��C��������=�~x���5����;�Bo���2[JZPdM�!������H�0�w��_�Mb1�����.�g�g$�}�/����$=����v,�K���P���Z!��q��L�h�ȋ�g5�ʝ�� �d�+��q�J%嘑��/s:}T\� ����[��0��`O|6V�����8i�~��!;�6׭��x�%�qϳ������3�#�s���������O��|dОG��>�:�8k�l��5XFE&��X���E+��X!ۂ,�UĖW�R��@Gy#���ދM�@hha$k�<\��n}���k���ƴ�!.|�/X���[2�I_X��� cp��I'f��e)����*()��9+�����߷��z���8��r��$.e->����f}a�~jB0Q0����9���Q��!�ͼ�E�m�+A�Xڔ��Q���b��B�AJ �o�Q�B�I%?�����[���V��f #�R�݈\� �p=v�F�P����yp夀�&["Sĝ�5/�"�'��K�.�b�o���]��`��-���?T����*J�g������HrT柭J�a�'��z�'��:^m���+�L���ׅo�y	xr��&J5�K��n�b%�L����2��u#(vRp�VϪ������D���w���W(�W� ��P�\��2�L���g��Irp�ڛ��C
2�׮q�1�^D&��9D,��k�����;|�p�O���vb�,D��&1������ų�@˘l�,��wĺm��^�Bd q�h�m^b���}���(�#������xA�ȰfO�GI�E��.���qd�26~�վ�*���xh�O����#P��7��������e����`!�(��s%%�K �U�FLa�g��/�W�l��u�8@#my2�4a�EMd\~B��������#�N��s�6�M�\�2�-����`�Cq�j$p�v���͉<"j@}۹��v4� B^a�N1D�=�$/�ʙ�i����y� 6C�ILr=��JB������'�S���GL��xt�閅�}5�E\�Ø��8�|�	61�x�K!�zPv��|_�u��y��B�S���B0�8)����}�ʃ\��ɂ�>��4r��B�D4�!tUf����:֚f�<�N�dG�Q��HYT;⼟���"0���N���o���N3+�rx���{#i:ڧ}��o������7�=�3gsns���l�A.�����X>z� ���$D��e���G����X���3��6X=�'K�w��.�<�r���:�>��d��\i�QR���ň���o:܄�I�_�q+��i�`%���vH��;������H����1��r��ww����E�c3��=�F����5������*AF���eś�8`�BG�ߊE}��]m~[�Nf���D6��6�U�Cݙ�'�3��<�eQ�D��<�r���j�k��~�]a�m@�+D�j�T��>�ӱ����U��+N@���12*q�S��Ί��� ���b�=h���ށ�Հ�!����P������e- h�#��,p`���Fr���C�3W8�$�ٙ����l�xeA Ѳ��Ouw��ٸ���ܤ�`p5o
���7X��g������v�l���0_D�-;dJ��\�����Rp(��fd�W��ԁ�[��q�+�����h�{.��
k"%I��i\bU��M�sN°dH����}!�$�M �0��8[��L�z����<��aS!�
�7��H���^�8�aJJ���$<�;���C!���JN�ע:�=��̽�W@���9U�2�Z���<c*/�Z@�$ J�9f���'�bIO�#�|�**d	�Wg�NY>�R3H�j�o�	V�EN9�����|�7�gs6A��Mn�q
,	O�h� "o\�l��r.X<�����|t�� ��D�ȯ����5;�z�<D},
u�n��6 K�S+6i�),}�vEB��j��#�b�V*@�_]$�߁�_bY���M�~�P%;�d̵德D��ԐZ�}�0'���n�ƨ�A�\/�=�$��-�o}y�T84A�2d��ƈV0�����`!�'zh��w	�V-c�3�������E�H+�~�����~@��]��"(�"΋'��q	u��:�3<�ߊ�廇�bșOŞIx�D�" w'J�´�x�h��+��VG(�� Q��^�/K���(p(��ԕ�@,/ܓ
�b��VZ)��2;��Q{LC�9��qu�)���g�M�d�"�n��g���j���
���l�d���=B� �L����DS1�Qy�����m��U{̱@S ���#�8��5�g��ě��[�T�#�G�waϦ����i:���l���ܸq��Ĳ�0jS���p�z|���2�ꝱ��<�w|��( P��9̢�5�9<�-L���>�|iP�UKM:�&DO#�Ậ�Mč�A:��#5p#Ϥ/v$�Xk�G�g}�e���?I����tA�8��:�d�-{`!|��k�do����{�~j4~���ؗ���m#�@@Xx-����a�F�s��2�)\��::��q���o �f��yo�C���	>Q2:-#�n�������.C����#� <z
��%YŐ�,"����3�����hk.Uxg�SzV�?�A�6w�A�j������� �c#���������6��Q	�a^��!��c}C�M_���5J��rup�
���H��^��U�6�Lc��3N��Yr��/���)"f.�n\�.��&Gb��� ��n� �#zy�'v��3Z~lx,�lU���}i?˄���,�}�y�0k�1��?h忪�k9��d�w9
����ώ��Hϛ�=��	��w�P?S��,�xq�@e,Rŝ)
aL��V�~;	x՞n�A,0#}�x�؉~��O�O��q��n�*��CrB9�ט>��Ý��/��hiF��{��K���/^ѩ� �m�E�p��"#L ��eHR�Pc��%��U�E����]�h<�a��hn|���*6QL����.�W�	�J*���Ԁ�b1 2X�-:;���xbd,
}K���C^�\�P��p�Ә��x�7���;3wR�%墻n�:YJI���!���B��cs����|�8t7��fJe�����I	�J�<8��ɘo�N%@��G5�u7����C��
��}�!��%G~t':λ�L,��<��csu�`tߗ8��ZB6$Ł������c���1ٶ�,[4��)���PTv�d�2���"z�Pp�6��Z���+�s�vX�89�ג�J��5ލ���b���y��`��k�p@a}�;��tl�V�ȫ�.&�~@>p{�~+�4���L�[6�8�����	l�C��Ԯ�m�b6�@��5lCB%�,��>�㑑�&z)$1�~�}�>�P�,�S�ځv�<�&��ӄŨr�g�*j�p�r�J�[پN~��Ȝ�D��]
#��?`I��_�-�52�b�f
:�٨��d�n1��&��R�� g��o5)~���/ѩ�7`��t%�ACY�l�w��ν��H�ӑ2ܑc8H��	.Orky����@����|�!f�����&v��؁��$���)M�*A1ďb�A������Tl��i����$�{"����lM �����IP�[��L�/~�BB����h����եۘ�t��q��t��f$��\5��oI1!�f�F�S�ޏXD��M$q��C�L�?j3�z���0'���Tg��]4�9f$���.��u�>�����U�_HI�p���[��l��Z9�iM�x�!�wݽ��o8�~�~B�7���(-�9���(��~���xF�]C�A[�g�Q�ED'b���p�]�Y'�LM؁���	Qtd��O Cc@���\��\��oЮ�����z1��VN@���U�@�5���\%?���O�*S�GeJY��Zq �gm����T�����Yڰ��p储���RB�NY�#{�#·KVM�s7Z�*L��F)�S�b�7�B6n�b��Ԅfp��#��g�6�&TV"�a\�Jb;�l�:\+v��=���)�}��j��L�N���1���%��|O�~��r�� l�LT6���8���M|����e�s&q�Uw7W_|=ld�,ʛW����i��2�ISz��O�A���D֮��J��h~�'Ak`�?�*��;�5#E�ŕ��%���$1�qw3���<`l�Z����V����x��LV��1�/yk�{��}N��1s���+�A��>�/l*�ܞ��� �譪]7����w����|��:#LV�f$��]nH�p��}�A[kZ�	'd�*C��WR�́H)q�����Kk����"�Y��d��pfP��E.�\���-��,�B��۳�G6/ Q��z\���.� ��`�q4#�*^%T�-O��w��TU���$;����d�be��>��	�H�-���=�w�P�g�ü��^�m��6����h�l����s<?v�vj��["�������H�;��ϲ���� W`OzYTd�A�����0-Bh��DM�'��tH)*�+\_�����6~�z�a������-�����'ך�j1�/`�Dv�~�_��S
g�*�gN�9Y��{�z���K�D�w�t��?ϫ�P�9�<��3+'r���Y��Jkڂ8DeD�����!Y���'h��slǥ@D�
^�x*%�}���"���av:2k�]��W�&D�L9�T�֪�?���/"c�;ڪ��Z��(�iSxq���DS�%�5
{L��=�"��z#Y4�F�=�ZN��<�O>kP���鳀�Ys���`s-�Opp��g��t�K�������7��S4VCb���5����PPH��:���wI�����o��*Β�?g\�&�uL��|�T�h��v�	���c�JIw~S{ڍ�M�CA���I�;e�t���/��2��(}6qM�Bb<���N]���&A��\�c��߱�6p�����wD
��f[0�W���mMdC�]l���'T��6Z�8�(��Ns
�-��b��i����k�4C������r��N�$P �ri��vH�QLp\u,�~S���Ih�J���_�
������� �6��H�����0����n����[C�|�v�#�klJg�-sw<r1���FٓT�A\+I���w$)�����O�T�0���h]M�������1MI'i�'��p1��a���mBM����C����&^
�E6{�����ѐa'0gP{6�p)f��������������*���E��)~w��J�=��Ҷ��	x�ؚ�o�T^"$a;+�[M����?��������m=~*-��ȟ�d�w���vx��H]��������ׅ@2�dP�?�C׿���F�b�����g����h}��ʰ��0�us�Bl�D�lX.�Vt��3o�w�"=�6B�QK~�fA�F�{lO�/+F0?�������&��a=H}�hp�p������!��1+k��A�p�b}��cs�����p}na�50jZx�U�Lu�n��A?���(�:=��	�T^��E،s��:c�!�_��ڔ7�8��)��|��wS`��Q��u��כE��)lY�,�앣�m;�E6�[�:���g�E �G,j�u��3Y��*I�]�K�>n�ӣI.h��̏Ϡ��P+y��"��A⥂LH@02{��pƸ zaܕ����T���@��&��I~���ɗ��ڐzmS�M�����V�����'U@�P�13�p�1�)t�ĕ�1�B��9G��,�;��<v���P�ci��z�ۛe�Z��/���!��m�������%��+�{��k�ȣ�J�v;�UGVo$�}��� ?�\&O/ũ���Eo��n�
::�v��?�{[R���.6h:�v�ݤʏ�Ӯ&HK���AJ���;ah��*%3k��?9^&0ZK h(,/|�j{�۳ق7����7j���V�l�)��L����-4���R������geЋ�$�ՠ�=_�33n4&+>���_?Ƣ_u��B�Ag��вRh�ϗ$�ߢ?F]w�c+�Q�ʣ���m��ǎb��=�H��8u�f�r��xuJ�I,_#��m���i���FC�G(bO��lD#�AGw`@W���ƹ�S��Ƴ#/�C��Q"�U�"ޟ|��E�b��
r` H���` 9���m�E�^�M:?/�X8w��S�w �6r���K��p���\�c��>!*�Q�_/>�!��΂��H�:�����(\/q���3|m�kv� ���,g���՚��L��b�"g�O��L��C��z�U2-6�$-k���p�W����{�3E0 ɟ������V<D��X4�Z)ԗ���dN ����c,�B��j���_���v@���괠�wƲk�v@��sxbwП�@�?yȅ��
�H�Z��k+;��H]JXP�`h����-�)����w���/��/�م���ף�(H�w(�a�)�Օ��9Iq�JD8؈`���Oa-�Fc�`���jT⽓�0��:�,��:�:��n�#{}#'y<�e�Q��m�h�!�G�V�PH���Ұ-��mS�D�=!�wc�M�o��CL}���5[�����Q��	� �V*��@�K@3�_`tJ�h�d�6��ܫ�4!��7�l4��o-g�%0}��haA���L{�~UT��8���H"^Jv��F���ZFq�91���)��K'b��q�۾-�QB��h����3�2�I�%j")#xD#@��rktڣ2�=��(�Ͷc!�@ ��-��b\��"�����F�#����ˣ�L��ܮ�EVO����S����\%�̷�[���L�ߜ��h���-�Z;T聪,}Y��+AH��ݧ�j��X���XzВȽO��Z�'����@r5�jH��qWE�O�j�!5�*���J���z�2����Q��|� 1�M>�����㱠|����>H��51c� �@�T^V���"�N���u؈�v~��y��rO�s(T/�/+&<RkO-z17�8f�1����^��ߵ�P/z�)�Z�dq�4G$�w��Q����H�&j\k	P"ׁ�a�p���C��O��&�K�:�CH�{K�hd0��Tr	ⴧC����Isʉ)��WD���D w��ug��,��/\ODF��۩P�G���Hoz8f���by�gZ�e:�!�Ծ���&�z����j!��?� �K�:���h+����d�����E;�2jBd��,5�ץ���]�P���ב٘�vN-�6^�A1iH���C��h�G!�7X~Ϩ[�Yq������2���.�ϕ2$��������8.J,��`y�j�tz�I�s귾|a��զ$��g��J�����k�urw�d6�ȎGh�wzW%�h� �f��.�ѹ�Tp;(
ߚ
�!��t"s�]|����P辇���n(������0��A�ǋ�*M�\q���@�^�!�q}��S7���|���x��p')�5,��|L�p���H��V\2��L���I�Ό��}��hxc�a���b��ne}=0}Fv�.`����b0�VRN�Eu�`̰�T6V�/�Ϙ���U�R�zT����]��7A�R�Dx����ꤣ������2��S���4�B��%�/��ƍ��{�H��{N�r��P�,��%�F�\�����N�ft�LI�rZ���!�εvF���?��s��nx�cJ�۸����T�g\�W㣫El�	��j^J~����W�z������h߮��߷ܣ�,fem���)O�=׉��4uQA���7d��l3a㛥򽽾K��,t1Z�"l������Xu#Խ��e֔c6�T�â�2Fq�-��Q�:lI�T`�ȭ^%vƠ#fD#D��Ae+�o�rR�/�	2��N�J��L~:�g���y{�a��fM�l��� ~�{�R��|֝5�>*��DNد��V�y��{���)�_�Y
pBi�X@�?R�8)s�^�2O�+(ݹ?�C��a %�L>���у��E��t��j�/�_ ?��m�h��ģ�ք��儎�Wn�)M-�~�7�g��:��*� b'-u�Zeti:"	�Kz��n��М����j�䂜��,4d�E��ֿK@�u���_���t?�A������ff�/��{s�1I��٨uY�2��g��Q��P �<A�������Ǿ{"� ��A�c	�&=,�Ǧ�L8ō���04Xag�M�P��F#�L�=��B�k�;�Is~1�����R<'
0����I[�R]'������n���0NmM��~,���u��g�Q�ЎI�2�	Aw�M��☛���><�i�1f�s���`���}ݶ��;A�sV�7�s�����o���K�����?"����0����b٧
x��l�
P��l��<��ӞB��&o���Q��鵷q��1 �y��aް�p�ŴhJfj����YT�]T}��cƐ��(~����Q�VT�g��f`�%j�^����NA��Zp9ȪW'��rD�:m��~�o�_ϰ'��AÊd%4��`a�U�hư����,��m���8'*X�m��y���~��)�9��-��)ۭ[>Us|��2�fid�ϑ�u�|��ݐ���ڽX�����	��@!]Vrdl`V��o���?�!���V� Fa����?t����C��`Z�p� �zlnffCO�'V0?I'�8���S�����b�z	%ODy	���JD��w+��ý��2-��pJ��UGA8q�.����h�:�K���IK��/E5��G���2$���0�n)�cxZV�=.���SE�F=�)㢐aO���T��$.�s��b���A�\JP��2Np$�^���pG,w���ǌD�,hۿ�����<�Z�_��\���bv*TH��z�XbK����b���Oߪ��[:�;Jc�9n!A�(�=���]L���3�\�Ֆx�ŸSQ1�����~��!G��mp��>�i7�8��C�hH$�����y5�Q��%�g�P)�3���3VA�<�G�?�i3r���+q����a���`uٴ�psg�ieұa��3+��~�ʕ~pO����N����h=����x��}��3�Ӧ�u��H��.-(�l<�Q�VK�M(V�Fc���jY!LwU��5&9�� �TTLv��n���N15�FX�T5�[$��V
� ����#���@��16�e��O�lA���1�2^�'��]�šÉh���$�lZ�5]_G2h+֗$�^��V@���l�U{<��ߕ����,�� �xEY� N2|.�~��G$f�.N���&���ܛ��ez]g/�1u�4���Oa�_ �7�v�@�`Y A���/��6�ى�D̈́��{�OFǆ�i��.����
'�
BpV��cQX�-��	�P����_��c��r�pG�*$R�9���RTUYS�|D�n.3b�y�2t��-��wN$S$��xƠ�j8i�� �钬�������P
Ü���,�}i�]�4����27Øۻ���̓È�4���4,&�(g�BŬ#�2E*L)� ��g
�>����ky��Jx���D��k�^v�x���Jl���뭚�f[Nx"^�`۾>`�H�x�FNĩ[󯕟�Ƣ�}�Yr2�z'�GJ�q��VJ�`V��F8��\��Ő��q߄EG�tM�1Y���1��j���)d�V1P��B��c�҆*#,�1��!�~�6�aN��r�G�ޫ�^Z�]��(�\�*;��������Ci ��_X,e���$�A�`����9�v۶T��J��ǿe�q1z?�Fy�V�!��7d�6��i�d�߹�.���k��bA��ejL�}k|�%�-D�$��9�&�;Gw�� �РƁ��j� ئ���-��g�C��B$}.6a��;t���:5a�"�96E�t#�^��Fl�8�탕l�֦P�X�N7��G���ם�!i������e$���CN$�="z�U��>�Ԇk���w�!:�<�x�nAb���=a�Mˁ��3P_�v�Eg%�ೀ[6�K��"/�6��p����c����������������<�x��,��60kzL �
)��J�=�i��_���=���Pv�'_�����<�4N�mǑ��1�=�7⁎�]Z���2�����~��V�e���l�t��h�-���:�F��fsο���?�j񞶘��'�h<�DyK��
�l�u�$G��S� ���b��B�*���.sWT7m[ʯ	CJ���D,AT�q-Ӡ�Z4�#Y�U+���ԖY�e���S���"kLe\)c��b븬�u�,n1�̟3�A�>l���	mK$�C}p�q�:W�b�$Е���t�u!}��x�*9p@q[L� �w��K��N"�٭ݼ����ǘ������-��yb�5f4w�6�!u��S�'*cE� Q߆Zl���"�L�J11���!�%K�	�f���W-�؞�L/�A�P�E$B�Nz�U�=�g�aeo��c`f�oD�uf*���"������?�)@��]�"��ya��>�Da�J����x��D�w�dt秾�Ȫ��th7�m�6��V��1�/�S]4� "��ʔ>�/�S�1�%aS���,��;�E�`VO>R�Ǯm��q�b�^�A��j�x�6�M�ʲ���n����5����靫�+b
3f[v��Ig<I�T�Ӓ��2e�4(\��t �g�y��� i�sۅ$�մ ^�)  �^Y��S:�Xܲ�Zz�o�_-W���*_��V'�@5 �P��vA���x��)�E�w�cCE��
x/����Ro:�N�JZ���=��e��p���3��x:=���v󚦷f�o�����4�5��94���5l����S�E�ژ`��[<yF0��-6P_�-�fA�C1q���-!��Į�� *8D���-��`F���������vx����C ��{@"�ת�,��pkzO
eK�L̲h]�6��*��;�Q�_�^y�;�s �rz_�V.Gw l�� ;�����}��|�h2̧Ӊ�{18/"y����^8�.S4|�K��8�8S����;N�L��*~�D�{}��c�po��c����u�j�\���[@X�>�󜿫I�H4�g]�T^����|n\����hC����;}H{���c2*9!��:���.�1����l��/~d�b��w��J�ˊG��_fe��mK�Z�r|Ğc�p�7E0��1��O*�S�e��.%��] ��:�`Oc���I�g)
�؅a�N�r��^�m��̾{��|�ߤ�n6�����j��������)��j;��+Ҽ�D�?/�hBܕQ��{%������>�Zwe�if�4��^�h�4+�w[��|��%�a"��z�	w�dч�40���<��a�'�R���KTqƆq��6�i�$��07B���6/�����ǐ�b��f��>w���Z�X�a����h1��,n�*��C��+�a�<k���.{��m�܇�,�[dڪ�������^׺�8�Z�d�M�*}���?Wn�<<��n0-�%�MRH��#�{��3G�Whr�f�} �~�{��ZP��fj�f�A@�$ �G��SX�:�`�8\CPXT�]����H��6VO�l�O�!��Q�B�w����H�ʐ��):�g��m��)J�?ӎI_+�0�@�*c9�#���X��í�vj�����^w�rgL����}^�P�Lsv�Q�t�ś��p�E�h�m�{��S�x�a��6���L�(����;�S_��j8Q|8sj�/��aׅ0/_=:
�_�#�(��<ϥ`�.�{��>��2�E�
3�am�@P��a��؇"�l�^m��Й_��e�UM3�0�&��h�%�}�1t��Fk��FU �'l�8�!��a<?6#�������}�+ʓ�J���Pc��`�C�&^�����q��ڲ^Z+' o-6̧�o!I���i���B/��m�H]��\� ����$ꜮV���Џ"^�Ԕ��@/�F�Kߖ~���:�*K��TU�J�� �'A�����0L<�B蜚���sM�0L��W!D���_���	ś	�U�`>�Ƿn�����>�ͼ-��sU��͔�e��Dd��Ic���Q�~����� 6�����O��������R�ıwa�+�He�v����������i����)�'�}=��[}�w���0O��l�P�����@�g�T�����sEw��!0V��e� �h��ХMQLF�����I�KNK�Z��]�%G�$�˙3�fB�bR&�0�N�n��+{T�E倩|��&�P	p�����C/�H���z(�u�K�rݧnp���ý �����+\/����B6�yU��8o���?P5���K	q���F�G�Q���B9�5�N�5���>2�h�y�әo	Es�E��搸L[��z(TTr40����s~X\���jJ�^�G���rl�[��q$i���> `@�	t!�7P�tD��RKN�N���
�跾��x�DeL�/���!�PR,.,a=$d)���Q�<B��	��1��\x�~o,��=Ħ�dg��[�:���gQ+�`S�Q��Ȟ�Ѿ�&�&+�/�k^T�H��y������e��/?
ny��h�6-���P9hF��J�8���3�}5��p{���F,0�G���+�K�s����3������Yܮ��V1�q�i-K!�"��R_�t��Qk򁂙g���y�l��J��Y�,�a��m�\sY�re}�����$�ZY���^��(��Thރ<<Fx��ݰh��uM.L��,
���N@8������v�μ�?߿1�9���+�Ds�?��:z�-�_pWG�~w��g�a�`�����*��<ރ��~:;�Q\j]�z�!���������O%�^5���M�+0���Oп��X02�(\��x��D!"a[[ʛ�����,���=��>4rE�����H��D��� �{�J�57{��q���g��ފ3�7�H�O;�q��w�)2ڀ�"�}gU���Ve�3%g�Y�����=p�2{E��WCV�+9G�2�G���t�T��6Lh�,�$���������iN�T�t3��69m��2ո�b�W D�Y����c�H�/xi��o�
�5-�D,J�E��� ��F�:Q����~EV�}���M`[`���U_y3�r�˵�7Ģ��t�}�4P��?ۮX�}ӇBU���"(�A�U���?����hｴ]����3wԳ�]���]�W5�������lK�햮ZI��u��
 N�y����g�6�l�e����v8[��>��"1޼�S+毁=O�@(�)��<ب1c �VB33eO{�]_k�AG��Xc������i&�)��d���/�F0�sC�8+�	������P������e��������g>����D�F�8m��ذ����v�]��^��)L��/IA���sKj��%�i
`<�p��*�G��X�z��MŪson�'w'v܃=�º����|F9dn��̳Pz�O%�F�J�����.`�}���e@�Q2�d��һXC�0�����y�33��]�!�f#ԣ��'�?���r	}����������U���?���נw�nF�hp�Po���������P.A,K���ݷ��2�o4	�-ሬ�~�9�7���5�����ƍ�ً�|�ؖ���xې�C����T��Y�#AD��8!�A*��6�Ց����
J�OK
S�F��
�g�������"��m}�c���h�`Z�Aot%��-¡4?� ��k��ܬ��Jk�=���~t�����vͮgϨZҔ-�z� �d�Ǘ��qXkW,�@�Y-OO�Fa(�MБ�mL#�,�L�p�ڄ�i�.�<�T,(e�7r3�W�_^���0��_�M�B��@~.}ط%�����*bҟ��Ҝ��J+�|��{�T2��WN�s�"����NGL
�n;� Xn��JW��{^uSjGS��ZJ=r2Rxvi��D:+��u�N{����R�pr� �>%'�d�xօ
*	�an���������%��ҡ}{<F�i,],I�Ѕ+	����FoH[�ν9�户t�3���8�J�*��R��RC��θ�d�ex/�'�V���p��+0��ǺtbychIJ�Ōo��q��t|?��0�xjö�8N���� i���H��P �{g{n���khLkG���
�&�s5�������{�&�l�l�/�U�Ѽ����`�~��<�$��p0�L\P痧X��~E�=�%6	�&��Ԛ��!�n�P?�����c�N���C2�zT� �O�,a#t�)a��$��g|��	�Cm�ڲ%M��z��$��H��=���?�v|jhI�쟝NIك �Ք�Lf+p��j��0��iJ	O=px�Yj	{F16>	H�l��F�y�Ǆ�����:¹���C��=3�R��H�<��鱥	��y�
"��s1�p�f}�aM����붉l�{�䮻��T���_@��"5�<QL����U[�v!nׇ�� u�W
jv5#��Z�{��?8m�K8��睁Sŋ����딇�c��C��|:��
eә�c�Cҝ�|6^��P�r]��)W�Gh���F+��)a�pp5|ȇFrl-��D�p�(F�9vs�a�@��%Ͷ�c�����w|�GV�U�Q�-eT�8�|��_K�Ic�͖�3M4\:#��ڛbWG�p��A��A��g?��nÝ1y�ǘ���\Z,�р��)��X'����p��$�?S��i�d��-Q��Ҏ3�f��%�&wu	ˏ� qlc�{�蟁�!|i���~H� ��jo�e&*ǘ���\�X�V�Q�,[���GEN���+hE/���^e�D�h<}4�\?��6��|�A����y[�s�lz0l���L���Y.xZ=Hut�܏5�3Ζ��9M˪hg��[^�������=hgy�)QLF�<�!���j�^�"8�����j��|S#�Qgo��U�w��?�T>�.��\b���g�ܹ�Y~�7� =3�Af�=��}[�6���A�w����.coL9k��	��\z��LpL���������3�ōj�5���V�Sh}��� �MQ�p&&�� �8�S�7�/��};�;���+�g�w"����NQ �m�KJ�v3��)�E���, T^��&��j2x'c�x��a�l���`��o:/�bU����ix4��~�� ��\ ��~,�8��qu�?j��h�RzǶ�*�b���zCA�/wf�Z0��zQ������祊]K(������&c�|euf:������~�:�j�-�|�P\$���ppƪ+-�y���":b�]���R����v�� 	��9��;�*�ε�j��=v���1w�KAXvW;��ߘ�r��^�{yH����$�)m�Qa�DA�;/��{ r�;'��Qn�n1���z9��l�m����t� J9��J�o�{��T'�WJ] �=W����Zo3!������jH�Q�	�N�� 2}�_����R^���Y�_7��f��-Bg�WB����e��<!�N<f��1)�M�u�x'�hd=�dcb7}�S�_^s���D��^��b=?������K���t,�
':Z���6|�tY������Jpyҗ=����}j�dR���bCA��2L�]5��}�@��j������|��$�%[���R����];�8�pqh����Qj�RW�V���d&����Quc�$�`	�q�v�
$�D�4^��z�s��9:���	�І
g�s�m|�y�<e?�ݲ0��o��,�.�Q��| 4�Z���iޘ#�,U1_h���4M>Kz�[Ķ�L::N8P�#+��$h�9���y��0C
��`�0����l��"�)bvg��i2/���ʀ�2��	d�&O�rkg?�ǆ�,\+��MC��=���w�gz�O�  5zK�(Ҷd�l*	���~)�H�ʋ+���G���z��
g���%�ak�/t�X`�!�0��7��W�e�T1���,���ߊ����O���������N0�:�`q�T�>�Jƭ0׵��h(��\���D�h�V8N�Xk�!�CQ�p�i2-
��D���N&�􄟈���Ĵ!��	G�D���e��+��#�u#@g��kzA�ȧr��a�2m! '�[�oؿ��	Ixv5��/�d����7?���0�~/���*V����ɲC݉��DE�����S����%�=YFV���I�N�`p<K�Y#�78��/��] �S�^BB[�/��ݞ�&�|�Y���d�O��_yᩥ���b;�bs��JpL�M �$�>�t�G��Ֆ3���G�hB��jy���������/� ?���n>l9�rѨ�3Щ�����u�w��R�J Y�Ќs��'�MP$��B��N�sz��75�'���I �V��Mż��n���C��P%����q��J�WR�9�N���_���B-��ڞ~|�:��9��>͉��!̴Z�@�/C$��^�" ׿�vŦ�D����Ο8��u��2��}��}�o6	/���=�Ӄ�nl
��9|ץJ�Z��ײ"dC�U<b��I�}�i�K�(�q�$)'+�S�YD�@ ?~I��?ϝ	��rm�#�V��w'�����e:2��>��l5'��yU:��zf��o����dI�pFQ�
��G�'cz��q�R5d�<�"���0�E]�/�w!0V
���4���$�Wg�(O��`>�@Cf^��K�ܬ��
=��y ��5�g��?'��PAto�5���Q�⢲,T�d�8&g�R��Ry0� ��ڥ�睜�όvF\���Gzԑ)!!
%��%���ܴjU���\��|K���������b�"P�PT��XF	��\K'���s[П����^�4��)�A���U�oOTS���S4|r��BH]X��
'�. ����6[B��`�lR-���)I���h��N2%�Mء����k8R��!�!�s���ެG�\�>�
}��9��j7fdi(����W�@���2�����s��-�l�}�k���xaje�V
����k��ٷ-�J�Ϭ橌1'��#����<��\��9�3�Bғ*�<�� ��CX�6:ZY�q<��	((�ڔ��j~������P�6'|>�U��͞��:��O���)3�ֵ&,�_bPr.�O>��>�G�o�O�&�P��}3��ܾ�+s,'���w5��=W>^U]�}�[���dÊt��X�P�SA�@��eS��lsOI�����@PҵX�d'po%C�=��Q)s�!�V��3��e�έhA��׮�.��B�y	�A֗��>�����n�D����d�B!?lG�M���Df@���h�q����G�v�����$ �o$��A�rmǅ2,2F�Zft,]�6�D�`*P���>l�m~�]xh�3k�ux�RA�K(*!M�q���d��쩁5tS����l��)w���3V���q/���T�t�a@�g����3�C��#i+�q_6�t%��a⠆�F�4������x����E1$9���>0ZQ߰�����?WcԦ����x�;�9{dC�G�SX��j8<�wV�Ց`;,�E�
Rp�c������P	�q�u#�\,X/uQ��m_A� k��v��5�gŖ�å�ӵ%���78j3��/Oj���1�L����S����I�D����_��/)#זs�~�r+D�e<�e~_p�@G{�F��H�B��KT��w���4d<z1yd�]��y��^&���:"@����k���gF�-!�R��ʕm�>t����DK�|�_����.��g�-ۯ�`b�+��������G����Y�D�|�&��;��q>,��|��	����||O��x_�!=%-���%	G@|U�z�sX&�<�쮭m.(5��K��`�:�Y������\�� s�>��٫_�U��f�c:(c����b�	֣UÑ�%����W�/Ù�a*��Xv+oQ�#/Z-lU«[d>;��qO@,l09_J"�
����1Y0.�6T^C
������S��ʾ�X��<���%��Cr<��닶'"PüZ;���9���bR#q֑2!�#��|�B�\��Kn�Aq���1'?&%�U�8)��}p���-��}�}_�3�{l�@寘f��>���N}���iNC�N�-Nr�BƧ��*٧S��B�N��n�pI�yԮ�-C�z��ZR���ܹ�	>���S�����$tDՎ��dV��������4�w���0�djP��z�⼮��r���:x��_6�$=+�}E:����y��	�(G�����e��Aڜ��"h:�T�K<-�M9I���N�PV1���CS��3Pim�W� HDc�
��q��w��w�VV��g�<ٸMQ �܋�c�l=aP٠+MRMz�	`-������I�n�_��'�jiZL9xqVd)X�0e_�ϸ!���i!�sy�1e���zcӦ�����Uhu�[�_�H������35�F����`�m�v6si��$>:�@ݚt����۫�]h����2�f��	����rN�؆k��?lb��!�P��M�%�l `�Fs�g��l�a�EN`�X�o,�'�$s\�f�Cuw����*��xWPC㌦�%�-���>�*�a��Ϧ��Y4����J�f^mlt��P�$��pߘ���S���$����3�q�u���;�����^�~ɕ��x䰖�l�ӹ�w4!�ћZ�h� s���� y��_"���l+�N�ga���n��c�u�FBs�n�g-��~���5eq��9�(y�̀�����ˏ��ܣF��[�^���q�i5$��cj�_�ʿ
e����Q$ku�uŅ=���F�z1_"6|S8� �ㅯ�8_���ˁ�x�ʯ)+��|�Z�}�*켹A.���?�80AmF��ߌ�]?{M�*:
�������B.Z͌��R�'x^���W��� 3� �7h�n�~�֓Pw�xI�}���E_� -/�~[wvrş�	 s�˘PF��j���JH-p�R@&���$x�{�E���lap62�i\�������Eyg��Y��;KZ�a.D{X����3�)�	�F��Z�	':cñ{ ���������8B����%�}+�&W����1��J��tE�"L<T�>d�Ky�$a��A�v���!$ɵ'9;v@�rB�x5�8>��3�N�/kx�S�*-w!?��Xm�]�5,򻃼�����ɇ�VI�c�^�*����_M'�<�Q���7֗��;#n)VW%x�BH0oq3�i	�ȵf�O�o�[�ʢ�b�Ows{���u����wd����"���l�r�&�87~!��]X��;����BI��t��󢕣��DPs	J+�Q����#�쓼MS�K�rH���z.WKA'<�9���٪s�@�����[�Ʒ1��+�Wu�6��G�S�·8�m	�2�Z����MbX�S<�8`MgH+��%��3����E!���6O�'d���Z4�XkD��˖z5�=��o㩩�HLe��Ӝ����ꑧ�|L��<C���A3#���0�Q�����BJHJ`����X�h�IɈB}��v8��S�l�/�0�֬���:й�3�����	�t�R�H6���ڿ־���?�ڙ�����Ո��,/^BA�V9��ڈqTo;ڬ^����t�A��^}:��WzT���ѩ������;$�(cKE,�D�o��н��lž4�̅�� 7���i���n�w6@Px�9ԡD�����lK� ������+Sx��g_6��#�W�=��s�|�Л�����^.B\;�ޒR^�F3�YH��=�9[��Ƒ챰���k<�TהL�I Z�:Smc�y���,�ly�W�2o�-PjɅ��\�l��E��bdA�Խ��T=g!;��ֿ����`K�{��VoI����Td"o�l��YL3��[Sfus���"#��*����x gY����"1����Z�ˍ������c㻘�(!~ܦ��W�G�ѓ j�c��=Bip�M�~(;�iS`k�1���{z.��ڗ�ќu0���a�[���ܬ�!�{U�iPoلX����^I%�I��s� PW�o��n
�`,>���~��;��"����3��#K��P�L�ln���;��'$N�_'b�����\����k# 8"��gB�@�)�E���XY�όxO��Ǖ�T&��ϽL+9�Ǧ gj��&��ӻU��r}Y��f �s�R"���:�wx�`��A�l�7_{�ۂ#EunzꚲQ=��j�q7�hVy}a�������D��l+X4t<�U��xW"/N���_~$��D�|�?zu��d�OՅ�p�A�z#��Z^�5h�#f�pT">�`4W���I�O��}��P�iU�O�~)�X�"��Jߥ��)Y����؊R4�K�5����\l�+���3�"�z;Q&bzl���9vn"V[�0�.�2�v�RvG�[zuK�͍�x^�{��'�G�q�s&g{�
P5ق�y������/4d��Tr&��g�w�!z���7_&"<��7��� ���H�o*�Ue�HP��W�k��Y��U�{�%��,[a��j	���n� \./�<���������a��_fLx[�c��?���U�#�/nv�6���C"?8{U�����ԧ��ZX)�ʞ��a����~^����:��O����Q���:NS���f�س�m���v������=f����3ԁ�o�z���~Ґ0����~h�Dz�`@_�'|��$>QA�����72M�!�+��B�S�C�4)�f�N��G�h�uY����L��aK�;�2�*��+�Q:1}��Q����R�!�����"��B?"9@w	�?�$�a��E����@{�:��V�kh( j29Fe���ُ����(��^N�!q�Z�����t����Я���`�픬��TU��h]^m���`>$j:Mkj��%v)K�K-�	@^k�'s�T�}򆀯�e�9C�D1��/�db�r�0I�j�."j#<��R ���H6�I�qĄZYlc�fT�(��/9M��F��vJS@�
e�'�>)�s�Q�uۚL����dU�y��H$uCˀx,E����-	H��-+R��|���
 �9�r���%o��bJ+A#�S\{�o1��K�O���<;�p��̒ج�f�k]��� +�P�g);}6(��׮v�����o�

G�.䙳�G��S}\g.�"푠���m ��	�!.l5L�\���_�m̫L[o������<��6V���ʆ��7=)�x���]�����U4�ށ���sZ[����m/l���c��T���O��z�J����ſ���x���F|�_��؟����΋v�e�\ʜɃp��LD_;h�����{�Muz���dv�o]���������S{��1��9���e���ڽ5	b�T�󹜊ǵU�g��8����IH��������l�"̹f71��!O�*zo�|��$����RE����sP��a��-
B�5��WkN��犔�(��U<H9Nkz�k�:�f5���g�߁E'�256���T�WQ�LǗ�Rs�9)����t��*%k=��|�<��1�5g�nt��r�MbA �ͥ)\���$�6�X��EY�=r�����T��9_ܙ�G��B�PSQz�Ȼ�}�Ǵ���>B�������W@�UP�~v��4���� 7)(�-��xa���&[�^��U��Q��T�0�������1.�c��������d�RRT�,�3q�MZ�Sđ��IPk�����HC�l��>@A��gO�U;�t78N�(ڌ{�>i�2lV��`L�q�Tw� ��晑���HS�Ҭ�Kf:KcD�P8�m�6S�x�8�k&��yj6Q�����^w(Ô&����拚_&�"�;�֙Y�e�eSE�����������}��R΂a��WBݓ}*J������P��֒�^�2E����=P�qPA]��W/�Ϻ߉\�:�\p����4\k�+��஁��y�?;SZ&S��.d8�������p� �}>D�FD�6cJ��u�D�Pp�j��Ǎ��=��s|k�ߎMi��A��;Έ5M��O<_�h�ڢo
�*�����#�Xw�Z��d��'/Ȫ���CA���3�A_�͸1-6�����J���A�f�ί�)���0�/\;_U�+������P��?��ǜ�P��C���̤�c}�$������c��q�2 �\g�D�9 ���o]�qɱ�T �׃�x�y��s1���p:��� nq���[����J�.�;�~�����p,b�s�l�}�"�p�:�f�����pșj���K()ҽ>�Ai^9$j��8�X.�l�37��G$n�M�s�⊰m���"<&�e+"b�EQOc���?�x\8�sv�dH�Ͽw��u��=������s1��}��d�N�׫�xA���S��wj4��J��8���K�ʹ?44�7sH˪��bȔ2�^�B��:G��T̀)�H�Ȯ7,�J�"xq�]�}�n7Q+\��v 5�lY5��������Ri�Og��|�!Z�G�t�0���c�l	sX�� w���˗^.�Q[~���AM9o��,�c�(���t��鷷gG��z���W����9H�S�����ϕ4O����_u�X2̽L����09��t����1�*6j�+�T���]\nx[F�ߍx�7H��F��n�<��x�`J����|4,�B�Yr��X���)uFٙz�m*op fXCm�)N� �6�՝�"N��do��zEP0�XM�p׋�W�+06/�3
���Ԣu@��ڦRl#����/����G�A���e���*Ò�5�F���u��J��){T�0�g���`�#���6l����ud�#���>-��!��UU���f�����"�-���G�Q��z�����L�s0e�� 73扠z���0�/���qK�j��X��:�,�v�D>�5[!FM@�Ne!>(�9��#)���M$�I����R������3M�)6x�G�E�wEqh`�V֤�)�t	/���{sG�PM������s��(�p]HMNL�<�O����2,�����@�[@�DAy�f��'e��K�Y/��=:K�(nP�ו5�<��`9�>;�7��a�(Cu*��_L&O���69��t
}T�X��I?`a7D���>A��fv�**NM�w�ސ5;��]�����5vl�t���m!L��䝊;s�Q��p՝ޜ&$�T�V�Ltw3���;�����X��B���XUO:����$p%7����Ay9�2G�\9�7�"*�XA��G���z�M�K��~�%)\���d 5�.�Xk~n��_*�&��<R�d�w��j`�w6ؕ��v�@�a�"������(�*Q��FU]�N�f]�xJN�R��h�� -��V�$m�փ����Sh�k��ڧ �Oa�����ȝx�":m�j�@\��&G
Y8�߿�Pp貘~���N��$B�;�ϮPN2�����Y+?\=&8�z���CԜ�Ǚ� W�NIŨ�ᇨ�77-P���W��[l7��/��ʼfap9�ul��$�@)�!�����?�hI�#cba���gR������ǻ�� �Ǧ	���d�/1Pgqٛ)���
��ɔ��nX����*����-lel[8��h��1��E�d8�$�$�M�SS�����`⡳������ğ�ti_���!R����_`M�� ��e���F`(2�6����cbgz*�6�d2cA��v�_��!�:
�\�^�������mI���g�.�nc�9����	lq�&z� TC�1���?%R�tT&͕)�����,ˇ���7�U0����a�����]2�ҏ�o�e(�c��#���/6W� ]q���{�ߌHI��S$P�@d��}Xe��g�뜞���s[p ��8�۞v�r�L.�]I���\�n�gۓ�nU�Ƌ�*�J���q�|I�?�o��k�� ^�L� ȡ<O��0�|Gz6�t�f�������ڌܸ�vco$��rE�`���J9%u���c膺�֣�Q�枹p[��X�ه5������0
w�ۄ�J��Xуr��؇�X+�EP9�6��6����W�*�F:��~f��u�z���{�&�z�u(Wg�P�Q�×Ʀ���."Lϭ�����ndMmp<G)U��pw�GA�i�sM䬠\,<ϝZ�$�:A�:<�iV�ߖ��fa��T��
��G@2��q��������/ѕ��Ms����C����Z!�D8LR>�j���}8�nJ�L���Qy��F�Y颞�7���ƇE5�Е�<?���o`>ڢ�8��n��P�愱&��}JB,��f��ۻ9|��,~�����'�t?����{ �zN9�s8�c������y%��g��rL���q�3�q�n�7���vGI�Z�I�����q�C.��D�`�*�t�9�)T�j.�U�F����c����A͒�V�t�"G���C�ҏb���/�.\�-t �9ۥ��ˎ�XkuM>��O���Y�Ud�M&��-6.��2��N����
�)����~y���r������1\ �nt Ҭ�ʃ�E�}��[���d��}�OYh���g"ZU�� �"����?Tz�|�L���PB��aI�Zz!6	�1� ��Unt�q��f��v��Ǽ߄v��b=�~�Q�{㗲|�]Xj#B	�D����$)�rtѣb���IN��Z�ވpʀM������T���i�'����pI.�w�����!�w�#^I4ꞗ01��y<Zv� ��z�=D�\B���m��FT��-�N���1f�����$�i�C�rµ*�<����|�ch����{1AH
����4Ia&xH@o�.
�P�4�������[��{�ҽ�Wu�o�H�B��ӑ\�F���/�R<�4u��ҥ���3��T
�䟝�;��e��~��3�w�x������Yv
�O�g8,�/��`��q�����O\��.2Q�m4W�~s���4��X��̴k��P��X��Q�]ߨ�8�J}]<ಇ��V".�a�Y�SM�B�4��J|}�3`_�$��}M%l�c����^�Y�>4bN��U�jہeIP>A�5��mH"�H�~�d&3���؆k��#��ǥ>~��AW�~&A>�䏋�a�Fʌ��R��P�!|	y��<��i�F��̟�.�y��&��)�F��D��.&??琌��o����Ω�|#�h�����p�U_�^�T���ME�&/ F�h���C��hni��FH�F�w��_Q����cU(q{��{�c�� ��3Ո�~
*�W���42�=�V^� �r�7j�x�ׂ[��&�����]�<��T����3 ^�?5qq�b�����#a�L0���9�"��%P�:�E<�������ӝ�s|!6�ehm�=�Z3���y2~�^�]��W���O�`���eL����)�W�Mo}W���Rmɉ���9��=������b=qf���9�	;o䏻��)����@4֑ݴp�]��FS�gKI��NV^������p�$��o����>C�h������)��˘)�Hc�/oTP�c�N��2��"�G�X�ߠlgx�����@h�hE'5M��:W�k��0=���f�pV,��>W���I�>5���{�I��� ��-x-�}|���78�+��=��tD�@��P�.FMQR�7�e�7A�4�'F��z�%�Ν�x l�Da��u�:~�Z��{f���5�����=[α�/����
/��4�d.c9��ٰ+��p �Ȉ J��5.�ǒ�*�=F�ߩk�������k>a+�gC)3͇s��4�R�=�W�~�Z�1�����$r���]�C�����������X�˩Qe@�5�֋)�K��Mi�^�v E*~i�i�[U!�5�r�a����3(�!b��О���-�P�j�/���W�坒�@	F��2z?Ot<2�����R��v�*�Dn����J$
	��0�Wc���q�H�vv��Z��FD:���2�<���3�2l��Ȑ��)Rv��\�O�sU�o���PM7�ߐ�GF�-}�31K�ыؿl7�`bA�g����i���DR��c)��=@G��$m�O�x�b��7���D�zV�^�Wfܷ���[֯]Z%(���@�L�L�c��?�ʅ'%5�i�ENS��԰}�{��Xp`啙�kX� �=� �b������,p��e��`%V��Nh@Y�{�����Q/��0��`�T�2x3_wh+܎[�����ڝ:F'��#~@��w;�p;�$96�a�q��6Z����S]�.G;�����MG,:Y4�����nh	xi�ץ��8�bY{a�����ɥ~��o��P�lJ����nmq������,�����4Job�V,���0�rู�?��\�L-]�=�./�ۃ�����3!ϒLo��J�\@�|P��V��ɘ���o��bN��+d�F�nC��S�����ŒXk@��un�Q�3M ��m���s�ǚ�n�5,]�7�%㋝�ڐn&J�º"-`��t�#�@�#YO����wB�K�"�q�7ܙǡ�O�z���\�@B����Vs\�NA�Yє�9��� ���1��Q9�#�d�忊(�v�Ӊ��{������ƽ'4[���F
��"E0>i/`̇��IM��ޮcn5us�r瘷A�9���Z�IW珙��"�V�kO���i^W�ҹ�᱉�& 3V�͈�Lv8�h�E�2x6 u��,}p�IBĐ��\��6�|�ޓ��oF�sJ�iQ��Eh]���'���5�K�@n��-�ձ�<X���ԁ�Z�Q���WI��eLe��?��wDEE9���m�|�&M��klK$JH""���ݧ�rRT�.I�HL�"�����i������R��(q�HS~Wٲz���z�y���Ȫ2N��pv/�K�����C_�Bjz�N5kh�"��J�f��j���N^�>�FDϪ���۴��;����Z� (�+�>iݢ�T'�)D�	=��,� A�i��Ju������x:�tz��
�0TX��'׏���Ԍ˥������`P�rSw��uG��<����b-��@����3�(P�M��:|Г�p?*b�����b�s����|����HN��`���k�nnB�q��ؘ)����_D<X�R��0�rc�s�@D%8���|��~�*�BN�E �D�Psr��j��Z�O����ݽA}J��^'�p���0Z����������&Hd���$r2ܥ����}	�z���L֗���U�撹�
j)!\�s	�!A��ߟ���a��
z�P;��Qd"fAF5Qe��l\��lS�P�L?�=W�j��b> �:g빍�Sܮ��be�4�}1�P=�>��׻M6t��cD���>��H�6]��8e �SG����gԂ��2,K��Z�ބ�� TC1�׭���'#����Z��]"z�i#�lG,���d�5���ګ�l��G�7�+e9�T�3���0�-�%=�r�	A=ҲVZ|-Z�T@�?0�ե�.��n����(W�!7�h�D�hjb�t" C�U�S����u �dkv�����@^��G��mdJ߇
<r�w�.�vnK�':U4���A㒵�l�����rG��#�����Z��2��\x��t~�ܵ���������
��x�M�j䢪��*	��`��M�͆��A���>�H_m�׺qMF]���϶u���˕�86�5������
���@���g�K���/�2����RyU�W�2�_^�Re�Mn�@�A�xw��M����~m���A�#unk$�F����y��:��Y�����+�ilp���%�2�<i�ľ��L;��v[�G�(l1��?<��%�z���tf��l�oJh���5�<M�]�2�ҕ���ܺ��ҚЌۢ�A%��&�}��Ǝ�q*P^��G'�L+��H�Eφ�߈������+�Չ��ā�>E����-q$��iy��SD��a��C&�����:�Te�v��t�������YE�R+:J���q���� `P�u5m��_\��`�[��۔�RB	"�x�v��1�Ȥ
����s���ڈ�z󑮥:,��|)�r�.듇Ե����'P75\ �U�9���ސū� _�{�o>��M_����	V�K:���˗ A�1���Zj�k�`���9�(��>�i��0�F�X�w��e��z��-���	�7Ub�����H$���z�7:�+@z�����6��EmxO�a��G��d�ѷ�������6�Lj�8bu�@�\30ԯF�Em��9���̀H0�����t<c��&i�x`46��]����1��Tin=�[<y���@��`��"4p%�G���H'��>򀻏.�"�d�eAN7<�fP��n�x�Q�Jj�٤>{"|��N��ڀ�	��a �i����US��[+F�k�}��W�-ab��R(J�ꚆRx����8|�-}��+wH�i��&�����=!�h�<|�7&dsM�n1��j�T�(���D�kRv{�+���k���X��)է���p�ZU����~?	���@���!fK�/c�+�Rk��3a�{F��ȭ]�ߒ�2�H�}:�9�g�>���t/��)����Ы �Y����veZKdԑV�1BN�B�Ҍ��gO{q��De��u9B�!u\�:��1�`&�,0E��!��.�/����{cHm�
��;�x�8.��8d�� ��-��3Z�JC��c�*z����=P4Rb3S�Vwi{��m �~��x븩\�x����S����b"IWpX�>/�6����/����Bƻ�FN}���`�؀9�0�- |0$�W�!�CyN"��^-�\
�-(-�[�u�ex�ֵ�~�5
��𚢂�UlAx�W�T�Wg�d ��8�\�,;fu_2f��/�W�$�]ڊ+pq:��ٖ�Pu��f�A�*�?��˝��b�׶kH��| �Ч��*1�_z���/���*�B��^�r�ED�b�C�/H�k�J3ؾC(Bn!�\�B�c�m��8˺;�'��g�ܜ˿ ox�dD���}<���U��8S�"�w����6�dib��Zo�9"�]#g,�,�2����rU�j��K�K�U�Ov)o��(��^���O��VZ�]��C��%N'KJ�1��kH.���}<�Bs%�υÀ�%���9�$<������W���h�S�����)l��O9��~h���$�w����LL�7���S�^}�MNh��QR�_�x%ƍ��{�F^���]�{���xR�Ǣk���T�.Z㬚�_^�
���g5�D�diĠ� zֲ�oc�g��X�.㌧��eMRnkK�F�FnK���wM�*�L˹�gf?�eOU�Y&s4�c���[$��A2��΃���h+�����z� %�bHg�~�s3�AAD(�n�p��)~4������uQ^�Vш�Ğ����A�$@�������ם}>�����c�~O�2o�1TD@�`p�����X�b5�2n��������%�s�]�x� E����d �`(�����O�[ �*R������0O�Vd�Y<W���&�ZXc��$����A�������� �;|��~��P�ƿq�f���^+͘Թ�pΎ��M�U�oh�4O�66=]�x�)��p��;���� $ػV{-`�wAJ'�]?��	�\����օȩ�S<�١입��2<����}��柺�%k�o�f�j[��IK������o��J�s�_�?N\���9<"����SG[�	Q8������d�ɥ;w�N���,��i�>鵆|��2�{��y 2��+��
�E*b7�XRq������2,�9����slQ�cI�屵HY7��<�\�U�ޛ���|o�S��)=�� �П���1G��/�+��U��;�&2�8���ꒉF$=|�0�eÕ>��*K��.�o�lf�K�:�V�t�Y�de^-�U��4�m�ܜ���)�
z^'�7g�ۻ���k����Du�86^6�I����7�u1Huו-n�q^�ꪴ�����X����d��5���-}����2���������ϢA�m��z������>��?����W��B2��$��bC�[Z���0�m��z�Q�QX��*���E�C::��)~ޕNB���C[��1�(�F��`<�Ʀnq7E���R�'v �_��)�P�H��k��Ұ�8kn�9zYPϼn�r�t����!D8��F�D_��쇕��.e@CE	lo��)��/�Qޗ;��ڒl�QΒ�{�"��Q}n���.F�r��阼H�d��9�P����SkEsX��[V�pv��;���j�X�o]�J���Q⩥�\�%���u��]�f���X-��iy�hggSY��x]U�7��Y<<w�Nd�L]�D�]��hE��\Ek��uI�IA��UЉh���K�eR.c0��4T�����Y�	�Z�#��t�2��\��'&LT�������t��Oa�W�:�ދ� =����Ll_FN#��| C�8�ß'�l�����Ь3E#2k_i��A�
0$�Ծ1�z !�o���8Lp2$q�u�r��ʪ=���i0���ק4�X[kL�NB?F^����Ξ����<�;�о��l�k>�`���_����e7���9���^f6�1Eǳ񜌡�/

�d�zp/��$z�S�t.�o�bK4�t
g�U�Ma���E隂��� DW��d�'�Yi� O���L�W�4ԥ���֮�)�%��[*��$٢Ħ@�X�iF%�J��d��ϟ8K�&f�Q��ޖ�v)}��5z�Y��6$�N�l��W������J�N7�W)6JE2w'-������}��Q)�
e�i۳�j$c��`/�h��Gђl@�[l��}��J�^Qr@�X�>y���@/gz�O���$�$O2S�+O�0W��������v,ln��w�m����Q�AY%����)�r�$@��mE�e>��-�mQ��q�'\���0�'rp�u�颉F��5�u�3Ku�Ӏ[��:�>�1q�� .�C���s���W�s	��	�[���;e���(u����?�BL�,��Ǹ�@[�bu��`}��X�b�	��*�Ʃpa�m�����D�ۉ�u�%y�[G�x���ϱ���{SB���gu�'S�5B�I._H��!�A� �lӅ�x��Σ<��0XЃi�D��,:_�6�5�9A3�	@�|]���:V��J�^�쭘�� fУ�[�EG��l�����@�E !���8��]�/��Y����]�̎0$�y�%<�ˤ�L`�.q�2A��N3���ls���ii�����"[�9-4�zvTh2�����IDYxٖ�ټ�57��^	��1Ǔ[X���8BE�������u+J��Lt#C�t+�o�1���?�UXU1+qϭ�\٠��Ý����y��i9�7�jnP7eFi��� �r'�^��J�u��W�a`<4_j��/�=J7��ʍ�@7&��$�g�N���C�i�%�bx�Wq;k���:�����0�F�x�bQ�j;F�*�J�6a6y	wP�Ԗ�J����	�*�ۥo���%�ÔI�t�75��ڨ���d3/J%��"�zn�A�Eq�h{r��5��b	1��S9�ދ���WE1B�U�#��#w��R{��h�=�ϑ�˚V]�i5�,�r���γ���Gb��0�q�+o�\�x��'6K��x�]$��/m��l�)�?=��:����nn$�Qȏ��	{S���e�}��Sߍ�UE��(�?jj;w��w�~���bc�w|��}V�x���f:޼�YR�a��0h�h�Ok��pR����� �ñ��C7G����|y�����c����v��y=�2<DR�Th�t�;��I�3���KK\k99n9�Y��S~؇)Η`�!���|ѳ�X�M��0U�m�n
czJ[�X�KD�+<x�g3�6�ڎ��4��y��r�彛��j�W������2�K*�]<����;痻V�?W��,�vx�7 |�g}�e�\�&yO.�r
��E�8�"N0L�ANߟC_T�q��Z��&1c%Q��j��,bg�G-��|����fl��-V
.CE��F�m�xsESM#�fۏ��xF��)�E��j;��*��"T�v�[�7��7���S�ʍ$��b%��d�3�Au� ,p��l��_�;��cϱ�s�u�Vj�0� `�=~񑥓�q�Mn�`s?1]��;˯��˾<#����t(�$X�c�l�o��efʷ���e0�B��>�������0��R��ɷW=j��C�Ԙ�0T�".���B��}�5�P�H @�6mgT-A�lP�i;c���18PU�@69xM�0i��>L� ��r��Þ���p��Tm��{xP�x8���<�Yvmf�9͑��% �~�Q�s%���|���Qe�AP��ϓh�_:�c׵�
DR>�ß���Uq�Q�x�U��K�uC�$�c'�',�I��zV�5F�ƣ�P�7�$'9��9��Ι�xi�e��F��-𑘳}�>�^2H�q�PMKک���� -�����xd����e�Fg�nK����+��{�A@0�/խ$5!������!��:�����0g
j�Q^��"q��
�TZ`��$�"\(��L�6-��Zbs�5�C	g0�e�F�B��r̠B�@�����q+��Q�TWaȗ���0$Sѳ�����CZ�6�f�����>�ԅ��jƔWA2$� f vf���DvHuf
/�Y�"!0;�ؒ�&�	:�W�8���i�n��i��4��n�I2@���GO�11 "�5ハ�%��t�1��;�z��;bh��>V��������m���PX�
���G
���^)�Xr����k����)�L��:�ptV���e��L�o�*n��w��ң�m��Kg9T'f��j�{�����;��U���HCz�y��=�;�$Sѱ.\-�1��]-�4Zi��U Tֳ���o��|��H��M�b5�`ֈ�2�RN��yG�v��m]�V��{:i��<
����C:� �H�q
[KE�d���\� ;�6�pP�z��1�՟��,HǓ���)B"jH6��5���w������'�%\a��&�q�$��M��V��6L����i+D~��/�b}�y�kU��'��(�"�Pl@����v�?�d@���zH����%i��8�¸��n�G���uME����ϔ�d8֤|�S��+
��I��{�c��iD�us��-@��M�w��E�!��IA�M�X.�»�{-$���et�����-[y�&f<�C�n�kGCܞ�/�`���(.?�S�&l ��(�	��m�ݓ��p�]�	�KS�Pz�:�j�u6�ֈ<����r�OKY/z��oJ���Ʉ��	/WL����;���"��g����I��ʎh�0Q5���q(�x��_��އh,TdX��� 7#�M�N;]x�Yq�W���� ���a��>����=-KE��#�q!iE�	�!f��JM�ӕ��:3��N�;� $.��Er*��":bP����[�Mn@q�5�,Pmd�&$���C��JE
*"��d��3(���FaZu��H���������t̢j���nj�˔iGOp*tC>����\r�܉��ح�vp��V��ȸU�Z��*ҒN�'8v�Q�0�`PX�F��X�j�Гݍ�d��v�P�W2k���R��
���5�p���J-�F�~� ;����G�ů�u�h�V, �[&C�R`�������p�$��.E�����)X[�-�ۻ��P�G��&�������,�GXߋ%Y'������=*���ac�xf��F)����8����Ɂ��;����zJ���_�,�A�J�B���?�#܀��yx����S�m/啺�d�ST����es��ԆJ�o5�7oYg����8�N��l�Ҳơ�.���h�.��2 hӰ"h��4�HF_C��Q^�"�Q";qr���ժ���-s�Z
}����3��(9�!2�*�pҭ��&�;����8æT�k�]!��/2u��A5�+�^��I��y�Y�_����9�tmf����="�s���\��P� =�~9b}�'?�>�:���s�(�I�.�mп�+�^e�L�a/m�c$JW���f"0���
T��p�3t�
����:��}){�����Q��S�z,4\�*��B��΃�)�{��՟��p#̢���#,��!<.S����
��-�#:��.|�����z���2˕���8�$���bb˂�g�� �,�� ��>x!��c�V;S����q�T-�������20��,��M�H��x��#F�V@YBS!�g? O�&:����3�ų��mFj`!w-ȳ d�ِQ��U�.((��+r��I�h\��ɱN�w6I*����K�y�xv���EE�Kx���u�M�3g�?�$��-���H�x���[p4fL���`�z�ϋl��Zm	
�?�J$�6ΔV�ˇ�.��i�������a�ËJN�@6�6w^���2����|��kż���E)��mqA
/oos�m~�1��� �@���Ԑ���'�D������8�N?�̇v8�|I�P�Z��Zv9
�O7�O�G	*���kF�T�͛�x=�B;I��_�K��0��S��]�f��џ�5����]��z�=�4<��.G�{��s2�!S�EV��,�@�s	�f��d�������M-�&�ԕ��Û���7�+�}N�)�wz"�_��ސ�:ղr��6�E}�26l���kY�g*-S2R�?�)��<j�۝��3�E/�{�.s�؊Wtaܹ2`Hv�I{�ꁋ��lDN;~0d�;���Co=��;{RO'�9Z�.�p���C���b�!�'�#��][�̓�~��fy�5H��F6J���Z����y�ݩ�|zl��؟'7L�K �`U�8t��9�0��M�;U�D#<��r���wI*�]�l�N���A��v���p�4 Q�Ʊ][F3%�m\Az_�2�n'�����?G��_��[� ����+��)�6N�j�^3����_���)���qyez+�%O�	Q(B�\ؠ{�r�����9��- %�_^jw������nO��8l�^�?m�zt��Ǐ�������7�v��P�0�*����#�!2����BAe�9��):^���d�u,�J��=,^�7>�Ig(���މ���C�Фy��bNv�i���)m8'�����Zða�ע��:q<�h'`45�%�H�c
@��A��$���T4D�0�<JO�9kMP���>3	j�_j��C�D�!�=�F���_0&R�J^Ls�c:E���e�
�=ɩe e�η�b�+h��l�
��r �*`�]��o�ʟv�PnPnT��ɭ5�u��lT��Ud�P���Ϫ��i�o�YT
����}'z|\8&�������V%�ڂS��U�n7Y����2����q����0�	�������(af��6�lV�q�&�x#Z/����$,��ը��p^���j��!C��љ?`���I���5����"��n�4L��W1��P��Sf`$/ϲ@\���۶�W4ݺ=�F(R0�d���ڝy���Բ��-�g=�Y���sѺ�(l�p��y{I�\��޽�j�T�1��l=e^�Z�ɀ{(�2��"�L-{�X9�v5�L�o�c]���#jC�D�l�&��b+��N�,�=��8��ٹ��aO��\�P��3cWo-eg�"T��Ͳ9a�&C{j|�|T{�_S� �CV�`�1�� u�!bC�n�j�{{|���OR3��2m���@�o�e ̰y{��U��]e 	��r�����rE-� a�H_�1��F���ʆ[:�B1>_�Ma\X���:���T�����������]����)g{��ĥ�(>����۵)�!Ә����m.�+~
;����+������)oeظJ(�qLpx����ݗ{����^�I�rYΨ�����W�����Y��6N?���G�.�?v3����lG$-)�O�.I�aX7�Ӿ���U�%jy{�RC':�}�p�������m%;�8��ν�X�H@���s#j�;�[\����s����{ �� �c�Ջ6��2��2�����tq����	Ξ2��pW�~�}� �Q"�́ۖ������[���a/��B�lln�*�S���M�|n2~�)�s�Z��P0������m&t�6u����8��O�;�r�.���=n��Pj�iȈ��x�*b�tcq@5X±���S0�N�,(���hw]t�[`���.��ë>���P-Zf�������X���n����7� �H2�(��/�z�{�a�,A��2dy��Y:�L���$wb�x��o�sj�Ճ�)=f�?�k�q���"�b�|�A� ��n]ز����}\&|�	>�Sб��
Z����}O����J�x�����!āϼ�m�|���U<�0F�E�Ѹj���˚g�H�C�k\SLx�`͊��)d�g�NWj� DKQn���9yŭJ�C���V�������8�D����Dr֛��8�� ��]B�f�\���{ė�0����F�B $ '�5O_KLi/�߽q@�Q3�h�pP�Y�.���h��g"�#g�g�o�ř��^��O��A���l������x!�
&Z7ob��L�:��G2����<z�+��'�<Bu�;7}{��桘h; �|�!��4���Ǟ��\X"G�Z��D�,�q�G`PV���G���liF:B�.ɳ�6._�pMM�"xj�w�F-;��X�	m�\76�8T�;��`d�����s[�W�W����lf��Ս�S�`�y���%�Lu���N"����,3�l\b�twd�Vqn/�7k������℁� ڹ�2��/pU�B�>��'�s �x<!�@��A���*fp30f�����D�~^�ΆX�Mn`\UV�a�w��)*K�[6���U�'8�e�X��z ��蕘���[��\�QY0�����dr�	9p$���0�����m���/n�px\LV��G �P�z�cII{tq��6�ɂh.Č����Ic]f��}/�����ݶ���A4��\O��B�>�V��s�;�&w������A��=ڒR%}#�f�����eo�2.ㅥ�",�vȱ)�ۗz����Xc��Ke3t�L����T�����@դ��R���Ul�Y���8��o��� �TEt���!A#�y |�
v ˹Qݲ��*�A�����Eڏ�k�ΐ`h~���;$�Ok��R�fkYBv#S��?d���Z��;V%���=J�]I�y5|���H ���sj29��UD?�bI�&�@Iq�ɵ�����fp|+��0�h��Yc�Ա{}�� �oDay�T�Q�Њ��n�S�d�?6��K��!�~�_x��Ȫ�ն�{�)&9�(7�h���KJ�-7:q���K�|�goM-���Te�����0�������Dp�b?_ų�y��2����AbS���ŉ��Z�8�����M0������&���U8jW�@!ޜ'N�z*(m\�陛��$�^|����5!d0�w���b��Z�����!�4G�ҏ+���ފ�P�k0�R�[�Wo�3>jm6xx��������}�q�����x��:�hǋ���:�#�4>Z�EB�T,.�-��a��F֊	��ӫтD�srG*���y �lI�~���f�z]y�ͮʯ���#�_��]��������~.ST̀s���P�0�j�-��#q6�F]f('�+��n��v�&�a��>Nv2(��rկ��2���3h2!���zQ�Oem��%V~U��a�f�6<�.3\������A��a#�S.�I�
���}_KkeJم.�_S^}(E�m���>�����s��F���S4����*�6̨��f���x�k��^2�zMp�%s{L�Qs�,y�#�a�Wfn��+ͯKN]�����V�!�vLф�����z�B�����6d�2�}%��8׮?�E�A*I��la'��18�D4^鮼[�\�O�����vQ	u|/���l�tv]o��Փ�̝�:���}v,'r<*rI?Oi���oF�����A�l]�(#-�>gR�D j�Z]2S��r�-hZ���rF��R�6@Qߔ���&\r��:BZD�
�/*�D��� �rg�pY�7T�m����ѢJ�7f���\M� �fF����w0�%��U:;�;s�T�/���"J����h�Yy���#�==�1i�A�#h
�5[�&	��S�u�;�����6�7���d!J�V*U�5�龑�Qc�]�\0�\o���cOA�.x}�eY�c���$zhh�z�+��4��k�ߴ���`8	�=i�7__��� ��<VW4eyFPs�:�
�nȪ42�����S�0r�S�ܐ�'�w����
�*��[d�*�ѻ����M�_���bk:Z<M��F��I��+���_��1�F���'��Ѽ#��:Z^H��y^2���J������$o8˝�*s����3]t�~4REi�����ȞxQ	��r�ᔑի!���+�<�K�@-�r#~᠒	�Wr�q�a�Z:�11�rBj7�[#��^�M}�Z��m2�|ŗ���o�"{Г���W�Yطc}"N�3���5�hM����Ʒ��ԟL��cLF�l�ԳK+�L�������I�u����J����S`��L�N;��6�'��xc���|y��-�;ꅚr������
δ��t��y2�4nJ �@j��D�Tl~d޳'`؉P�W���	��T�pqh)7K���j�c�����D �q��7��M�	�Lݒs^'C��&�B��R���bŵJ�8L�v� 󪟔a�"Es�o�Բ�E���?������l�������%"8),#�B����F �����%o����%��f��6\8{Y��|q��4؄�+�>lۚ���tWrq�0��B��g�dLw��dO�dc�	2v(� ?�(���@���P1���O짣�1�w��۟>O^�*���d<XT����I�7P�OWR�Ǵ�򋈷�Jټ���%���8�̗��M�:�	;?�·�w��W�	Y���mm[��R�Tt6.�`��܎�%���E�hō)*�G*k��f#))�</��۫�W�t������rBl :��ƧN�!�V��ᅱ�R���x�h������p���J�K�]U�e�<���@'�̊�t���G��]�<H��z
$�ҁ��X׾�k4φ=k`R��S���H��V��O%�N�B�M����������c���T��Xw���ދoJ<b�;��Cn��n.@�Q�
�u��q�xr�w�sgR'��?�C;�P�����,Q1 IiY�N1?�$ą,�1Ze)灿������zy4+z=w4��栀*�g;Y�Ɵ=��*d=��N�q���P�B����CV|z���$���uu�������\l�qaZ�myo3ROY������M�V�6�����R*)�	�]��l!ո火���ڍ��t�����	� '�v�T����A=��PO�DN�T͢bē妡����v��4,ӥ���iʳtH-*�f�	��E��PC� }�����|�݆�*k��|Ӆw�+��5��^�[�I�� Ub�;�U�����U�����4��%�@�_�y�zs�a:<�+?y��s���׫GX;Fd��J�b�G�('Ph��߈uȏ#kN'�6�
�A�$�;��qo��(9��Jkl���F�Π�A�!et����/~}�W;4ܩ~1�(��uѰ�B�`eOF���Qyy�ZH�Љ�����g)d(,(����(��z4���i5�:������B��2�Ç��=^�&Hp��/���+I��>�Ԭ��)gyH��~:�P���D�Kѡ�=���E��5"]��K��<٦��� ��t�8g���	��ȡ���-J���pHu	rS���F>�Jx�p�VJ,� n�W�˖�	q/0�sFԨ�f�¼B8b	 �v 5y~�e��Z��+Ȋ( T��&{Ļˀ����ʻPWS�L��/72��u����5��� j꾢|a��U4�ŏ�����U"!��;qi�Y�^��u8`�JrƉ,sGs%3�PQ����3t�N����Љ����8R�c���Гu,f��8�lp�#�\;����U��_�X��rjSl�ǧ�lV��h���K���޼����K� ��(oř�]#B�f�J�7$�=������ӡ3!�8��p`���޼6��:(��5�st��,��H|����H�}yy�����Ks��q#�vw0�-q\.A5*�+�[�_UW��<t O#V��}\�k+�e{�h��9�/���L�ue�������<к>�7��S���E���
ӭxZ_,�<|��)�7���W>������\`�F3�T`�P�X��e��b�92)�K��Yƞ�u�PM�	�A�XA76?�1gnϊ�i忡	(��>���j]��Q�̠�Ǡ�D{�Q͓`�X�
=%1!����Ժ}�E�X�=��¼���1�]p���)C��%�������Y�!DA���_����zA1�3��:�|��ʯ,�W��Ç&�W'��"�,��\ټB/�V�?�_�=�`����L����;L�E��vĉ��&Զm(6��!���5�g����ֻ�?7�G�U����_.��1�TE a�r`A�a��
�l�B�<vEJ�|�*�v�w��Mfڴ/
%'�g0B.-WXMe�Kuv�=��/�R�q`"�[R���/��6S(��Yf��ń���Ȳ�,j����cnR�J����Y}0��8��ڌ�-���R�Is1��lh�|�'[Kظ	�6�y�	m�*�#O]Q�~���%A���@�E$�1��8�>Bp*|�eڥ⭧�eri��@V�)�B�q�ܰ龷FT�+�"i��w�'Ͻ��x=����(�����1$�(���A �=�0zd���n�5��I���y��)f��Vq #� �	�g�`mˤu�����+�}@
�R�x�F���<����z\M�`�s��5(�d�G�jo(}Ғ~2��_lN����9nS���"[� ��;�Z2�Hg%��ѽ>E��o�8 ѯ>+��)��U�@�Q'��4��Ԅ� ek�2�Mp�5�wb�kp9�X�Պt�M� uW�i��PiNɡ��3��ؒ�����3�2`B��ѣ�宊�%���~����C/ c	�D�V}�Ώ�P��v�iP����剁$w��%�����Ya�֫i���MPh뻳0GS��.���W��+�?µz}����qj�݇Z�珚=����N�ǔI��aZ�oY$�� �y���DRZ1+�c߷#�8/�PO�-GvϦ����}f����kw�L:�����2��av�'��@|����mN	��Ș��ܢ�w�%C��)0X����s�7���bG�x�Ӝ�(X�p	i�.#b!��>YgPᲑZv;�+�r�^)����0��]��H �/ai6��ݲ���JK\L]$� !�p�+���d}@���!�u-G�(ɛ�ݲy�r�U^������x�e�E�}= �&�qT�_�eD$�P��4�ųЁ �X/�d��]?$]�"�Cb~�ǩ�K�-<!#ok��>8e+�ä��:}K�M��$���`=������s���\�8�1�K�;�Ԧ#�T�*�`O�@�+?{t����{y+�Nh®+��:ʩ9��jEWyeS0�\����]Xj��7՘�e=�`It3đ�p=[65~���H\9Y*��I�B�_�\�����쨄'��dUj*�?�� ��e�/��_5d��1~U�����[���*�)V��|��ww�.�ſ�ەVC���k�˨��'�g%Y��3sKm���~}Ϭ��R$�ߞ�{��Љ��
L�=�N���1�����:G6�EZa#��8Nڨ�Z�__�ő8��Ad�>s�>���qr�e���ZM>�XЁ�F��<Ti�C,x�`��,���<�O����A�:(�腡���&n�<�M�\7�
!�L�D���	�Y1|[�����R��A�n#���8x�X9��mMa"٘�d��4����n$22M��������'�J��^"��]e�W�GY	]���x��l�`�!��H^ނQ���x�{�6��(��S�{u�y����߲�w�R��?|c�cs���"�">��[���z�^,Y8��	���򤆝ջ��EN�Qj�$>u��+���P����I�U\�5�SNE�XN�̤Js��슡3^�ٯ{����r��Y�8[B����`����v@�:tk��������W�Y�G,�1X�{A��,󐼎��� i9¿		)`�Z0*�J���H:�� �pk��rai���'m�g��oN6�^�~\����,U�-��m�u��`�n��HL�'������ѭ��W��2���������f�����o�>�N�T7�^���C�o�y����ҫ|��I}1(�'��>�ך�K���l/Ď3Q"����_�H�G�O3|�����S�2'*R�#8¢�'[k6E�����mut��]^?�[���7c1�Ta��nGϑ�}�����h��1{۲�ʛ[�fv�U����h�dDr�d��f
�S�9N3��;�8�}A�0�p|�-���sf���gw�Xf�[��Q�4!�
u��#怢Kr%s��G:5g�����Nd���� �&��J�"�=���a���P,�σ����^y���W���v3|Ì���� {�	r�#�h�h�!"���U�qCC��U~nE�b�/�u����F�s?F��b��> �>���b٩��Vr�6�6��|3����L<�E�3�'`���v���$t=hd)�I��3&��Z���]@(����9]�le#0�O5�" ���Z��m
A��-U������▰fW���\�D@kAJ��C��}�நQ�k�S�ǇPE��"�?յ>TE��nm��|ʊ��b��p-k����в�8�&��6���/&���-�6n,;3�bS�k��;�r����/��Ÿ�$�p}Xn '@���;ĉW��������ņgm/Μ@������_0�@ǯ�"��A`��@d�F�?��Gkc^-���l#�����!���p<�k�:2�D{�鸸}�[����_]�7ku�"�*s�$
V��m�_�`NC�"�5��w�4ķ�a��f���3D%r�Q��o3��RqB�;�T
��7t{�1[@r8W[��V����SG����E{��ě����]���`�z��w��>^�<ek��q�h��*�a��.4Q]�)�ow��̡���������m?�?�����P���%�5�@���yH����'�5񦗑��:�рV8(��~�B����|�@l�W:U�L-��zv]Q�����R��QV ;���ƽ�r�+<*���Ή��g�-Aˠ{N4�瓵M�W��]��}R�z�[G�;'��{Z���f�;�����1��4cO;GTDE;*�M5��M�/"�Hzm��w��먛�4�����aO�}�U��[,��߻s���[�� ��+4�_��͍Æ���(������Ս*�E&�g����$S���C�)+��#�>�����%L�9Rw��ҭU��,?&�!��ܣ�_*�8�
�Z�a���;�`�}ϸV���茦���)Ut�*A�T�Rங��ؾ	�|���Hp�!+�Q��;g�K�X��C���a�g�P���.�i�qf��9�"���n�iYg.���8���Pe�r��2mlU6Ό���ŢA�}=����YZ6�A,�6<r��ǎ��� 紋F
N�
ŷ�{DџŇ@���W�f���6y[����E��#k]n�Y`|��J�v�:�r�2��FŤڵ(0���F�=���E��҂�U�r�RM=xD�\�[��!����F�ަp�x�����誧���'�R�S/�������fa���<��c���Z�f�	�b�R���K:JA�Ӯ���N����P�#p��O�V���BH�P���
h؀�OI)���0��Sd��'�uC+�C�L]9�-x���x�s*���X8�R��{��o�}�K��Y���wA�	S��d޳����hKU,�oo-��$8�kUÞy��'�4Vq�ܣtmSj$��c�V�����h96��Uwg�����e�q����2q^�OY~(���e>�
l�V�#�n��Q�s85҉�GJD8�C���z����h�R1�'#	��k0����K�D�gM�f4��W��C��rܬG��n�^7&�_��y~[$p�m��y��NB��wr�%�*�&<-���旲�%���:V!� �9TU�G}o��O(����SJ	:d;�t	�bң�ȑ��/g�{K�YHoq��)?�� RHiϲ�78�����B�y]S���-G:�c�b�_GE|�W)���G�ه'1;��?'"c|��]�t,09�JF�g"5��h^��ˁ]�ݘ��b�~�S���;'w��Ӿ��ȳq����n�;jb,;�B�:�˟��D;�	��=�ȜR+���js�4{z�=�Ė�tP^J���Ó-5��V��tԲ�G�L
��C��,ȱ����B19�`������z�E���W4w��m�r@��z��>����`�B�wZ��8@����H�w��ʦ4�7��8�����9�м�nEɼ����hjh������\4��+�qɮ���%]�Q�8����X�kQxK��:��>$�,|^��莱h�W�Mx�\�������:�]�刚aE��QH&𡈘��1��q�$_�g�T@XV����3�q�zT}��D/Ĩzfis荸��$,~}б*A�:�U�`πU���!�(�	s>����XA#ߌz�#;E�z�P��7W‥����y�]�[���og4!��kB�M~W���И�\��S��2�����;w��� ��;Pi}Si��v�:|�Q����;�"����B�/���m����D�)�+�F,��K�?>���0\�74l��̼�dO��NFj�b�"�.]��#WCn�������u"�uʫ}�!�o�K��|�W��$�mk�����;"Ѯ�ܴ%�g�#u��p�6��E�{�KL�3����i�����D>=���/N����?:!�'H�#���V�e��~����|������eK{��.���Ȉ�L��,�_�Xl s.9�(I�np������[<^�~�((�?�ovn�LټGॵsw��p��	�!(��D��'y��͜/l�Ѣ������l��I~X��)[+��C����Q}*~k}x�W�ßFA$3\B`&�F�T�r���N��*�^O�]�^��8�m)��q����N�?�3�/��_g�ڎm�$��Ҹ��
���`Me�'��r�a��ŭG�-�P�/�&9�z'����Si�*�w2�ʂ����{��{�\�%Iġ�Y��n-� �>�[��O��X��E�>�
��{g��'O-��B�g7ʴ�Q�vp��.�i���T� CQ��S	�Bc*e��ډ����c�G��%�8τ�)]��6h!�R��&3��I^�	�Q��N�j�Bv^�u���j��(���\L�!�7lIS�!��_���há���5bo��D��#U�yR��*T#�.�#se^#(UB�^�L8�N���n)bE%�0q�\��Ċ`�O��n9t׾��I��m'݄�����*bܼ�B��ƭ�\X$i<:X�M�,J������g`��:Zl��RȦ�w��{U̮��G6�z��ހ���g���ԭ�	t@�$�׮�|�$H�%'c{eI]��d:�I�����|��X���Q��zu���@I��})Z�6Q��6�2!'i	����b[�PN�X �@��w5(����Iw�R�OG�
�1	�ߗ$�$�P��X��E��A����\�VO�U�P`+��ar���0@�ڡ(a�B���>���OT����l@�iL������ni���ߋ�ç�V����3��� ��i��(=Q��V���d'�E�/���k���lׂ{��'��>X�:6�5��c$J>.<�i� ����r=R���q��:��e���r}F���|�h�+�G��Y�0C]n"Q	��"mLoHa`9�&��@R�����$�MYI��6wl��Wެ�=QB:��l"��M!Yy�ݫ|��u�b����
2�z�  ���b1�i�mr�+5?@'¼R?_��P�v��r��CG���>}�D�&��W���s���թ��1��j�=	�c������1�G	<O�!�'XE�d8~Ǖ������ ����|�ff�g�t2�vZR<�&��?YZ�����t������l"�U�i�ʴ����,亦 �9vl��H�%go�>��3f�{D���&'�E�8�E����t-�5�Ɔ�l(���h4��uOm	(��Ȧ#����=2[�:�V�EdOr�R�y2Q���t��
}�7�唌��x��Jr���k ~n6�:�[Mn���$U�3��D0�Sq�1N��{�P���=��)�)]���u�N�A���db��#>#I"�^��9f��y�{�^wXx!ZDnC�=l��3D��=.�.��c2ID*��yېd����ۖ�K)`���u��IH�ssO,r��$JdL%A�)���A�EB{+X� ����+�V6cK��Woq��t��������F���e֡Ɯ��v�q����]?
���;���NH��
#���Z�)Y4����AB9�� +�'�������
I`?�s�z$��S�� C\]�N	B�˦g����brl��eW!R%�U�����ꪆ �T�,ȟl�=�9�> �;n�C�����9߿��R>b`���|f��W;`��}AR*��p�og{!�DBfVU�@���_���t	��Yu'Lj��/�b�i� E����f ��*lX�.������a��Z��Q"X��8�#G$6����Cw4!6!���Όd<c�� {TO#.���T*���^$rj�� ���,�������V$���ʿ�⢓c��P'��e�u:8%�����jԝJ�m��6�k:l�e��{`'gNF���9PlR9Ն8��V��Gv��W�E(9��.P�E�����a���ti�J�D�T�u�����mRۤ!�dJH�p��s����8P�������)q���#/��V�K��=>xyJn�Y�JG{�G�~�Z��SՑE�>�ּ}-�h�ajY���k��-.頂3��w�2S�GD��ވb�ILM�E���u�����,���zɑC�Lc$��˝����u������<�0��������c���5�~\M�[�,����F�'H�?�ǭd(�a'X�S��.
�j�@V/�RoQ���͜�Lrg�6���,�"M߹�~�z�#Gz��6Ie�@�O�Mzrqb�D�	�L^�;Q���Bk`?��[P���r�ة�o�{{����_!�b�L�r�V��B���dF��M	���ˎ]ԇ\&fTƕǵ�m	��>"$�F-E��q�dt� f`@,H�K�
\IS�"�Q�d��fّh����n�r�ީ��N6�J�>}�j��E�4����P�P�$�)@1= ��������[�Y������d�z���sD�S큎�l�n�R���E��.���xRȺ��cP<𱯻�);�N��*۵$�	�è���W��.�1)�>$�����N�"/S���6�_��S���g����c���s������s��B��L��+��[�3[��wഒ���:"~����Y��/�X�M��;W,7?t�����+wY���ߊm��=�|�#3�9��4��`�tC�2͞�/��0�K�>���m�{:�?�oj��A��X��h��H�!S$�i�}c�� {/	���i��A5�f�c�mj�.�SV�n����e[��f���6,�9���ek x�j��T!��XLc�O���|Bpȼ3��e��GⲘ�\�*���e�L�9
�?�
k3�boFUI�Ḱ��Dܸ��d����p�8�:�����X��\����)!�R�B7#�5�"ǃʕ7��d:�oh$�?�5����b�\����j>)
iv�=Fqp�SNߵߡZ�<d������ƾ����'����"�ʯ���*_:��*D�m��PU��.�s�^8�<�Kӝ7�
��-�([R�H��C��V�/v�l~f��r�Fr��,�]@q��h�@uO����7[�9�Y�5?�(���7��&~ ?��meM��[�[��I���J�x�n.Z"�G� �Xs"�#���le�Zwf��rD��<�k��	��^�B��.�bg;eX���mDړ��pQ�po�qD�\�R���w7��u�]�2��j���7����UՖ�4Rb�S\��轌�s��)�}B5.��[DS8���h��=A�����P)�Dt�F�Hx�o�T>���d!�؝6+���{�o����ec��O��)ٓfƋ3���7u�\m�h80�lw���d$!0���Gr`���x��r��M��V{o�U
�XR�� �U�	��Ĭ����Ȏ�p�γ[�Y��9�}]��)�F�P�k��đ���� 8�fk3Y(�G=9����polv��%�\#��b���	��)r�a�?u��H~�4&h�b	@�"wD<u���1|-�����\H�N���Ff��4鬷\Epd�!Edݻ� Woz(�"�g�A*�
]�8Yuhzq����z��;�$xGz�D)$���)�*Vј�[�M�:?��v�/~���)�+Ʒ�C�Z�,�~tO7��*�W$Ԍ�_QٜD�m�R i��95j���'�#�~�h�(Ĺ"8�:����C%��n16�9����g�
�J�g�*���	�.�'㷧~{h��������:|)v ��>�O3A�����1(D�ʚ~��t�IG��%5�#�iEd>:'�F�١�I����r�����R�B�|��V�JFG�c�ڐV��}�+���D�����#��T�>ǐ�Ƨb�ݜ֩�����-�h�z*A��h���}��n6��ʨ��}��]�/�k�)�9�<=oj��v����PuT�M��v���2�%9�����9�[�j�;0�P�Q�!F���������x�C�������Z2+�!���R�c�K���E�� ���h���2�Hk�]8 {wQ=���Z�=h��2˟6��������EZ`�/N^��M%2��n ��3�_
fp"��-s%��)������}�M�]���1���4�O� ,u��S�iE�PQ�RQ�eme~�tY��(��@�)�����̉�r��4g�c����Wxp:�"�Rے�*(��p�t�4՚@{�IA]�tkO�N*��`q��Rn����ebֽ�K�!��K�nq?P��y/���\�MwZ�uH�!���XS��C A�T����_�;8)�=�|��*YWmq�&Z��T�?�^��py|F'X�[32zu���y�������rizX!Y1#�`p���^�0����'�Zٚ�S�)Ά��bڦ�~�x�6�f?d�8c��Q���Po�=����<x�&��%B�H��e�q�ԦL֌�"߆Ly=���eS�K���$�w�Nl��~!}QP���D�}$��!�TM<��xb�D¥���_"�OZ��!m��lg�y�/�^���öms%`'H�*�Q���"!܄y����?=RBKEs��Ȗ��+*�Т�!��(w�U�M���R�N�3��$�y0����������[��)�k����{y/L�'��D�8��Hczk$�����y�
�q�]�!����[���ŻZ���A�k�7�S�q��D'9r���TC�?�b<�nn�"lb���xj��wk]�8�e-7Ōp*�p���l0�8k���4�I�8�&��~���ǪeqC��D�Tu� ���D�����5�H��:���L��-��q��R(��!7%�*��m����5,R��`�p�2�7�_���|����	F
2����O@f���c����E�G���?��u��P��1D�S��?���/Gg����SJ�x��\ܨZR��Ro������5�o8��#��6%.���n`x"�����Y�ig�rxv�E��G�~�mP��)f�@���@��׮���؋}+�y/�����ds���2ic�!��UMHx/h�;t�L�N�d�B�G|�0/��+�:�f�2iZ��4ƨ���)F�;��gԄ
�F��,Bx3�iÉ|������+�0�����0m.�·O��_���5p�.��yA�b���LW!�"i���Jf��õ�s""��5���x�����7l�������q�y>/����0a��x%�w>�.�Q�8X(2��O�����aޖJ\n������O��_���㑅�6l��N]4-s�v�����0���}��	��9��5�R$d�t�|�	6�H���n#`a
��Q�W9���6��:d
�6T���܂��,kf�.�2 ��� w��g�Χk)�Ό�������k].���4�xwe(E���Ȥw鯔��'D�cZ���A���y��wV�@-�v�yg\����p��6`�Jb�ۅ����N�C�"��8>bv��a���z�?�+CfI q�c�s&�Y1�=T����>u7'|�-�-U�cDˆ��Q7'�M//�uy��z��Y?�2]���t��7�\>wA5�J1˃�U�bO�B�;�RC��pm�����6��0T��vv*Q �c����p.uP�]��Q�b��xu;�߬���A�W���Ҍ�5�h^'P���[�kc�k�Y��&�1�V����Y����r|ўzD�(��|}����hĽ%5t)��Ӟ�|$����q��¸oOtj�Dɝ9���K|�0��Y��Fkt� �x�8�	��4[�O�qw�����j>S1)[ [QW{�*�,u�M���A����ݹك�Pu�~�k���|ab{.b��V�pz:$�;g���2x?�G���H��hѓA/6��xe�&������O�}&�hb&L�ס��+8K�J��ڽ�AǤ/6��ևt9�*�@���p»�q��v��}S�Q�v�bdB�4�{:���*���<�e�B��\�?�:�롇�V��.�ӎ�z�Ԕ�.&@���9���o���h�=QQ�{)�v��-�W4����F�8�#����[���Mۣ��d-����$��b��� 5��U�&|t^�T�j���z�`��t=���S[����0I���ZV�о�o�y���{��:�2�W�]>�+�W�>V�I��P�\��l|�p@j;��ȴ��ؕ��)�v`��+)��q�9��u���sh( քP��:�]��3�} ��s�5p��&�4O�VP��x���ܚ^�C�#}%�QX�!Ď1�D�s5��s�r�9J�m����Vľ����}V���d,�F%��ٺ�Xd�|e�I��i�h�:��;�M�J2��_���璉Bm΁�;���P�g�����wUu��v��iޖ�6�&V���>��b��5��#		�� ^RQ�v�.AM�xX��:s/������9͋�ˁqw�?�텼�:3Y}9d+2,|VQ�e���|gM��M-)E��w���9TD�]�S�E�����R)9��Yjvl��T�]V<"aP	�W`n�Y��|qS���U��jI�4ps�0D�X;�{�0��^��o�Vph���#�c^�S�=�
!u$�0�)m:3�y`)v�����U�n��B��4�!���{AN�cK:�PZ�G(�dp��zve^V�x���k����:LL]�<��["�]=���D���8����.�=������x��'�x�%�t �9H�<�6�={n,>+�'��ZΪ�0��r@�ݒ�$��?�����q�<Y85J��Cc)���J㋛N���æyѶ�d�S�F�m�uZ�|����䧓��騉�V|<�p���g�4ZC����'��T�$���yH<�(O���G��as+Z�:қ�]�G[b�v�_BQ�}��a�/��1� U����X�9��i|���eO3�,5;���L�g'�s�bĊd���~Fh-���n��0�&`�e+�ӻ���-�dl�ʌn��+"�@Nɣ���@A��SksU%A��?�≯�>��x�#�;�e���r�l�֮�E�zm
��)���YH>v�\+���y�n���V���`o�F�E,���,�a��w�3g8d#�l{�������:j�
 �hz/�ؠ��5__���HC
�MpU��w���$�I; �F���7o+<0��v5���.@>�v���4mG��#<A�p�Z+��~	�i7�bW��ʪ���$�j��4�����l����� Ѯ��j���\vk�[�(���,G�A}���⸉�V�n/ѮU������q�g_��-���l!bZ�̯�VA���8�����h�3G���������{�:�쬱�:��5����e���V��,��ܯ�D+��HA��lW�O[&�x���WgK4�aӎE\�a�@^� ��?֧A؜X�������Hzfe\�w�����<�����M_۝��4-^�r���D��w�]�k��DADK�z8kn��������z����b�u`�����`.G$�Y���`�M�f6�����w�/���L$���Sۉ�)�7����A��6~a���u��8_I���e�{	�y��I�\�c�,%�2�e�5W�\������+~vE��<4y��T�L��b6*[�J���B��ҁ�GT!;��r�)���%	A�h:��^i�n)��N�ֆ�^�f�a;)BSfߎ�ɾ� r-YO���L��L���i	4�X�x_�S��>�E��) �毛]����\a/$b���#�Ug�����gU����׎o��t�TQͨ��DG��XO��`��a{�2�h��xuA����ifA/�P��n����s��A�G���񌚵���0�?S����^�g�9!�c����Ry���� C�4����uM��ݸ�[���N,��8��K���ay��?w��h�(���G��FXe�}5k�+��	\��=�Z �&���ej�R�w%q �`c�~˩ ȍ1�HK����}CH�U�gkE�v�;�{
���n8���h��AJ��t	��qynR� MX���v�W�f�}����(Ԩ�wX��7���2���r\"M�a� ���v	K=�"�������k�X|�VtNKk)��V����z������v��h	U^�yKf�dZ�xw�L2z�@��o���� �ᾳ�I ����餏Ȥ{{DV���G<4
ɿ��9��,�K-�R
�]���=�Ȕ��#?���N�xo��̠/�S`�ä/�*���&�P<���1�l�Wc��[���u���h���{���8�+J|�_[��b��GA��h���;A�e�hy�����K���$��bD1n!\����u��'�3H�XjVx��s᧣�A *H�����Fhޟ�nz�^+�7������{���@#�bk,����O*So� �7�%w��4������W �W���<��0��X�]n�Ҝ�gBx� �Y��u����K
J'�CVJ�x#\�jX�uM�K�㬊���/+��>�"Ϋy����6�%�-e��L��שq^o;����m�8�3)���sˠ��8pо7��Z�	 V�2�{`��`�~#Eʏ�Q��;�hg|��^Wt��C1"W��dQ�\�M26!�p7{�X���$�SA����O�N��Qj�h��TZ�hJ>О��|撣�*6�WuN"t���.!)Ws�z�ب�x�o���x��w�1��rb���U�#�OXEd)�?�῎_b����� BʙM;�'A��Tf�;92�3 ��w(e�����53�&��I��vz>KX�*l�3X~i吏���:�?~h�!���oi�����V�X���3�� ����]��ء���I%¬%s����T[�<�e*�;`�A����y��£ �V����Ą�nx��7��2�m~vf�YB;_��H�<!��*X^�=�^�O���%,l#�j��~-�'���������}�jg��p� tS�G�i,n#ϭ�WHy5��q��R�=�i����̀�/����*�g�{��~"z�=��U����[��]��Oy��
�-x�V8���j���#4֟�+�p��о �-�)>�.��a�����E=ھ��`�(��D1���1���zc�8Iـo��s��_���Z��>�@�,���$�R[Ea�T�k�6��K̍r=D��Jz��T>���uI��t��Z]JcS��^�Y�o4c^����E�������Z��U>'�]J�XO�
a�󑚋���fe��~z�<�i���9��'��� }h��ɐ�P��Ո.�A{f$��O>�Kk��DTr8��=���_N+|��)� � Xu���Y��-�;�nu=+
�,&�\���15����������b�ynK���l9V�"4��Ak�%� Z� r.p�>�eݓoQ���̓�u>��'����L�U�EzK�;t7Ͻ�3�o�a�r2� 3��KŞ��R���݊O�Ţ$}J�t0w�*�b��l���ͳ�����{黎Zl~����&i:$��*�K8Gy� ��+��k�N��3����]��J,G*C|8�|������S���M�V�h��T[����*L�,|��m��c����BI�v�P���.�r��2�����
���� �l�ڀ���:u��]�h�\�o0�n��A������BN���E�I�@�&'���%�ܲ��eP�$QO�s��\q��!����l������rD��_�q0��L6�+
�Ȭ@�'�bOB��V�
����&�[�{w�M�s��j��3�V��{���*T��0w��c�%	���8�!������puX��P��)����iҀ�aUy��F"Aߜ)��qd:6��s�"h"j�RZ1^���������U���*���7���8%��4�7l����
��(��#�.Еķ��f�:�Ry�P݋���"S�&:�Г�\�G�e���A;f �Q1�d�:�R��8��Y�a��
��b�>�G&���'I��v�}���W4�y�_�F��
R�Ut{w��W�E�� _��F��)��6mh�v3E=�;�vǇ�mb�ZQ�\�HiP���~�a�kM��"���7J��Q�;��P~�;�^��^ʖ���S�٩|y,2��A��]�D�t�Z)P�=��)`\��z�R=i}���/�O����:c̩�p]'6����y@M=��XT֬���`3�3$0�Ct!�q����]�r�j�,A@5p�� � � L�=K��H؈�((�M�M����{��;�#Y�ڹm97T�S����a1��U�
,P1�遵�ǌ��X,��XCȣwK�����7��^��ك8�%�?o�;�d.ߑ������d�ga�D��Hݯ�^Q�zN�^�� Ԓ隢���,��~v���{1|�ܧ��iX��*�,�(��U�5�w�����L�����t9"ǂ�i���Tk�a�m�ڢ�۬����Fhy�X���%��g2D�Y�a�W���w/q��=|T��%�ڱc��ȿ���ӗ�d!�$x ^� To�<*j��/�Jeu��ev�A5�aw�=�˷�WQ)9�i���і�:��]���1 �B$���Lq����M��b�Q�T�n]�e%f�d��6���|��&e�Z�����"������#��C_q\ÂL�����?���L�5�e�69���>�/^5,Q�v����a�֩���1t�.�&�1�6Y.���g��bS��؋�(�[l�����pJ4�w�+ �a�u���L"Fe]Z+����[�G���'��9<)���Y�XYht��p~�zaLQs*�J����Q��ãb���D%O�Er�'@D���reR����ԛ�h����O����N���-n�p�j�a�;�Oؼ��R� Z 5�2�8�֯�5��V���A�X���ċ��z�Ptn��"+l�L�^�kںP��o��~y�F��V,0.��������������v��
1H��Go���K�0�ݵ���kA�t��<.z�����J�~ۃ�c\�m~�����z�Q�Gn1}�Ό���Y}S�&U4����*��IF�H�GlY֥��IM��Ť'���R:�z�y�����U�zX���"�6{
�t��y��O��$
v��!��l�)�x�!�-�#x��\�\�&�B�"�'J �^�Y� ����ޓg��]�~���>�[�jp���	�*���Z]���$6�J��4��
X�/O�J"Y,����;ў��֛p�Iʶ��ы�}x�b��^��C*z>�&���+ݑE�.�n5����k���fj^���8/%����.�ǧk(o�g���1�'(1K�H��|���t�1/��+߳�Tߊ&c���H������z#�g[�')ooU�o�����]�y0DKnõ~�w�����w>�>�I�N��r����hS�~=n$<��E�P�u��3���[8Ҳ�%���|��G�$�<h�]ke��d��Wa�eו�����Z�SAƵ�/rf��tdM94
U�o�E��4�CN�2�D�@����o��W�������
�R�I�S�г�����\,�|��u����4U�6
�b ��S�t=�y�ڑP0d��GE�Z2�\��aiкf��G��g�"����
�D�>�q�j5f�$K����y�2'��f*<�-����TQ�P�:�E��Ä&���<<gd���e��3����z��ׂ�G�}��h&cx 53-�wf�Y�O!��%�pP;k��hK~�>ʿ�;6%�E"	{*�>z�Kt���p�+Sd�uJ�d�z�F���]%�����aWö)z���m��u�FqIb4�/3�����O�+uk@/�I6�
��F��N&!��s(O%-�`he�ps˹�|Cr��xUK/���{�_7-�|"V����.�E��t�9�H��sx�9�"F�)�����!����7��k���wX�fG�\���ݹr�G:,�ڕ�g��bi�D�i�S��"4���B�r�梌Ao�M�t	:��?c�I��Nf���R8"�{ڠim-B��@w�����R얓���om�*נ��]�E�Z�w�s�C��G�L�Uf �>��-��I}G�*?ra��oo���K�{�3� .���}@&ݞ��4W/h<��_,�x���D��0�Yى��tb_���^��8i��d0]���S´��5�:[,G����w��*�<��y��6�FP����J���Z޶[MvӰP�W1eA?nEީӌy�&��Ԗ~h��ȶCb"��򛋬-;[ƸQ(D�!�ZÒ��w�]�&(�`��!ۃl���s�1�>��G�Bh����F�ݾX
�W=����_埂]�7Q���!�����&�f������S�Tb�$I���$�5�CS�bt���N��P���a�)�'2�`.&��+rO����'UN��"BT�Q�R�ȩ��'����M[J�#؅�KAR�uoz�u�&n4+�D��qzҟ<K_H����*��<4����15�4-��0����ʈ�r�J���αW���ĉ��2�E��M����7����q5o]��m�	Mjb�H��ͪ�-�}w���fs$�5d���Kim��rώ�mZ�Cq�먷�Svj>���#�Y���A�04�:�)���J�������<����Ľ�)ƷB)~�Ƙt��a���Ţ�*�$c��f�BN �F��?r6�J�<��3�'<pI:�{,�z3萁#��|	�/&��͠�`�b��ȉB�G����#�d��ԖQ��H_M�^�}˷��`S���������b�HF�m$�5� {�n��ҿ����
Gl�����;� �t��9�vWaJqj�� ���Z���^r4����+�%���9��Q��.��.H��u,��L�ЌnǨ�3��&���R���Ns}��2����?�YS��$�ہe{c���2�w�kԲM��,����b2�����}��PRXuBp��B�-h��P9�|�0;{�	T���G�s�`�F�h�ҧ[D
���h�Id"�u�t	f2M��D��te�|�*���y���Gʂ�X�)���y7v�J◼��%��Y)f뤔[��T­-P(�>/���Ko�I MrI^zUͳ(�Sdx,G�߼�E��س���+����H���ˈZ%����AD��W��������5}w*��/�C0K+-���SG)�U����J'��W����n��� E&��/���0�J���	��jnUv�%y�����+�[����Zd�n���
����r�!G/B�ѪJ�<zB-��t��:9CU}*T/��9���MƳ���C"e��k?�5�:�|���W�Qt����.�e �V�w��"LVp�ƙ�f���@�*A?�p�F���Y�(���ㅆR�H�O�u����@`te��7kQ�n+2�W�X9���P-� ������*�":����.��i�N�Z5��D��c�D՘QsN�e���T���Q�~���7���\H�-y��7N� �3X������x�_+jq�i[*�G�F81����d3��>�q��kFA�:��>LC�L�ס�f9���oA�Z���g�&����M�S����jYwذ�6�� f�W�h;�3��J03��l��o��H��>5D��1m��Iqj���9Ku�!�G�`��?�e%���C��?�v1�7iJC߻�,t{re�%@�}ux�j]8���	��;%XJ���H^~N��&�%�jP�߸#����Y"��ӳ`7�lu��"B>��]B�����W^i����"�t?��0i����������4�N-0ZZ�J)���K���Sus[�o�]3e�L{�5�w��
mXvL�]1(ǹ�div�g��*O�$�F2<Ȥ�{�~�*x���G�%*��ḧ́�L�f�f�Nq=%z��M(������ߧ�%�����ݤ��9���OH1� �Y��fX�"��Ӕ��t������h5��	v`�`R(�6e�6m[�j`�o�q�PW�54U�׸��y *!B]��� ��`�Ro� �3�RV�tK�_��Ӌ�>���dH	��E%�8�1��/g��ήz��y�QbiW���6�=�NE�a��-H�9N�0�f�Ƀo-�+��YyZ(�45�!��ҕ� ��#\�@����J��m;�g�W���"ڢ[���H��w5pN\$*H�l�D�)T�|����(�,ŀ9�b@�]�-G��b/�� �� ����C�AH�"�\|]#�k�2���:*nu�zxfW<�$��\�g ~�t��/5���į%"�w��	���D�Ƹ]��+�z&q[*�8'�:?�L8�6�-af�Z*����3���b�����֗Fx�Ps�oK��AҲŷfC�eu;�<d��ik�F�{��W���g4c�P��ޓ���]Aɏ����S>辸�D4I�XF�t���#\�6���٨������p����g(Q���H�qE�M�ܢ5�,�D����&*���,�J��J���^39.]��+YHy@��k]�xb�2�,�t!�[��ߕ�AWP�#�~���ζd�A�^J��{>^��+u�e��ߐ~��D�`X��@��X����[z�?��e�hu-:���g�D~��>̏PId��˗}�r�di�L��Ϫ3&�߳B+�rq��֘NF�6eB֡Q�eM�n]tV�s�e�=П1d� $*�4}%��5��A�λJ��~��aGu�+��\������'S�����W�w#���xY�����qT�`p�C�g�9Tdn>�e�b��5jSᡅ��72��ze(����K���={���r���,��_�0��WtM��������P����z��[6,*��Ɨj3#nc�gB'7K��;�T;�mT>�1���|P���C)�X�~��x����[JDT�����*>d�/$��	�*O~"��0�4��\�ʑzO�[���͗���gR6�Z�^�W��kc֋K����O�b@�7���=t{1�-1U if����4z�WC�	w���c���]		������Vؒ[��.��Y}`Sx��qj��X�:��ˏ�s�8���4Gܪ�3q�q-����U|��4���Ɍ�7�R�,g�G�:SO��vx,��܈OKz���>��AUi�K��Ъ&��hn����3M �8��3�#��m?��/���0�ZS�1E�Y���w}�=����3�xr+6�X��H�/��&w�Kn�����L-1^��P,]*����if�P	F��kćĆe5�ç�fϒ��$��3S~��z:i׭�OVQ�e��6p�C�w͟��� ��:u�,������o��������̧��I�^{1D�ށ���V�����_O��ޥ�ȭ;������b٧jn��\�p�1v1�$|�zJ���(Z_k&;�'��cMi�sj�i]��܌pH�f=U�$��J���LkW���z�U�g���b$��j>�Y��Q8�-��"��"�ք,ū"aҹ|pI ��"9E�}ɨ�>�H>>�
��~�SkJ6�AE�O���=�$�-�CPl]��J�Q�k��\��kB�B��xn�D>4��q��H�`�n�R�Bo�������J����}���z[&��@Edu��yŎ���{PN\�K�i����3}�*Ih�I�%Kw �
�܈�b�7B�|��Yh��/
K������.9۲D��y
@g�L)>��0@���R��ꯀ
�@�4��8�.����; ���L���҅f���������m�eiߵ�Wh�A7|�V�~�2(T7�1%�4�Чu��������"lu�.ff�L�[~p46/.׷�&��T������(9�e5@�%�ۛ���	�����Ҭ�����(�+�ʶ^�)��栁���m�����H^�4�.���5(#��f_�3��Q,���OD�CN��1�e����G�YN��R(�.J�?S%R7���f*�owpI��'��� Ye}.B�u�o��n��HR0�n����ɓ��J�H%,�^�2�{o��p�m2��X�<��Carb�4E
������=L�W! >go�[�w���1�;'C�?�EŶ�
��}
.%>�c'�лq�a_�w�&Q�%�l�C��E��M��"���GG	z�Z���z�/���n*�(����'yv�s����8٨�ʌ�����M;oW&W\���$I��lTyd�6R��s�,���o�K���\��L/�0�W|�D����o�Y����)��!1�%Jq��Y�������|.�4���epsm
7���[>>��l8!�࣯��ل"K�t��JC�>+���G�>AV��H�R�C��kw�Ӣ��#�H�ڂ�ϧ��I�k����.xFM���:r�L��D���p�����;����B/z�6��ô��d5�CoK�쒦vp�y��YO!�˦��ZϷT)O�»��ǰ�?�l�u�sY�`�fE�\q&"]Tow��6���,��e/���!���3�����㑛�`�^٣֪mOD�����7b��l�|�8��Hg+�h��yBy+^<Tk���0��V7<l[.���3�{6h������pĲH#T��NO̿�IHt��%_qw�^(h�$���b������t�zX�����ڀ=�Q��8�֠�������D^���#��ӃN���CX�����FNe�J��q"�&H��\��z�ظۻ��l�ؘ�m�i�t����ʟU'��?��!����u�y����'��V�buC/�� ս��*�%<7�,{�-V ��mn���ï�ɀ-�\9\�����.��W��X3�1C4P�P�N:�Uw3�08�] �d��{�*���1RL���{w����?�y�X���N��	����2b^�ގ�ƌq]i�e�x��>���0���9��̟�=w�K�إ�#5,��M�����3;����*#�g:E�"��ʫ�� �?��λc���[A�B�#�:I��/ulH�BS/cw�-rϭw�h\�Y���yEҊ��t���sѴr]�յ��K�(^fS�G�G|]C,Q��;?�������־��q^g��5izKB���O�j�����XI��Zo|
�s�yǎGqV��A��Xo<�b]3�Z�O�Q�B���Eԛ+r}��-Ao�2n��[�`@U�e	�������C�xe�I���#���' <���K���íP��x����gd��=���9�1
lUJֽ�m�W5��oAO��L�Ei�����.L�r�<���0���mAi��>�
�`d�X}5��=�qߖ{��Wr�Z7&��6Vr���.F�� �O~ )������ē�rߘ�$'���q2H߇J�<C�SHU3Ĝ��t�T��j�c�22�@�)�dj?Q0��D�E����p���S@�#8%v��=G%ߦN�4�;Ċ��H��^��
�n",�?B>XoJ���p{\VΊ*����ۋ{�x/���u\�kQke'��=�M`�7A)wC�C�O��6M���כTTZ��^f�tjXU����F��-��Z�>(Ƌ�+Z����k<�@��Ő���96�h�Z�'��-���y�/�,��%"�6�T 0#�xE[�]x�VޟL����Ah��4d���fȽ9d
/��lUٻF~��z�_V�)��itf�6}w�.����:�L賲�`O�M���W��e"Ţ�/�ҵn��`9�=[�	 y ?�*d�؅�,�Z�@a��_�B�ɶ��D�b���&A7�,���˖̀�,�e�D�F��~��5ƀD�8��/m�HD�xb����"lۭ:M?�94{Oip������)O�)�HBT�Ubf�=3�X r7�a��0��5��ź��Θ��nM���.Z��3��><�؝�1vk�����0�ܐ	#������ĝ�k;��U���L&�H0�Tg��]�3�� �9,�3�&E����N�������J�ԙA��1&��P�S�Xa��/��~:��F#J*�cGTd�f8�z%J��^��#&4��Z�K汣;�\�Iov�p�K���.��(��z���x{u
O�Q�Ӷ]�?��� ���n���߻������A'�l�ϸB%��#K�c���(a��H���bK&X�Q�}�!�Z0�3l���0���g���^�vhd�;@:��n�[}���� F�t�0BB�_U����d��2P6NʐQ�*�Ѣ������@� �+���B|�[R��1��J^GC����Ȁ5��R}��Й��$]W
"���S;r&�uPY�����. ޢ��dy��=�̽���>Yּ�t�w0B��6�7OXh{�?����c+��Mw4��/?��?��bFЌI���p�8
��[�
D�u��*��݈�������i��/>k�a�'��.f����8��p��a`����X�|�#%��94ָ`��E`c�r��8-K�H���J�{Ō�<\�J�/î�� T`�JmP T@ 9�zxu0��o5�A�@؞��5��nk�Ǥ3��w1���iH �#s�?F����jkA�g8H����c����ۭ�6��)Ī�i�+����i�!)�7��m���'����]�ށ/�|�M`�!�����~N��L1��/���#��ر�Uǡ)�''cE�Hܗ���B���֢��i�ln���~zG|} ���]\t�򀝢8o��z:�
�A-xwvA�fnMh�Z���h�N@^���g\�ٕ(��Er'��
�ו�+�����[�C�G8�N��Z��b����P�;��C���H����ɬ�5����y�����f9�a�����g��d��	,L��e�/���x5���s�+�Ʌ� �1Џ�D[9
_3٥A8�ָ,[AdveowR��,|(b��� X���o�[T~�)kTUd�2��h������=gQ)(>m%�q����ͺH@4�!����
A������r����1�x�����x�b�L*�G.�`�i�
�!�s�����w���?;5c8�l�q�lV�Y������y�3(���JR�`��\�|�쌄9���c��B[RF�[_��NL:[;�}�zȐ�KU����֜��#S�(�]��~\t��w�m��j"���,�����M"����7�os�Aɨ`���LTV��S�����הIG�舵�n��)����
`�"'ٴ	+r?���*[D�W��9PJ�\]3V��4L�<�M$������?ouE�Yn��_pc�=.�9����;s&�,!���][Fj�u���5G	#��.'
�+v^�	�GR¢��mU�Ja�?�b��&xy"��^A3E�%�?�O|��+Sgo��Җs��tQR��H#�ȵa��8֏�R�y�#)+��!���p���]^Tc:J`8���F���a�(/R��L��O�E��$�/}XVZq�j0��RT�?!ױ���n~��Fi�1P��x�#4k�^Tz|?+�_3�1eF�kt�I�\*�^�)����*��j0P�yխ*I@2���$�1�f.�!<�n����.�b��͐&�	���+J��QaVnE�	,�Ɗg�Ċ��qc�!�U0��>t5ox���u������}��L�J8+���da�σ�}�$�̚��+��wsj@@�]2>	�+�s9�+�� ����hV���&�6���H�_hʖ�LW�x�!��Qj������䅫0�,�`Yg�.�e�#����xϺ65����!����Q+{[[B��3�������cJ����=<l��c�g8%_u�:� ���&������Jq�ᲂRq�J<P׉ڳ#;I�
]��=vcE/����?���ń>V�20.����h�͕d\��|��$�˻)���A�s~c�r!���7�a�~�[E֘�(KTS������JW��j���T�G��A�n�һQ��x���|_ʔ�PX)��W9����H�w��"���({�����X�aDxb3lE����	�<���7;�x���x	̼�
d�0����U��D.�H�� ����˞���3�*������ʅ�6LG}"�"�dV�_ͤϙ
�B�o��[���Y��%���+E7u�Y+�=�/�:��E$O��[9�Q�o�:��ɞ�b�Z���Ɵk�2��${8��r�
<��0��S���\���`<vN��-�r�gF~��r�P%�=9ښ���h��؍���y�����E�y�i�U	�|������WPU|O�x��SQ&j��K��Î$SWX����>{w��g��@ըa�`#�r�f/�E�����=Ul	���4!#@�b\G��<mt��+��v_f���En+�i�Uyv�oX,e�3u���H���b�w�x�����>�J����P?Hϓ�zҙ���֛��3����Ud��AZ���%E��Ŝ��. �����Z����j(�I:��4��o�5#m;�995�Q�R��IAt��VMQ�}�wJ� ���a��n�dֹ�3�O7��u@��4]�s�x�HAc� h�kL�܆�DɔH��$����<Cr�TB>;FѣjRIKa��wt%��������G�yH�o�9G4��JӪs�d�:�7.� dZ��T�#L�"j�6���*�a"����_�W�l��ɣ�@��Sѻ�4Ӕ'���+ 86@
ԫ �?��GY�B��_�^��o���8�	ܹ�U|ɇ���:���X/��9��"����}e@Oڇ���6B��CO��sZ�L�����^�=�"Dk,�(}@� �Ռ�����C�u2�P%�7 ��}ޠ,8�F���T�aЛ�<,�Ϋ��z6G���+�2�@� �?v�+��&B�=�MV��n��5��Kn�7ZTZ�d^����?`�c����Q�b$���a��	�eD��݌�~�Z� Z�+\����K�'V�	�Xr�/�����$�F�_'�~n��,��?�{t����J9��=���8��&�/�)�୍+�K�Cã�dn�x�n�=d��Em����ᒒf?/�=��?@e�G���i��T?)��	[LM��eu�^���ֽ*w{���db��|AP�7�� mP�����:�D��)xu��D�U�|����\���!��1|Y��3���Ť��,"	����`VD�	�T��W��l���Jd���I�`	��h�/u����/ lXm�2��~���5��TE������o�E�V_>Ia�9q�Y���b��qB3��'s��靬�5�{ ���}�z��<����׍��L���煜̦��!8���g�/�%s�,�'S<��)��I�*k��/�� �?�h�V�:��ME�"6R8R>�[j�N��*�LW&w()5SN�V��G�����E�l�S!�S�{`"<����i,oaO�F�%ce8�!שxj�wz��u͸lܷ��I��$�X�o>�8�oe�|�j��t�d��*/����+�h�f��Y��N��tc��<bZz����?g��%���7P���s&�O:Gtj[�O;M�5rU���1����M���*ڄ�� 8�Uw���=G���K��IOCv��K��F�/�]aQ��,#i���x!n}�y~1B>ih��7�(� 9�D{���xSb��֣�����|#";����[��n{�}5wTaT�ɮb����u�6ɴ����j�#�@D�dy^�����v|v'�j?մR��![a��p�֤�\���F�Ax�Ef]�#YZM�Z��u�0Y�=���q�̝�!=�Y��%��0k���Ng*(?�R��^�L�c�
��v���O��b��>7�<�㟉8�yprO��ԉ�y�A�@3�R��y��4�x�Ч���ٌۨ���p9�	��pR�*�\�F<9Kq������m��3%6� ���E=��K�0��S��8*�a���l RlIvޗ;:�0N�njǸ�F�;�5(�V���I,/�UyD����I���W��伸�r�i�±����a"_�\��U^d@0߹ *	3v�#��5Ll,s�N�EPh~��Y���*�yw j�5��X*b�ֳsE�L�$@��h*Al]�(��"s<N5��K ��Z&��u��_�w�	5���荺���p\KJ�q�zA7���y����3���kU �.R����� !�6ǣxTUyY��-� �!�N*Fk������珧F�h�AW�1[���*3h˺����;�jhR���'��̘�i%���ϻ$}yN󆆵6o���ډS,���$j�  fi4sb����*�C�������6�N���q�+7w9��]�r�ٻ!WZ��ۼ�SM.d(��B�6-��&e�m�9�%Mj5x���1�J���9�'�ށ;���)����m
�~�2S4��}��L�K;|wQ��2�>��U�g�G�S,�{8H��[�2~�R8H C�|�uR�@jV�u�-<��g.9�\���;���ђ�Um<�t�'ULU�Y�$�����W7�/�ʨM�� ������@�ZԠ���+�A�\�VN.\�ĬB�e^��d#��4m8n�XCO7l7�/R�oD��u;A4��,�����w	��j}OT� �-w���Ŵ�Q�1�e��,��8�:j�������CQ#�Y��]�t/���l`p�Z�a�aR��EzĎ�;FY�K<�ĩ�	ŴYQ H d-X' �32�I���//݄чF�3�:g��f(\�?Yl�{�LY��U�g��M�����
�^mܻ<
��{��ov�t���ü����d	�K�f��M���{ �3f��}�+�A��	os�-:� �\��0�њ�-"Ԋ|�_��֋�Ǩ���7�����u�U���4���
0��T�>x ��1Ǒ_LP�� �����_���9�,G6U�����꧶pXU�(������^�W)sƔM�LS:%��r�g(��9c7Ǩ�.�"��/L�� �M�G�M�q�XKBF�ף+����jn�SUg6�D�a��ԅ҃���_�ƾ�z���s�m�͑�r鞝eT���/�z�ӗ�i��a)ɦ��B�J[�}�� rGP��#�dr
H�	�L�OX�&ڍP�×�q��o���\r��䕉KPVo�'3Se���xh>�����l�4M��3��9y�,�'��dGkPd�+�CTZoc6�H�\��=��i�A8�y�'(��5����kd!+wO�AOV�P�Us��K�Xcw�=r*OvBU<�%yGO�������+���-���F�M8I�]����.��������5��6�Ŵ���,n��=�(�t�g��MO�ܠ��@OF�>h�&^�;�\NU��}���
�d8�3�f��V���4Ɨ��'|Y]������$QTl��(�.��J�:�h�(X�\���ﮗh-��#�d�+?�Ȭ�b)_�I��X���K�6��B��ȅv�����h���{q9�5�;o�򕆦��+3�������A?�?ͤ�\3(�>��X�h��C|wR�/6�����M� ����z?���q�$w�h��D��|Ik� �\��B�TLf?�1y�-��:�T��e��\�bIV�26��}�hQ�cZ�g]*n��5 JdC5��[�k�,�^��g�W�Ca��w��c/#m*��łMR ˰?.���C	���̲��v r���@p��;0����������.oY����YMD�y�M*7�ѧ�\y����?�g�	S�i���kv�����,}�������y��87��ɇwHVa���#l9�Q��)��i>ע���:�z�A��V�ɲ�RvR�h3�Yb"bԄ��5+���Լn}C�OF�زy`��N��w���K��9F�(�i6�|9�L?"��!��ox]r��V͕j��+ ���D��֨/~�<4*���:����q��JBT]���UX���9g�[OV~�^��
���}��F�WR|�5@.�gDR����#��فZ o���b���:V�&�Ѯ�敡�eT��Y� ]����W7���#ƸtQȴ���x�c5Ѵ���Ԕ�`�9?�F�RQ�����>G����K�@�d