��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P��v�"<ߞ��&'��k%P碶�R�ӣ�sĞ������FY&��["3�l��-�n�t:�NP��Y������2��Y�FMv�9(^5��6�kӚ����6��G��A0��85&{�[�$�J�?�Z�7�ԡ=5����=�Yh��#��g�C�{�TB�ͲEl�Q�ŧ�m1��%4�<+8������&7[�ɱ���Y�&���k[�05{���ih��(D�+���2����c���
[�.bg�ķu,�e���C�w��S���4�Kd�L��<9F�9+i�A3��� U6Whj�N�A�8��X�@��-��,X���(v�>�X�K���<�J�6���Jɸ���|�}U���&��/W
��f�Rm�'�(���\������iц�vӝv{b�s�<f����Rd�K��ۖS��+�wd��Ĭ���m����-��D>.
�f?��CX�drr�-�i�Vc����NO9�9O�70_�,K�m����Y8�Ӥ�m[Bh�e��/l��c��!�v���^`�}1Ҡ���ZB/��5����ί�s�#�����$�&�����F�.��8,$�9��Ɵ�ɨD�aT�	J*څv����ngN(쭝7oE�_h��>c�yg���UN$%]�@1��u܊Ֆ�0��v���C*�G�.Y��O��^Ɉh9�P��[{G�� ��E֙$)�YA"ui�ӡ��D�_eB1�{y�������U��-����I2
�\5�{7���&2�|��.��&�O�4�li����s�x���n�#�5�2p?W��1��c��_<
[Zy����@6}bV�K���95��;"f���֪0$�S2h����u��0�IQ��*5��@��c�N��;5/S�s6�6�3��̣|��I�z��Q��+��D���Ӿ@�K�5eM���S���������_�8�l�S��(�O�Ђ�����6�g[ �I
�bS(� �%MD�p_�-��4�ѐNA2�E+K9k����g�,�&��S����1��n��[J���C�ɇ{�����A�ب�(%���TV�
c䋈�N����? ���nhD4�:N�p� ���(J�R�D:.���
f���1P��@�Ux{>8L�Kc�`]�|-������2xt8RSĀ]^
'7�����C*E�E�y��X��/�%Z��\..����G�����~�ȣV�P�8��̢�X��ń~�Q >3�~p�^Yi�:��&�Dw����	�,�>�ڲ�|h�l���w���BЈ�5��������	�&OD�����'���bC/���u=Ѵ�LѰX�jpi������.�^��#�@�1�u���@��2��7�r��]��e�=7d��Nqai����hv��(O� �zZ�!��JI����K�f*�o�wܧ��?T7�%��9`r/'H�\,�@�F� `t��v?𰷉s���פ��[zG��{#���*�}t�sZUOB�� �Z�.[ڭZCF�Y��M��]
��0�<gdW�=I8�������w�:9��¸$�ԙ�L���'t ��6�}�n0�v�zc�T�����(O����lҸ�lF��A.���]/IŖY�C�5m�W����}0[��D����W�x����=b��$n��4�2*�'����0��R��.%)vIq�)���a_����[�IM�Ux�p�c� ��1_�|<'u;C/*�C�~B�C("�V���/r9��)���X�h
������=��Ѡ��<.�������e��:����7��ZD�}����!ӊ���&RN �!K�9���ګ��V�s����Bٌ��@%���Nݽ����+|����;C/tM0Xܳ��L��h> �TaJ@oGi�h� I�c����1�j�X��Z�(BW���~�����[�
I1/������i��j�'ق[�2�pm^[r����J?�AE�+�"��/
�W���j�EnN�owXV�d�p��b��<�@f�q�T����S�}�S�:�jQ���M���FZ����v�D:�2%�`� ˲�6�h�sg�hU<"|���l�r�W�UT��c�����F�~{rU��[��-��WJ��"����JIt8p�
}"�>]�g�i��^�b}�8P�KO���gZ_;��a�dScQ��M%L%�o�Uz[��l\��`P���݊�"��]G���A��Imz�1�l�$A>���V7�	���MG�"6vY���8�@����X��[n�w������Í�S��n�&nu�7�����X���m_���!]ˣL��ڞ�@��ZP�ܲ�.�'
Vd���L9���!0�TW��8�,6� ����>\���E���k��m*0 �o��J�.�����BNM�����rRux�F훹9���__rL_A�˻���H��*��FY� `�t��u�~S�H��4�V���uMKiy�F��(/���5%i���#�?d��v�!]4�C�j�t���|�Z�2��N�u������p5b���8�/��Y ¹�8ÆE� ΋)����>�� U6�;[�4&��y���ٳ���)!.��O�k���4��rc�P��[M�F���Fya�)r�(��l���I5TSsQ���X�� ',؍�k��s����������m
��q����<3*��4�#�j?��f�F�]�I����j+׶�l\��bA���9`b�=M����+lB*��n��(Nܻ��+;�{�G��>�V��l�-ʸٷ�R�Z��a
��f��.䤽�w�`����~�"i�*�����^G�xzh�����I�.m�8�f1n���3�Uݗ�I� ���	~\��������v�)�^?Y�z��5����jgֿP>�2:�$��#�d�������a=�"8J�� ���IE%�i'g1w%֐��9@�}���%�f����ۗ�}W0:B���yV��e��dn}łs�U[��Ϊ��&��f�����*Zo�gSٓ�������w2�օV���cv������+ɍ�����B|��.CS���7��O$Wh��/�P��N�VȎ`�Ζ˿��UZB���3�]�Ws�U�[8�g���c*�G�=�+�Z(OX���;� �T�[~e��q �%�_��_��$����3�{��������6Vs������p���+�)�8P�lC��=�S#
4���yB���6��I�a���	)鬜hע�\L��9����]t���u9��I��"�x�b>�Y⫂�I9�/y�R�/��ɝ����s�V�C=$rx��$�$���������'�e*2��069Jfh��=:�Ɔ�����yJbZ9=p=��qCu��=�It�~���غk��I$�z����%�c.!6p�of .JV���՚?n?ſ�^(`h��&�@)��9t��{iM?�o��#I��XE��2c��w
{����w(�ӹ��޶����b��z��2�VK��r���1�z?ן��fȠ�f��P�������.��ƫZ�O���Ae=�b�Es ��闝4�2w�����)�u*��i����DK&n��5Z���]s.jM/> ���-�og����$�������C���~`�C����&�8��Fȕ��ɟ�*f*�F��客��w/h|�׻6s�"���5:U'B�ohA���ڳ��a��$@���שqV�،��Z�U�����:Y��Jk@�2rk�í���R^��~Q#���ۻ�HR�+(U��w849lƳ^�� �3�ک��{{b���(��I�]�����6cY��&��;�5���r+�}���Vl�E���F4�֐](ey1i������^z��ؐj6܄��f;���w}G��h�:0ɀ��aw�ٿ>u��v�a߀y��{ČcZf�"4DA6n�!�a`��d/�˻/ᓐ�9'�~EcTni�A�F��"<ͨ���D!2���B�PХ|9�I��*�9mY5����u	�c[� 4�S1E�_{�;�x��T����\�dy�_�$&����ߋ�;�2����r遛쌩�,���!y�b�^�H�ĂA__�i=z���T�ud;v[,%x8VK��y�g���Kо	z�����Ybܰ��w���{��Q�2����}��4I�x�B�Y߼�
�d���c��4��!�\R���$�,����')�k"+`�jc�b`'���6��n�у�"RO�Y�>�I��w��#u֯�sĥPA��9};���a��Ys����H�k���G
_�L�����;���Oe�rc)o]\��Xc�ޏJ�ڃ���ҭ�F<?\��_�q��&�Lk� +�C��*�e,�;lV=Dt�ʴ~w�o�P��ޟ�3�^lnw8�y\r���cQ��$5B�������~���0�4MB�i4wތ8���J�3H���1�Wt�2g-R�$!��u�X�AY8�����Lxe��qB����Og�Tn��;|L&*�.ʠ�~.h�Gn|+{$`�6H��6��p�R{��ߚ�0���e�)�̳�~^��}i�g]R�{�J���2aB�X�^�����8�d77�͖����Tq�"�ڑ��n�
xx��CEp��R�o��M�ӿ�P
�K��NA�j�L`�녘�W���SJ[��ɲA�V���ov2��ù�`J�.���BR���;qО[4 �
��ze�v�x���)}�2�4���#��Q�n����E8pгUI���w����!q(��p�4c����l�@?[{�LþsE|tuI.+,��o��Hҍ��Z����V �]<0����Pn���[��^ʶ�m���H�yVh�:vB����>�b�޹rs\�:��I7�)�JU���z�]ˣ`�2A�@B=89̄�����m+m��f3�UA8-$����
�E
�bMX���.�b�2-X�:�F�tSYN�R�{\j�SE�9H�u�0k1P��w[��Aެ���X:������k�Y<:��i��^� ������<���i|�W�XAfn���Z��>s4M�H׾���h���&��ӗ�����yx�w�"y��)�p��:k^GG��Ly0m��9��~33$��nr��w=���j�E�G�ri&l��4��R��"@� r��>�X���iF)�&�|�&��'�~%@Frn��$�x��n���(����Xmhɦ_<��ş�*���(Ea	��X�䀉��<>��<��B�`���;ZQA�ؠgd����𡏶A�,L���Ay�D�%�HNǗV�-� Kh̎�.��Wh�� ��j�f(�����Ѝ���'�8���}���g���{l*��.X��g���-�{r}�Q��f�_���=@.׼��!��B�_��W�p�~����d�*���ߥ�S�ˣ�����h�;���N��.�	�Y��m���Й�'P�]��z7�`㧠��*+��?��(s������#�YZ�g�A�\Z��Q�(ͽD����RJ����M."�^�z�gf�gQ�3 	G�j�����hܢ��N�	�_9�¿��l��	w���ʧTۿ���e�9��X:�U�V��b�i+>?�e:g���!l�V��N9�B���I�i���@�%y����;���]������zd����%-���O��M��k/�����딅�D*)�I-�=0�!)�,��K����h|���rx�ES[��-,�-��'5g!�WQ�D�#�x�c�� �k��A��Ra��WKX��Lw`���hj�ȼb'-`��7�H��nO���0 #|�B��t"�D��/���V~�lhC���/Xv��t4������5QЅ�z�6�2�٨(a�Q=Y5��$���_��M�p$H��݆\��Ӊ�e�7ˬ������_�����CXTpE�8/�d���8��*j�	/��h�k`Ģ�����"��I���s���6����.����E�9O��tW�|�R����I��cz�/n0�2�D�'��6L�0t��{½�Y�7�ݴ��^َ)�		��̞`7?ì�8�mS�w/�i����ƛp`ʩB����k"Y�7��������t��G��Bd|��ǐLF��\�� n�-��z����E�����]&�@&��.�oo5�y�*�l63�G��P�B�Hc�/x�1+����K08�k�{�f
���5Y��"�.^Q���z�@Ǚ��)�6Yo���c&H��t}�-����Ǳ���N�nP6^\����],��DjY@�䨖�ƃ�~�����5�@�A�4h7�����1\���Ti��82������c 3J��H�� ؟��ȃ��n�ψH�IN4���EN��ng]hd��1���oSǛ˗�A	�X\v��1/mj�#�m7u�.ˏ��b� �a,Y*f�E��c.�>���3k0.�=��)��*�bl���Z>R24��v�1�9����S��UM��Q�}C���w1�b�x/�=��r��h��%�a����*~S����t��&���R����{r[L��H�*K�2��`U�����8e�~:�Љ��"�I)�ei�TWKH�1����l��ī�A��@@7^1*�v��<��/��A�����+9%�^�jj,k�����WPNƁ�\��Il'-��t�p���`�$'�n����1:����[AF(���A0�9Xt̮4� EϞ�ӿ�!��u�l��X�����^D�w��L�8�t��S7�߶�������Ԑ�P�����-�X�T�>�݊T-5�B�p;�P�`�kq|�L�.��9�����X���J�J�g�}t%�S�S�w��6^�t���N��TЙ7{��,r�U�ė)�E��Іo
ܭ�D�+�T��J����}H`�(�'s��Ye��pj�	�%�$1X9"�p����%�ϔ��c�2����N�,����s�8D�{)��Ƀ�{"[T,�8���V�#Aq�cD��ȯ�`��;�^oQJ$(�A�C@	"��k;M�A��t�z�2L��/���@bo?�C-O�����s$J<I<�k5�$�Y/��׀N��#�~s��Rx�)~�loN�A �ŀ
��u���\�$��X��t�$D'v���J:���[��`��,���u���鳫��¸���n�+�NM�K1e9ڡ;}����;�Q������6̭@~��!�D�T7�O�8�Խ�T0�����Y^�wI ����{�H�f</k��,��~x�dNG$�㒨��L�ѹｲ�>l~ 㪚D&�+�7_���1u�+M�e��[qF�	c�kJ���9�������қ&��j<��ߒK�ow�|��a���J�����鷙�\�kXY�f���ҴR��4��������׌+@R�E�+�,}�)�]wGtk���;J��'?�Rˤ��zi����>�S���W�A�O�EdS��d$`�ӰD���b���Ro�o�~��a��Osypl ��ڶUM�����t_ ��<P�D?�t�vIr����t�G��B��捵.8�_��F����ˏ���8\.�/"m����+�r~�_�j�����`D�I�'[��ˆl֖6��0ǋ	Nm9�g���%�򹲄s6� ����|���ɵ����}?��|�b�f4it�T?vK�
I���v1;NJ��O,�~�/�l ��2w�<�ퟶ6$�S�!"���F%8P��~"�۶aA/��ә�JR�\B]�F}S&}ͣx�]4�)��,��w!�H3��I�/��0+K�v$=��N�Om���i�=��`A���c���r��� �H�n ��z�OF�_���b#�3hTO���ӵ~���rT��8I�I�+� ��(ry%���.�� �+{��|�uJc�3	H��؊U�5!��ۆ[��xB*�/[�2~4p����q�f�t0}l2�}������ۖ����s-�DEː�5Q�|C�s�i��PEШ �`�	ri��k�E�z��`�P,�p.�.�ǚh�[��Eڤ����{����'z�鼢�Y���z��b�=�a��a�Y01����^~�s������]�t2x��~��H�����)�[5��P�Χ��0�J:����2{�E���\�Gi�R�y׆����.���:u���P�`�L���c�E�?�U�T�d�w�U�	d�%^cF
�>b_$1(��g>�-���&��J�+߃D����| ������.���z_L"3}4��/qԂ�x�x*P�l@��s`�nt�>Ftb�D�@a���y&y!�<a� �����X>1Bn��q�^ ��)�ў�7ݕ�"��q �N��M��lW����ZV�1p�<�v�GͼO�x��>�t!鴦�-���Y������P�V��W�_�#�����:9�P-��8�<��%S�g�M�2��ƘE=;$B�������E�81��Z�i���b�D�^���!��A�#��hr$�b��/�J0 [H��q�nR4ii��Ӊ�t� 5��'���!["��'%�: ��z�}�s�+;��B�7�ֲ�7�p�������z�������^.�6�2�/�ûcF*������Ȓ ��k�H�AE���T�A�H2�T*�nO���Ϩ��3}@��bV����9�<s�X<uYk�k*ӖK�qy	}�eZ���5���;QD�ޡ���T:��=��'�!돤t| �p ��=�D{���X��h3ɝVj�ZLҀ|��������%Լe��WP��Jދr(c�"��U¿�Я-�Q�-�s{�1��i1�V��[�p�K�8Fw��@����M�yD.X�Pp����o8�@԰��%:�Ar;����ҿaqtʊB��L���bx�oy�(
��fTh�m��l]K�[�������FTЧ>��},��3Djԡ�M%B��>��͏>po��D3,"`�h8��u~�es�d��I��z �ZL�`� ��%31��51k�_$��FNg�B3e���g=|@��֘a-e�I#���ρ�W���E�<� ��,}�9�e�t׉���؋�n	^��Y����C�Kp��n7� l��u�c%˛2��.��L��Pi��J�ǡ'�*S1ʬ�������7K��|���t���<�@�����ڟw��$�]VY� BE��Qyֳ�o:F��u6^�=��ڳf\����?d>+�\[�أH�1uj?�؍	W}���)r@�7O�wW��F&������T�~�P�>�d��Ǔ�;��"|��7:Z�n�Qc��J����HU(� ��Dj�U�C�dTӽ��3�S�֨c+pɥ��v��U���~�����6].����W�1�S���1	�V�9�+?�8~�N���f��G37�o���l�GŐ�J����cSsܥ(�Зn-W����H��1xw��ԪG�����`��A�;
Q,�Q��Z��m>�I6�� dZ�����������ٹ�^��jV�q��Y��"%\��h��Z�v��P*\϶��1��=��ṜCͽ�-��%?��  �� �oyܗ�$�RY2�qn����Ҁ���<����{Pi��9%��N�}8�-]Ӣl9n7�{��X}0�=5%m�O+��S"\�x�(E.��\���h��Ps&hT�r1�y��1<&O���P0^�`�,�LX��$#B''i�Y��\�<�0�%7�����^-pQ�ω�����-�o�Ky���$>h�fp��ji��X�~j�n�]�X�IS�#w��5S�C�}���I�T�&*cwOA�8|������ߐ�ŴG\���떑�6ToH��9�a5{$��gI�!�݄��J3��m� �[/��1�������iz��L��e"��5g���{�v����Ŭ&A����\���NX������"���E�f�c��l!M$U����6UO�%�+�����I��KqSQvg��H��=���痥Q���-�N\���V�k �R�F���7m4OP�6�x*TM��:��Iz!��0Dp�ccQڦ9V�aވ"�8��ao����{���㙑���F�����/�XCT�&����&�u�G{��nP Y��ø�Q��__nA�҆ X�I��iy���UQ<M��~�A#v�,���
���5ح�}T�V����ï�G�Z8ǀ�R�aC�I�F���4\J��cy��!��TX����F���~��ZK4o*��([ŗb�CA�H2�8���I����͔� ���ğV �`��أ^Vҳw8�.Z�[:Z�-�ޔ�����w��AV@����Ln��j��j�qG�#P~eK�w��|�RR�˅W�4U�wk���F�h����	��V���՘���_����s��,#@u(�U��ا_�{/�s��C�FF ������9��C��H'��0Y��+�#E�����#�a���44�8T̰�|2�3��_b���\�_a��---S��GX*��`���l��>��c�-�E�l��k�'�Op�2�Ѵ�����rh߭]CU�h�萑K]����ca��<)�8��Ia�/>�Ǥ����03g�����3�ZL��>�R�ʚ�{P�MX�:�f�̋D�'�1m�"R�
C3=��{��s9�H���V4z7 4.�u��5�g��5�J)�,�O*���='f��/�b�����9:�j%3s���_��M�-���u+�>�� @�MN����Va �LV/��B ڟ0�zI[��H^qՊ+"4Y# �g�둘7Ƕ$��d��"t�%3�r(����/mVO���Z��|��c�W���_�k=�1�7_�U�<�W��J�{���8����IIi�5��F��#/����H��Vԟ8��
���� ��
�6�j����sF�q�4�u�I�}
����;P�
���v ��Cĭ��Y��<��j����ǩ	ˋ�(���5״��O��Ӑ�O�c�@E��ht�x6����(Vr���� {�	�
��~ii�v��������NG���X}9���2)O�SE?I{9���
A �-J�z^��\�ڿ��5;E�v�<T(�#���b"ԒZ���U��d��g��W�����C&J]���,��zC�I��J�4�7^�c�
���1߷f�>��d"0IB鬜)3#Jˆ��>�p���>�k�W5۴WR�;l�Gt;ۆ�����p�쯧r�� �c������$ig����`��ҴI���j���'��	z�Q��SsAĒvK� ������y��R��J�v��4������z��Q	'��1���B�A���	�53�����h�F�q�4����̅�-r��&Gb��iOxӢ�v6�d�Wv2d���F���+ŀ�:IjV4�ׅ��>0�`<�`��XD��w$ߜ��v�_�>�;�Q���gN�2YM�P̓�y�w;����\I�l�e�Z���^��'b9��O�#w�c�E�q�xsJٗ���l���<��ѳU�ډ�G\�Gt	������s��v�nGM9.�SpKdq;������o��1PORèJZ540h'*#_�����×]���i�*=/�����ec[����؝��wJ�桱��z6�}�����_\ߒ�eK�HD��Il�%������1��lk���	�B��Y��'���&-56e�\�R7�_јJ4��D�L5�&��U�����|2�Yv�z�a2I�ؼLS"�k��$L>
�l?(.%=��3�	~�	�gj�*��G���?lX_\��_����|�Ƨ��Н��ӏ1����S�2�i�|��������3.f�k\�/,v�莀5���dYU�o'��ϦC1��K��&M@��?��D����꺱`i_v�o��
dн�����`�{��\9������k"�h�^�@��Kק6���+K@��,�F�6l�|��4�����A��q=�$L��1�$��&�d��X��Zj�A/H���
'F1C�7_�x���ixh\�e�A��OTXc:bc@�`�z?��R�_��A�`��6#����b�jgu�������	 ����=q�P$�yAϺ�4�y]|)��>�l�;��:.ԓ�p�sᠤ����ߗ�Y���*�ݰҲ���odu��d,\Ω*nӓrER%��ߒr���6Eݶ�z�"�E�*�����Fe#��l�`�i㄁�}`t���	�o:q�I���{�R�a�Ǽ�>\�Ӵßd����j����7u��sQ�Yvn��g�" {���!����ݰ���K�QDN�V d��C_1L+C�������P*�-`GD��5G��"����qy/�F4%L'"$h�Ԉ6��EX���o��� �8��xs�L����{��8g���[�������?����F�����^����������e��u���'S�$����d��$�G�;6�;�(3���y����O*�"<�uSD�UҾ"s�+p�ȓ���O�&֠�g`���=#5�n| �Tk�V��P$�I�fK���2e��Ӡ��*������oj&�R�ˤ&E�H2|�P
�S���10�yn��HA��	���E���$\K�5�s$T�Ԅ�o.���y��eG��C��$������N
´�e��9]=�T�b���b�9�Hw�h�?1D�:�&pxS��`�_�fPWw��˫�D>=�8T�#y�������ҁ$��_�)����
B�O�c#Ck��ǞG�Zr�n	���nڑ�F������((�ӏ�;�.#���^���`Cv�,�B9�Q����D{P����j���P�d�~>��U�|�a�����Z5�F ����mD{��3�=���4}�ױe�DՁ�ٿ�ha��5ԏ�d�~h�Ye�,�.ϩ���b����`r�����k~%�)&,�KlE4cԣ��Ɔ��µ��S_	kQVA�O���U�*�~i��hN	��;Vw#�nZ��|����m�ݡ�~��ū�ZB�hL�Mf��j呗�/t)d4��Z��NR>ZR���k4�f���Ζio_�x����r ~%��ub]�EVG&zSS�P4�+�B�3��)r���x5��F8�@�ѡIl[�=��j% �S�����2�/��I�� >�!nP(+^�7[���ܣ1�8͎�c��,����%�A<�p�9B�.FK�0ы"��s�8��Ա��ͥ�!=y#ۦ��T�Cٓ,����ۯ���룄��t�����ͻ)������x	�k5<E��/�	fd����Iŭ�\!�o' ����%'6NhV�,� ux�:Y���s�ȿ����o���	�zcn���puez���SH��<�oZ�y������7�^���y~�c��0���A$� Z�*�>��=�	6�:���|STU?�N�O�ɨO�2��搆{<Y8�X���^m.NHŌ�*���_�f���ã.p|�$��Kd�cN���9�0]�Q��k#>�p�C'Me��T��q�����H"�ȓ%ē��IN�<��%r�f)!��Zf)%9�$��NwNZ��l��}�c� �	r�DW�����c�Xg�/��<;Q�A�ɊK[�jC�/?;t�����0db�&��s ���R�8!�w��aG~P��3�	�q�Ě�G�b�� A�H���t|���F�R.c��
�5��`��������f`����f+��\�i.L5y�C\�`��Z����[ix3%�IXϩ��!�w�n��,�
���
O�O���
c"n�41#Ĝ���r8T�`����;���� �7�7v���UV�Ҧ�o����9Y�r���_X7��PM�>Z�x�#�N'�\��N�f�:2�������:�4ֹ�}�L�/e�l�#0�B��z�jM�󲽄n�:373�6ȗ����ķ���:Z`0OW| ��"<���SV	�<��ת;��}����F�j��}�@��?�%%mK&큖W�wf��ױ,G��������T�4�f��R�*�[�����e~]�
�������M&����++<�)N?�,�ˎ@��3�崽�,�X�k��B~���ց���Ȕi?��V`�Q��$鬠���
����Pz4^�	O��y�{	d[p�W�3���kf� ��POj����St��xHX�̻�-�Ά�>��*'�%t��6)��~h$��Q[��B�O(�i���f��Z�������'����߆,w�&���>�ٌ!��S"Z�R�Ȅ�uu%�����GB����"%	xN������;��Vl=�y����>�}^02Iv[��ţ��n��]��L)>n��f�5NWF� Τ"����v��������F�v%$ܑՍk�wx�(�y�K� �������8Z��J�,��p��osbS�����f.W��B�t��T09N8�GERy��dYӤK�𮪸&K�9 h�N?����oT�h�Xh?)G��G�~E���ʼ��1g�[����T��@(I���sx`*˩�'Єm;+}�h[8@��%��j^s���k[p/��Y,Zy�0����W��-�_K1u�I~ة^"����<F���&i�F8�m�Ѵ���R�4]2h}(�/6��[@谗i���0�������z�rܚ2��<������6��F#�	��g�
�m��܎��mV�tC�K��}p:CL��h������ŭj�0���W[_W��؀-���{�����?k��jĈ��{q.,�j��]�%_��^`}�\
F��՘V�t�CQHd��~��m'��N��D��c�)\��QgOv����j��C�bg�X��	c��%f����B�v�?��;���me[�`Z�ٹ�cF������_B�� ����xy�N���
d�G=���[��%�ZI�����oT�&p;���4��
���X�?4�|igmA������@�6;��a��49������!����/.$�RKW��"�[�>P0��c���֕ce4],r�(S���"X8(V�:��Cr�t7���!hH��G�����σ�8����G,���av9>xbsF�4��P	��?�)�����}jD�"�tZ2��+mB��Y���:�3�JXI)���3Y�I�%�'sZ��+����k`j���(�%�Iq5���:��j��\<gG�A��cW9�̧���V1��:��/X|�;\��S̥i�I��\O8����z>ڼ������V�� �n&��`���P�c�Z|J�����������D��ژ���mz&����_	����)�Lb�����f���� ym�f�=�C0"���H�����\т���\�1�F�����!	(�����S*��
�S������ϕY��QXGV��g�0�w�C�?S�9B�?˓X��CC=)�&����#��"�p��i	����٢�:$T��_i����H�R��v�o��	�\��ɡʂ1v���Z�m�Wx����Ư �e�oʈ�����ӛ{1|1U�ޘ_�X��Pf.��5��q��Y)�c$��C��Zyo�_�����oM�S�	�3�#�S��Iˌ<b��/��O;V��bT��{A��<��X�Io"u�	�M��$1.�DҠ�y�K�R��S,45t��� ��ݕX�R�Nm�;����\�?��A�F�j�VS�s�=g�4��,�t��=( ������0*��9�u7��~X�{�]����=��L�J��
�]6Sx��U Z��:J&��]�9�h��'�-�&v;��1I��pKW��*���ǥ@� D�L\7:>	яφZs"�T�Ĉ��w���B���խ�[]�;>�]�l��Z�$���"��!R-IBl��s8FY��eԦ����z��5�bv�iu_�Ȏ�J��j\�M#BX��r�MaK�_7.6_�%yT/��5��t��bb�hp����pѨKKG�AS���**�o-�q?.Z�F,�gd����t�\l�&�͠�
�&|¸ǥ�3L)4d��$�*o���@�p\�#m�w]�"�D��*T�Q������L�;s%d��?������c�P��� I<�m�c����m	gsyb�S�9Ê���@���d�>�W�{s& ji?�� ȃ���Ct�Kl	oJ/Lϋ��8���D�j(�)�	 �Kd�=UUF��T>�\����>n�:̿Q뽂��s�~�čz2���t�62ڇ'�P6_6Pa'�N�w�NPH� ·����>�����7�l�C�?|T�\��JHF�4q^���FN�8]T�dA�ǀq՛���+�N��!Y�z��b�Lu��M2��@�%���hƞ��az�Ш���`T�VD�L��D�v�'�1܅�����X	�f�q��j}��r
6�}sH�v̢@L����)��?���V�k�n/��[��n���):e!;�Ⱦ(bS��R�1Zؘ$iw�d?��aLF��`!B�\�'�T����T7�q@Nzp��u��x�B{�ės˂N9��A��{Izv�	��Q\�NQ�z��o�"��5�?������ؔ���|�`0�@�X�`�%�<���I�Ɩ�ٟ��T�j�)ѸaU��d�<�v9?�$�ގ�^Z�
l����y"SwBC�n�DL/}O�˱�c�-%��j����9�V��/�nԖ�S���+�,@�Y�7Ԟ�B��|=M^mi����p*���h�x�	v+���Sk�s�fɩ+??*��*G0Vm����ưg!����M�X�Q��I�nIh҉�]D�7?�d 6�UΣp�Ӻd�[��F��Hpo(��r��Ź��;�(8յ�K���p5��~Q�Nψ#���=�=�e�����3��3��π��^��`߀��c�t]�m%�a��Ơ����08�6�	zCAYS��u�9�[�\�P!�c�PR5P-O���/����<�ß�@J��1�H�0��NAD`Ψ���cn(��F�V�r�n%�0G�ȟ�Hׯs�aYB�'�c`�ܱ���x\:+������Y�����opY�y��4�ۭQ*C��2�r��cBLR����(ޢ��r��c�qG��q�֞���E���s$���Hǘ�R4�	�L�p @��l���$�{�.Cy[��a��3u������+�=�B"�O؀�\��ɹ_e���9���C�ɺR!f��qG�:!��&��w��F���A):�j��@�f�M܎��8Ȑ=h"@����|�d⫁e?��e4[ߙ���nn�`�?����}I�M:�)���^���#��b�Ex�A�rE���:7O)E�Qڻ�ʠ���\J�ੴ�3[��X�˳V�B��hnwȤ��U*�x��Zn�ݲ=5�C�#�?3�>������?�ЙXLe�7v���&%�;^E6Ƥ]Π�e�ǵ�&�<��΢f\kr)&3;�(�J;G��?� ��`�%�z�+L���vQ����1��h�>�n3�w�k fU�fV M��	~�L���������JWP?��6NS^�����CN�Ni+(؎C˧#����h�'��/O��ԅ�e�����7A�!�ڰ�U�_��z���r����]b:G�oY���ŭl�ܼ{��1m�(5�����t@�5�7��쟃�	}��IDO,5Rto�&�z~�w�r)�=i�|)C��(kg1�0,#U�wM;<�E~%��":�ḧ́��jLR���4����s��0�������� ������C��#Tؙ�2:���Av�(�Y�U���wd���E���E"~��S?�\1g|MObb�����(��G���H߈O6��*&���h�Y)�
��i=>d!����5QJщDn����(���F��b��i�*�fxm��6RPid��p��o�����ɘ�\ay�����rl��f���q��V�"�lր�n�FB��Gϲy�b���{�1j(�ku�2��D!��Q ���ۍm#�M��i�mY' *��#Uf6����谡�J`88�WZ69��w
��O)���(��TR������~�Z,�矽 ���G< �����k��?b�*����\��Ut}k�bǳ
-n_���[^7"�.��a�*$���T'�q�]-��O�3��㌸u���Ɯ��*٨�y��0A�
Qa����z1��c�Tj��Iq`gM��*�����'�ay^�$� �s>�q8���o�"o[U���<��i5'�V-�MK��W���c���Fq�޿��;�;xN*t���([�_~0��#��}�[܍X��%O�EF�m|ھ�	��:����\���o�CЬI�1�ʁB�V�e�c���$h�^�?1qSv��ۧc7��aǼ"a��U�1i���6}QkH�"�ل=U���H��ӦŖ�^������P��À�O>��ÛD��Rf�|	*� �H���0gKԑ�D�m�`V�KT]OӒ�Ȧd���F��	�:�
I�o�������v���-�Iw8Hp�tA��d0���(4�i�S�����5-1����xЃ7%N3mB����]�24���K�կZ-��H����(�/��R�?�V�����0�+���);��/Sk�T@���uR,)�b��?Wίu{���1��H��#P��/��*��=	���u�(k�4z8���ij7-�c��f}��T�U�����Q,e=�}���~�.��b�|.LB�3��&�;"e��;��q���O�H��
�e���y�ּ� Z��r�N�6���c��*+u}��G^��A4�e~a�wPBV��sc���]��#B���9b��f�R��`1��o�5�n��&ɗ<N(��B��f{O���Tq	E}K5m�0g\�l7��Q_R�F1iV;��G�
1��0G�Z�r�Y��1�F��
�F�c�uXF�wi��C�(TAf<'���!�,��v���:�c#�f�A�{]��V��97Yn|�N�2���+T�.${��o2��]T5�!q_��.�N��kUS��E�e]=��T7}W�w Gy��0��$P��♅q�=�����e�V��>
�b ������@M��N�?�G��\ξ���O����AX��l� a�de��(-��~�.�s ��ޑ)Ak���' �h�<�)���c&��=�M�����?C��(��B��q�<���* UV�X�gx�f�p��@!��KF��d��Hĩ Se��h#zP:m+�iW��i�
U�dő �1��@v4q7m#�{4 �8����R��׿!�B�%�;��m��px�g�b�a���_�W�l$� ���͏�1֌�d��2ш;b&q�.e��� �LX%��B�£�Zz��+d�o��ьG���Ո�|�0����O�Vny\8\�hV�.B���	�m���ϑ֧��e�74��'b�-P�{W��<�`���"D�a�)�h�=��=���S\�P����C�f���b)ӷ��V�S�%��慶�ihl��K�޺���ǵ�^P��y�Y:U���$�����Ǖ��4h��(�tG�Jy�8M8�5�
+����w�"D�g?���ۻ�v/B�pH	Ҍ��pt9_���긢�����姘�4bմ!Rڎ�_I���׳��S�:��F�|$�#aҳ$Y�Ω����]i�v�WL��!F}pTZ�r�龳�5n���i"���X4��#�WG|�<~��YK�xE%y~��l����,YNlJ3ec���̡��{pٍ��Iρݚ����.��wtm�,O�n�W�S�@Įh�)�C��H8=I����a�&\p����)\�7����/����`ܥ�k��ߒ�B��g(J�R��p�a��w���t��9מ����nX���ܽÞ��́�-�+j{��l�$\��������X�p�zs>��|��� L�u�tVAl�k��s�sg�l�gFi�$N�Y��`��rc�,N�2U�gXz�B;䒻FA����$��	���X��h�A	e�.���d|]��P����*=�n\��]q�<}�@����y/H���H��j�/݆���b��=R�v�hi��r.M;9���5.����RT6��3)� ������L	���V9,���ZO�f�j�5p����5�~�ay���X�{�8�����fJa�y=�:Wp�K2/ۙ	��?;��@G�/¢o;�n�fߡp�}9�.Ô�navLF���^���?O!f욋k�B[]Q1YY�)F@a,��IE��E���Lsg΂Q`����kּ��G��E/���"b�Iבt�x(��l��[ҝS����b�u���ͮ�	��W>4P�u��GV��cm�`QڳWj=����Z(��Ui��� �/�%cAԻw`J%�5�å~��*��p�:w��/�<Δ��-�O]�_�W����i?@' 8�!����+��̜���eR�#��j�1sB!���x�_ �qd�Hd^���!�P F~�I�,%]�.�IrJ���)L
� J9��{K��U��|����F�����N�Qʿ����"O��&ASO2��ۦ�_�J5O��q2����+&'ʁT$��XTOএ�P�s/����v\�J0�t�9&�u�z2�� r0|SQB�u  �n�z�W�+
�Z��~`s������g�8��@[&jd޺eS���8�£�.I�ɣ�[�_�[�WvYgis׷�BەG��S�lV���^�<�$6E���e܌�s}���*?{wi���H��H��E��¼�� �NɆE����&n�lÊ헓���6,HZ����(��5|�\k�9�/!�D)��0��(��$8���É5�w�-A����2nr��%��SEh�M#ha���ɿ5�wi��ޫ�Uf�r9n5a0�9泠sɁ�}�x�a�i��h�7� �?�ճ/>��Ѡ"�����nv^�mx��'���1��Ĝ�(�N�ċB��u���� ���^�W#�	/�_B�L~����ͷ��!��e� ���~�jO�T�w��bgwa�!I�~b�,G���E�
bh�f�E��*����{�m�n�ú�6ʀ���%p�eK�Sp��"# �W�����^8�a#ǺK)��v�!��Q��츉��ɗ��*��X�Ț��m.��$��U�kX�Q��s���۸`�w��R��uJ��KR�L�����m�.��"�"Ex���'Nc�5��G�WaqY�E�.��=ߚ;r��%H�������'�s���8۫-�c�z���#�ʐ {xz)��|jk@���{�:a��T�nbX���~h�ޣ8��
�uE�Y5��8TKf���;�_��Z]hi�m:b�d��P{�����47Z��R��܊w}����wi��N�r�I�A��mE>#¼�,�>8x�� u�\�S�Yp5�U�&��q��I�5�7��~��|��H��`�8�/�pQlu)���5��I$m���?Tc>6E@H�Ƭ�1%�,�dP0�2֚G  ]rw<UGS�+x�B���`��3*�n]��h%�TM�� _���n���پ��:��K�es�x�P竆���=�2x���^����G�&O��d������=R+Y����S{WXޅk��z���}h-�܄����W�:H#vb#U��ZIٻ�F��	��oI�����}��:nX��:�Ԋ�w$\�-Hx8�QĤ�(D��S�LM� ew��G��Z�Wr�6̞w����4����*�C��#s���n��\�\z��Q��1�&�
zI����((,8�I�-�6��wj��z�9�~�H�t��`�d;5�L��cQ|��T���_�_�nK�����h�"ԅ�7�7�A�/~�l�G�v7а���jKd����UR��X���\�mʴ�
�**��	K��Z�M����R��A�=A�����t,/�3�F��Eȑ	>� S�Qvײ���!�����((�Yן#ͅ?틃L�@*3���b�İ�Ήhg�x���H԰]���U.e`}*��=������`gFDh{��C�pj%��#���ϟ�� s�F�}�_U�=g�Z�~A�B6K���ߘ����&��P{�����R�����G憦^�{B�"�
5����  A��k��(�-���	��j��l���]*}�f5�Z=��\��k<�p&�g75�ǛE�l"r8��:��L<��h��$R��<w�Z= �� "j�8j�7�c�z����V3�4��}�&Vț�l\+�Mu�_��ݯЉlh8\T�da1)u�-%Bk�E���G���ZW|����n�X����v�e���RC�a7B�H�8����%�F�e��ZY�>եAv}6[٢ �������`L��b�#�ET��J��ZUq�o���A����z�!jos,���>�>���B����9hl�u��1�UI�~VG���@iq��R�*ݼ���uQ N �D����Z^��},����/6���A<di���K!7���jױ����	��Mp������ ��S�Wm1W�a5}1�u,��oW�I�J�d�l%t���۲\c\@��+{���Ñ��	��V^��6�h��Z���I�w5�T�� �d�NV����?�Ȑw�̈́�%��������k<������� ��#��'�f���!�o�T)~�j&$H�I���({[�Υ����n�ֆu&~ݧ�ל��D}@����^n,�=n�Y�UGr�5{"0����i=4���m~B�E� ]r�x����;�@~��w){�%�\.��?��±�F���\�ʩb�D�s�L`�PZw�K��&���/sgl�A�������F���v�!�G�=0>�m_pUB����"sU�M��4�
D~�e��CR_��Q�?|/���'$�'��~�|��m=��2��F�O�.v͔M{�X^{���u��<���ԝA�u��몭��ò���4�C	r�FY��C���XHZ�M˘�
�㌂J*l+�଑5�r��
�qR��*C�B{�B��Sb���&,����G�N#�h㎼4?	���S0wu�Z�]�Ur���Q
�7Sۿ��zv`B��<~΂��8�A5ږfϫ
&�m��r��H�ަ#D5���8���ј)Q�S`�W�^t}�����d��b�v�j��P��P�X��cz��9�t��k�`��E�5��I�D���S�ai6Ls_�}�\W�1K���i8�P"�AGq�e9�S"<�ܯE)e �%9�q=\��犰�����)�*�~�<r�<��@����F�=ݐ������0�&s�d4[�a�Ȝ���� ������cI$#���s 7�&���c�؄8 z�]|߶���]$2.�N�-k�߽�����8���,��+o�K�5��Iך��ۮ� �'(�T_�T	?"��ր2�%WKm*�L�cK�Ug�da�<
�rQ>k��k�q�+����������.(G�:�����.��k%c���C��V?ʕ) �f��F����'�ߟ����!�`Շwwu��}Hu��ٟ�od;%���S�5����r",�� ��
���6,����6����^T]�Ng�߶G��3E~�-O�;�.��y�^�
 �_���׳9tX�-����i�7)P%|��K�&^��b �))~@��,�{`Aȯnzo�p2����Fݒq5�k;\��f"_V�0JD����TA	;cʄ�g@����u��F�ڞ#Tc ���8�j��\�&œYI���#@��ie_
�����e�lcwo����Ky�见(�n�ti��&J��EN�P]�Y �P�����XS��=���P1{�R��ks�.In�Lo���Ϝ%h��n9t�0�,��%���3����(O%]��R�(T1@7.vY�S:��^�K{�2a���c)����U�|��c�bP�_$��ϲb�*�ׂ�t,���שO�=���_�cyy����щ�p�@"��}[:Pʜ�
 c�}�س];� �K����'�T�+��u�"��j��"�ҍRdU<�G�-h;#{iQj��  Ď{K{1B圞�{(��l �s`�r��70��ƽ(�\1Ǘ6�� �� TA���v��%B�1�%���1f��PN~-@����G���{c�,��>��0#���`����k~�n��ƣ�X�'?��q���10��9�?<ŪD1��j-�WI�s9����Q�z��7����t���9�Q:s������t���t�Y�d��|1h͝��ժ�m�z�X��B.9�qu�6���7�?}������tNA��f��q�y#�ɹ�[�"�A9�!ҁ�6�S� "D��"��p>�J��o7W.����`�,j�p���>�� ?p�����Q-ݑ}����UXk�G�M�r~�]vӛ�1�</wG`<���A�"����E�zt�:ۨ	Fn��}���0sC��(\��J5����R��u�\A�<,Ԡ��eO��ǝ*�\�>v�a��p������jt���w���lJ�Z6XsH�y�>�ۮjhX��N�����N��S��}�����~+��n�̈!z��i���q�u�}�sI�f�f��ҎrSPm��
��{�v�ҕg+�G��;G1Ll���Df+q1�Y���s�f���:J�R��R��94�Ӭ
X�}GuB�gm%4Ѱ�������E���2����&�&�adSm�]"/pX)�[�<fCLi�4�	��4�u�㢛�kH��5tfF<��������:�e�9abR� ��Y�2\0��d ���|}�'��OD%X2i!q�Z����+Nx�.�Gj��8�� �I
���I0�X$s�e�Za��	�jn���|�[���$n��Գ���R՜������ۧH~��g�p���c"�G����1&����Yp�A�yޢ����l\p�\9���ۅrx����z'��ri��%[��?�}�����as~�dTe�I +ӗkM;�q5����5ϸ剢��,�Mݒ�r��$�)_��wg�_�[v�(�i^�]v�.\sgZ�m�>�g��.=�@L��/:%ϻ�����z����O���M�pH;X>��eW$/��A�����&������Z��H�eU��/)l������<'c{��i�F{�7����5�K�Q�u���XHj�D���~�Dή���t�D�j,�eH�̴o�s��dh���ߍ�qxӦ%5�Kqw��NArᴌ�Q�n��}m:Ӻ�R-�*�M��̬����L{x�d�#�\�Rߎ�D3Vq�U��M��8�Ȏ%�t8�̉�`,\[Rz��
��z���JUu��g���s�ܬ��ֶz�N���)��q���?�R�3���\�m�W��n��s��8��j��M^�[֭]k�|z�H���h�_LdV�4$n{�S����f�ORwg  �|򣂫~U�d��e�Vz�?Չ�uw�_�ŧ#��?g&��L�C��~�Rf�x�u�e����;R��x�2�.]��t�c�qEK��#7b�^Z��܍���۞�I�%	���S������%�Į���ݑb�B�?��0�,f����$w%���~�DyX�����+��1�M�ć��dM��=�#R0`���k��V�U���<��b�ɇ���Q��{��V~��b[���$��jBs�g$��x��
�6��C��P[a>�S߾�r��MsS����P@���PD�f	S�.	���b ��lѹ�;%��؁c�՗ݶ��>v��b^�K[�%T�y�K���I��-:�R���Čf�߭G�ŗ�.��ԚU���ܷA%��aĕf�O%3�}�{������Y�������� /]����;I�_ɉZ#�0��~�&`��Y%/��۾�:�������j����橊�%pH{���N�-����X.i�J"���^�!��|g�3��+f`�#L�u�fƪ�zw�����V�aZ.%'J|3J:�n�R�A`�Oml�c��lHUx��2Q���CisCX`3��:�BJ.����z�}��1N)a�����2=ٵ3df��Sz���J���S۱u��~P�z���I��&v��k7�Q��N��,i�t\�aNE����5�xZT��r��{�i1�Q2u��:ڌ�fC�y`XO����D����>%R�W��,�ٺ<3�iq�v���Ȃ7u�__G�揦]�1.xv<�L��4Cϼ���:6Ɣ�QY5���<��\�oo}�F���Ў��ՙ�l����J��9�3ie���z>��ui$�6p5w=x�݀���^��;À*�Cn�6�� J�NlI�T�&���p��m�5v�V��9-y�s�J��~}��*��q�O]j�]*������R���6�%�+U�1� \SOI���HN�J\����z�1����ܼ�=��HT�H�{���3��Ȣ�h$f8�RЕn�뾲�'1rӸ�Z���QU������Ff8.�Ca���-ٝ^�:��q@�2b�ٱ���=�������9��j5��d�j�]���E�p�����7�Gb�woFy��5��W�����9P�j1�I����˧uh����)���,�o?�8/��չ{��w8��3�6�CV'�4Vb�P;���VǺ�: �Z�.>�+�^c6Y>� �F@ь�5uL��;:��AC���˸0��D�Gt��]j�#g�4���p����k���l�X/�m
2O�dO���5|E��Y�ѳ�q;p"�D�$I�EN5�(�/��ޫ *M��i��x���1햍 =q��N�#B���K�"�VL�El�/A . �{$�&k�A��;��W��)	Y$�WR��ڸ�Y�h��WN��݈����;1����<� >�]<<�K
	���Mqmߖ�K-ķ'&�!� �z_V�_~�m��/��=`�@�]��M�KX�k����g��lL	ׇ��?����Z����5�ؐ�0�Q��/�"�s;��>�z1d㻝j��'?�N])Џ�/�;���[u��'gXNpf��<��yV��#9~��;WmJy�!��`A�'���ZA3���Z�.��� X�6�иE����=mf�Q�J؉�<���㶦ޗ#��tv���i��r`h)8��K����9װ?���|�Ō��zw r�ºl�wV�xM����mgg=�|�_�ga��K~��<Po��J'�r"����j&���Qv޶�'��l@܋��6�4��wG�,`S㞫���z�X�<��)�o$M��d�X�r��a��~fWW+�f�~�M�Az�*��<��^���v�ݿ0�y`)vW��B�&>\����`���� ��M�Ȍv5��w��&+�K惥E�J�8Wn�
��-�$V���`o"�oV]�����fsDI���K.���Jo5�u�G��z�U�묎ȹݯ۟�o��/��� �Tw�v�� ��9�?y�
��c|����E{�B`a�p��HΉ�TB&8J���ߟϦ�직�4|��Y@Ҭ�GZ�<I�S;e	�;��C�j�a�_z�|��,�BA:5���g޺N�q�RtI��9���p�E�F�Q��'q��驒��%�{�R��/#�NT' �΃cfڃ��v�t���E�?To �g���:+��1)���FƼa6�����O��>H'4��������a��n1T�O�j�^��0q�K�>���`m�r��mm7���8�S�J׼���e\Q/�U8������6�׶T�r9�&e�7�j\�~���� �6��)����B8��"��}n��a��4y�`j{����˲I�y����s�Y�puWqB�e��0h��l�����&#7�]�����!F�{�c�ğ|��\�7
$��ݟ��<�E4��Tf������uJ,���d���C�iTLM��e�Gr0��W�!�