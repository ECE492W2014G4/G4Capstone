��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P��v�"<ߞ��&'��k%P碶�R�ӣ�sĞ������FY&<��� H�f��G����h�H�xI��5�-�v�Z�qRG�8���LK�J��_��7���l:tl�-N�a��A������ʴ�/K�&5�g���I8�W��^���_d�5}�L�3�%�k�5�D���@qc�w:P�����-2��ߔ��؉8�P�n���i����X������{z4�ao�n��oP�B�����f��E��s
��� �kǱL\�(�~�6X>¿g��զ7FD���.0���R{x9b̿ݝ�Oli������^���^���0?^-{��M>/_`t9��pƬ	�+i�΋x>�"nkq7���a��=Y����h6�A�I���Ukz�h_�_"Y��U�fW�i�!���R6�\d	�=�9�a� ��W��ᅱ/���_��:�|.�}X0���@K����~}��	<����nRοK] �?EC�b"��������Ґ`5�=�*va����W�.4�yY��f��L�:SQN��]��TD1�8��J������G��n����w���4S�&ZJ,bW�%f����n��O �B	��bE'O��a���H
l��*�\�:7T���Ej���nH𣽦�P����.�rկ
�;�&V�g-�\�ߎ��W�HE;�L۶�Z��M�m�ήro��`����~�Ϛ�`M��У^�6�}�,)�<{����˞����$<���J�����<��R*.��6���&LVr��RtQ)�Zg�i.�T�ܰ��Q��{�0B��M�cxޞ*��H0�-I��F�R@���T@�n-)���"�����]�҈�I2 ���y+��3������j�#ّ�����!(�{\7�	Q���L��6�jXU�U��H�DL����!ң��y�Fg��	jd^��e/�+���% �=�����/�Q�h����]s<�0\B<%�h�j@����?7Y�X�8$���|�� k�`\����z�����y�Bac1L��O���6K}��8�X���m3������]���.��m��։��c���N]�d'�jY}����Xq];�ț�/�@��Bߐ[��Ml�$�����]Q�W�<�/�0CY�o����T%w<����ciK3��t�=ƛȍa
V�U���_.ʽ.�Q)2�/�K�z)�3�E��,�i4���Ό�08��16G�7g��=�<C����F�"'���x�͉{J�*�B]IȪ��ħ�ߨA_�+d(��o�w~K&��Y�*\>����bNxm�q���$��?C�a�,t���4�c��=TVQ�벸=q�e�-�>��x�E|����B6tiOW��
\4/U2�+��A�KD�s+�$v�f%>6W_�h�A�E6��¼��p��Cl�\RI�eH�����r���zN����K��>�^�ƍh��J���X����.��̅X´#[��N>���
��OOlg3��p!f����` _�y�P=v� 3]�5d�Ya!R��y�{kE���(( +�2XXf��Җt��Bw��2��=|1����.*���8߅ų�NU����.���53%6�*��:T]��B���M�oɛ!$�vŻ�,����jW|>��k�&l''A�E}(QzX\�]I`����$�����2��#o����#}�뙀��p�h����q�pV���D�W���(���&3?�.6R���E�.c=��Dl�|/�r����xHY/����#��K�vT�A$�{�ب����A�b0#�8ߖrP��,�������(�U�����X��
D�$��s�_��)i�'�\�}�mm���$� S�,Fj�5��(|wȨ��O��>�'��V��H�r�pYbu�]���,Y"Ǹ ���dr�h�i����.pÐJ��HP�dX�]B#Z�<���0)�n�Z64��.7�qptY��$�a�,Ao߬��9��`�6��=���]xr{ι��|��Պ�Eb�9��:;�}vL�n"��(���bбi(�����u������9�j&U����K�CƎ�܆�ar���s;yo�'Wl�G����M-�����)MV��[_۲�����u��0�Ost*us&�[�t����2��?p�f)D�����9=�8�U31�n�~�n�$��t�p�n%�V�A��X$�=(K������[!�����J��PK�y ��%�ު��W��eE�fo��3��d�WGǋ���!���.HS�ˈ�Z
��0�j�;���Bm����ĄF]�^��\޽XX���ԅW<�_i��sB;$9�=e��m �`����~3����gg��C���q�Č��q9gXtM�]-��e0uiK�M(�:8���6:��}s/��5ʕ��Յ���߇��p<6�۬�`r)^j�	r�c�H��_��[]�3_F!o0LoF8���xӀOk���.�2iIׁDh\�d�
�u`@��6<���C��;�ŷ�|��&�S�]\>���'éb=%+�*��w܂��n"�|�2�T�r���6�!�43𣰚��#DZ�@��C�����\>�+ۼ:�{CG��G�l6M3��8�v�to?�L�F�f�'�`�A��QBw�X��Jn�����g�b��`�+}��:KHK��_��m���� TIɲ�2 ���4}�#�|fꌌIYѹȁ�����ej4�=�"�i{�'}jֶ��a
��#a4�7���D�X5=L�юBb��w#�ՙ�D���U�[1X���N�1d#�	'Kv�.#�7�Oe���R,���>�a-_x�OP c	l�I�!:}5qd��WN{����P�yL^3�g�h,&���7T�����?�X��JR�,����r�c���b:ғH~��v�����ޗv�N�Hz���u�d�:l����Њ@����p[���ô$T\�uO,�~���݇�9�`����k�۬���]�(�e����S�ud ���Z͖����7���9��y�fI��4��	I��OV����:��)�"^��U���ϘD
������}��Wd�w�pM��dJk��3�	e���W���#��X��B[G�k���q$�lo���:�S�ض&XE�<��e��ѬRb�NW�"}}~��$��U���g_��<���T��vYi�F18m��c�������£��yV����;�`�=���B.�ѽm�7�g��C��}�GZ��Wx�XO+fB�R�GZo��n_�~���ߥw�]׆;�D�}�2�"��i�~ �f8kk�Ҁ={g��W@'%p�0�2?�H@�HO�R[�iׅ*��@�<��F��E���C�G��G
�Y�FM��S��rg8w/�k#�Ϯ&���X�9?�.�Ƿ�y��x��=�9�����U���P�W�+�KB"��O6%��Q�:� �X!�������Lٲ�j����b��Ч;����Ԧ{����}m^sy�I�-�h�#������\ ��@��+��A4�'�vP��`��n�۳��~=��E,�Y뫾�Om���9�8�~%`�|�tDr"x�J��YT��%�gGx�҇3n�76����~��^bO�Ԅu2a��li1"���|�os)��a�� ~�\�Nr�S�Ű����׎I]I�${&��$���ī�E�U0����VG������r�e��"u(�ۓ\vQF���O�2VOeBj(	b��\����q���ߑ��keA�L��P$!){�g�� �n-wCh��6v��\���t6�
B�g�U�tq<H
&T�oI(
j{%%y�Z�b�D�<�	���5�;)kUrPk
&�y� �-R�1�M�]���v=�Ky�s�cJ����[���۬� ��A��~��"�{��+�13f�%�n�oR�F�8��)N�^�s�Mr���"�ص���b[)�k��Р�x%�3a��̚��$�e�.vRxܦs�H(_�ÇN҈�)��w� ��	����n��ٗ�徽��&K���k��&ڴr!h��<�����R��Hgz�L�����`�vS��6�����!��)RW�v�@�b�&XNj=wI7��fFm5Q������>��WA#�֦�S��ZU�)��+�5�{�]l�,��w���m&��w��p�D�����>=��4�ѤA����|���]�\���U��`aP�"���b>��C�Y���6�a�
�<�;"T�+���������n]��zV|�YT;=q�=���5�z"���C�C��dI���m,NE��Ń���S���>�� ��򦞟�U
�dWR%����c�iv���);4�ԆR�@�4V�;��b��s;PG�w&�.%�y0�T2�l���W�6
�����ŐHb�8�0���ؓ�-�Y5/�i�"��>��9��#�~�CW}*����Ӵ�_����%N�䨅q�Q![�S��҅I-5�hG�a��g�!ַl������� D����.X��"�#���h�$o���:.���Li��.��W�@�)� �����ג	1rr�h������'�(��~�FFg��m^ �رGH�f-����Xg�#'\�"�׵"cv���>��W��m�E8>L>��b�~M�tY�4�>d9�t�b���ލ�ϕ�9�7:���>�K��2�)��9�GΌ6��S(�X�X�1=<z+�3���:��*;u��O�0Ͼ���j����$҂&��$A�X���^�U�%�(,L	�9�@�=�b-��W���իo����ھ��.U�wv4�+C:x��>r�g�u�J���=%'�*����s�#�ܳ������jc�ӛ�N�3_�]�@@����%|<������S�P���{W�z��4����6�F��F�/s��7�7���g9_�#*z���J��x�F�Ŝ��+NA�S��ɯ�IӺ�?C�~'x�%Uۜ�;��"�r�2��垾P�U�:�H5�NZ�� ���-�1�Y+}�t��O��R�:l�%M|)�[U�h��T�A�䡥d���-BW����r��niUvz�1H����3��(�=�v㔠u���q�V�q]����_�d��y'�F/�?ե]�R���7��&�E��SE���t�/J�*ȓ�ߓB熁^��=���WԹ���I�4�:N�Dg�[��i/V��HW:K���#W��y�V̓���Z%L�ֵ�g�w�{
p(]�	Sj6n5V����8�ÿ8��ç4!>�d�� �Р��7A�����y�½��I��(��i�*E�r�����~�� i2b9��0Cb���W�mӁbt.����U�JPMf�����6u�AN�նG�DMڕ��[@%l�w"�����!����^�u���		�<��c��b��U�p�'k���L�_�l+o�P�l�TМ��C���PYR�a/��)�ᓟ�G1 *C���x�It���'�x�a�؞ў��m�y^�|퀊O�79��C�:%�K��}�S���=�G}�q�W�@��E�L9=X�i�aù����|�t�qOq.Z���J��l��G�}������WY}�)�� Sz��R����b!��uK�'�\EA�u�i�\�<8q�FHF==!H�'��ƙՕ��0���M0&�2�8���@��T]��L$��Q��L�O^���EF���_�W���ְ�z	���;�Fl2x�M2���\Z���:��t����ͻ�#�l���P3lb��%|�pWf>����3�`yϸ�C~�N��Ƅ�$N�H!y��m��8�g��E��W��p����7��}v8@5tN�MⰚ��)�Ѥ�a'��(a^�G�v�~�(��\��Lj�-yf��;n,�ޢ=����1
m6�1����D���y���/��S�V�ǟ��0�5�EV8XB��)�����٘�m �E9��6�]<�*�$��՟Ƨ�b��zȚXF�j:���z�Z��*����7>���9� !%܇L1����������Չ�"�iZY4ئ��ĕ]}j�a.��A|ݮ���"$ e�V�Af��S��c������:? ���6��[�8ȗ�y7�~��׃�I/�e�+��|�'��L�#�h`1����K^�x�F�,G.�9��X^�o�yN��daV 2��fI��ć�<�2�V�QW��;x.�R#RV�?v^2C���'=l����%�#.��L!X�6���OBÖ}��������nw����L �j���?�ǲZ:6���2��Qހ�-��f��6Í2�����#Jb�]��db��`F�p�7�19�d5�sX�/�87-s�����jT���X��-�C�{�(ݢ�JyXdr��8^/�gƶ[+�Ka�mR��r�
?E�1>^�Z5�Q�aj+Ɯ?vI��J�&0��s�."��R���;�C���)���6����ʙ0�3�7x	\���
6�n7vo�n"d9듽���-	�;4��@�0;�<�1
fXГ�~EH�7���*R�`ks��Ho0`퍉�n�|�	(ɿ��3���`�"�����d�2��o ���`�iTMO��W��Ŋ���n��?��'��k7�/G%1k���5:`��hD)8���b᫏Y���u�l`���vp������'��_}��0����Ad�'�5��Mvc����U���o����`�g����Kll��I�I�������[�&��S�u�,���/s�dV����w%8-"pi�G%PEw$q�뺐f:�����V6xH��m/%[D���<�oP�T}��6�1��#<�,IB��d����J޷i�z���>�8I ��_�};ˮ��>�u����%@�49%�}U�6iV�/���Z�,<�!��|���8�g-�c]
��S*��I�e����o�{�j6�G�*�%o<K��e�����P�.��GْZ�*�������[��a�m֐��y)XLڝ����Ne�yq��P"�ܠ��5���_z�	X-�E�a3L��o*:C	7B�Z�gD
;����A��[�$����)d�CZq��7�*����&�La������i�d�a����y�n�rh�y�ϊА3��)e�y!R�V?��������U65>��`m���]�4�c Ґ��mk�~��nc#C�y�����,���r
Lj=I��u7�xѷx����������j�"�sC�B�Z���h�J����Gn�,-�"�%�� �2	�7��q�\i?BP_�d!��ݬ(��:������N��f�}�C���W2��_��f������U�]`��~c��!�@�L6M��%ox���g �gf�3t�O��?z��	b�R[��T*�n=� Z&�:ۦF�k��AS���v-��aO�ł����%�j��;{��&%_ R�f!u�+L����YY8?<v?�R��D,Jy�Z7u���9T~�x�p|b$¬Y�ǘ��^�K����jm_ֺfϭ��VP���߮���9�-���R++�أ~>���R�Γ
��Y��`2P�5'�'I-12*&�}ig[`f�:�R~�J�n���a<5�랈�ZR˧�0*�S�z�=_�E�m�.� *�t���`w؏�������2r�z��:F�a��g@���� JQ$U���voB��ipf+^͵%)B]~�nA��ǌ��q��c���霛 ����Mz��1�p��lR��O���:2��˯a��@���}T�06�1	�?]<��0^��[	���v�4��f����cCof0�z3)2��#9��/�)��r��C'�vu�� ��Ԁh���G���j�Y���oL3��s�7Q��0���"A���.N���ߌZ^���crP(��kb��?��S�*3�֞�E��
����3{�j��R4��Y������������*���М��u����x�Qc"}��r+	>��h(�l��=��r�E{[kt��)/^#��]����u���u]�y�"iSFD�����Mj�� �vx�i��oG`���3)�E�`����8�/���������,G��5H�z����O$ý�uG%��Y�����e_���V�8q�i��@+���������zFð�Q�V���7�Z�hߪ�+������rnְv4���7��E@$�� 5}�?舳� ӯ�V�Z1^r%GҝQ�9�aNJЯ
��58B(	�{�L�
Y�Y�{Y=���:L�����x_9���׈eV�e��;�2i�`��QC��Ua+^�eM�b�	g�s��$�{'N�N鸇�!�=��E �% ~B�y~��������xC^�ͷ��๟�	|4b���V�ߦf���)\���Ŋs+&QԛܷL��(!6P�p�#�z���=�9nû��I\���&{����>R"����E T�|�Z���5,o�N?�W}1��yUN��e��2�9�����Q���]�D�ϏkA;���7��O
��d��j����������1�XXifpxu}=�.�z��� 7�o�������(���I�rו��j9��~�'mwLk��=:���h��W�Q+f@��Yv1Q���B}�ƣ6��e-?;+h>L2%�M ��l��*��B�AzV�	0|��63B�O�Ȩ��nn?D�QR>�jx����0Zga����`s���S#���@��:[��n}�my��=˴�=R�e����-I��N���F$i�B�Й4-X4��RC"�k���F�(�ךr��ժ�<��k�7�����+�(嬝��N����>�(���9/�Vw+�uM�~xa�j��m����'c�mR��I������>3��������Nߡ9�{3�6M[{a��]{eoo��Sy�糏}�z�ܚ`��g؞�TO9��e�%��!�F*�T��}�I�f�'j���H��s˓���P�!�(	֜�SW!�p�ԡ2S!m�V�H��Q�̨�{i��M�&�HYIn��j*���G�7�q ��9L��	l����C?+�:[A� X��ѫ�����x�C��b�֐�2-��#(� ��ҿ�BE$X��X�\��ϱ���+X��˼����ߙ_b�I	���px���ot˫dw�m���������c_ޫF�+6�?�`a� ���,�Ǣ$���/.n>[���Mܼ��\���q�N����j��JV��#S}�����%��l+�"�I�����Һ�5�0���і��N�|-p|j�^�:󷃕��D�\�W�A��P�����B�7c�0�������Wk0$�a��_zH��c�T|�]?Wڢ��:f~�y�a�(��/��C*H%of���#�C�,P7�/,�����4��9M}���}�[I��g���?2;]]�����\g1䓀]D�BDF��K�4�cs��K3��3�R��5��árY�~�Y0հG�v�i1�7�w�����MQRi��<����`(Ƀ�"����S�=|ī�0W@�?�\7 ��j�s����KT�}�G*+���q
@3��U�"9.+��6��I[K"�ߩ{��(u`��E�O�mxZ"g��B���tRnl��5Y�"U��|�#PjI҇����BVs����yU=�ϫ}�y�w��P8�8K42��[�1��O0���6�;s\��(���Pi��������ZG��;np;��ޫ��^����!��mh��u'��I���EK��#TN]&5���W�-Jj�<�<{��4h��Gmd�(jY�i���lܘ�5^>&!_�d�̂��������T�A�瘒��5[�k��H
��*xDlR����G��&�	��X�h�t��c�9�J��D	g�P�1z&D�#z�Z�������Z�-�`�i���*Ed�"�c���D#ĵ:KT��3�M�j���	k����e�jպ��CEa�*0�FP�Z7F��g=h�ox�'�4d��LY�Q�'���#bu&cκ��ͺF�E�ƍtw�<SyjT�d!��U�������ÄTѧ/}��,	�ڼޕ�N
�A�O:���=�m��?S���4�K�OGY���LTy�bkq�ʀ}g�y�)V�CV��H{�S��EO��l�N�>�yeB��D���L��\D�����$6�<��`�OT���_�_�R����L�Se5�nΜ�P7�ή���rȴ��M�Wfo������ZN�.O��{��LAI�:�h΀FO~��L㎷ו���4�<ٗde?�-�F4�����F�R��ގ��޷�����G���fK��RO���4�g��.���G�����nʹ���*u���"���N�|�̔�;�e42.�m�T�[���y�!�:b�h|�A:N-�$���h����_��3X�ʕ�_�I�~~�Gx�	@��&~Я9tz�5Z�q�t�F��]�5M�]�=�˴�!z(�"�Xw����)��d	"���&-8G�W�jn�q��@��b�#�B��l�uC�d�K�*�D]A�b%�5�܆tٌ�]�B���=���Pc���� lG|��5d��O��8r{������ċ�=��5�gs�5ڊ��k!�k�ܽY
7ҕg�1{��Y�L~��H��[�8&Imx���F_�rN�v#��=(��[/����^ͅ¿��Őp�z>����0͊�g�E��{�Vi	N9�S!(>��tp���t��q�(i�H�#v!�D(KN�|}a{板PN7U6�� k����o=_�D1��d�hIl�`[rmW/-[d��s?I���l�~>�g���&����0�uL�2�:Я����,�060�<�c�m-�tZ�<��?���J�-�˺�$Ʒϓ1��Z�]H���7����ԨoF���[�b����Q�`�࢞)��EZ�����
�ߚ��B���p#�{����7.�0ߓ)�
%���3�(LL*�8n{��;n?�O�l�@�֬�X�0hJ�4�	�ʲ�\%?K������'Z��$:H�[�p��P�ɂ�[��^b���]{�Ƭ1�.�J4������_�,m�p��c��T
�
�O�1�'Ab[�oT#ͳ�9��O){!�*�3�ë�moQ���#� e�-	qA���y��I)XՔ�K�2�_=��/�C��Z��