��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���2�U�z�[B`�#�� 3�����E��R�=R��1��TH�G��N�����` �۠���<q��c}�޼Y%�(�"�sڙ�AӛXG�{|��AT��x�PL(�]������r�@�h=n�O�^����	�{K�*�q�a�T�FV���:`��Q�օ�H�m�Z<A�=p�/R�ؙ��a8E?	[��C��|_EM!���MP��� �R.Cw�j-1�,?���Mׄ��E��T��� IZ$\��h��I�d���cL�mG }������3���@T�G*C��'���"t�a�3kM�����p�s��7�Q�0�[0�yS-*e��۞�`4�,u H��{�k�p	O-O���I\��vC&�] �oV�T"f��.�=�-ԙ�v��vd��__)��#� !�zL^�Z{����0�(�ɸV��腻��]�k�\���7ET�z^��g�b�.�����3��#c��sO��Ԇ;H'���50���V˧K�/��v��3"�c\Oֵ�����uN�=�R������9����dd7�Ndj��q����/���Sa�d9 �0�Z����"���1�1p^L�����3��Q�Ɨ͘XeZ���cՂ*�I��7��~U���y��	�_��%h��z��r&�W'�p{\�4�0`�oh��������5+4�u>�h��W�Yi]���3�>k	y+B�g�77�ľB9�S4��b91��R���i�)���C��)��!���oz�MFK���>x��J܊HO�arG�G���iؒ�a�h�R�M8���)����炖�L3�Lg�սg��b2�2������_1X�'�Y����*�0 �rt����?������|�{��Z+�X&T���ep��eB;1Jh���ް����*D��yxN\d�Ut&	A�
\Y��a �%�i�"�&m�4��˩)HO�i@���Ww��T������҅h6��T�AǼ�
2:|��r��Q��BQ_3g�W���l�Or��mm�?I�����Oy�˰&L�}n8+�K\_؄']��=Eī�����t�M���@M�ߍ7&�D������������Ɍ�5*��h�~^�#�P�u�ǫ|��Bwu�������)̳vw�`�e�CTxc+Nn��.���0��}��0���C�7�D�"R�̱� ]+8BZ2������������\ܮx��8����� Q"��J��!����B�����T'�K��J\�7�*��_� �	tH�4�_<la4/	�r�oV�1K
~%Dt� �M=����Bq�SങZ�.�|�n�;�Bђ�m���_���n\Z�r&���s�(d�P�`�w�|�w�4�vN�HRwuʊk�:qs\2f�' �G"�|�ɲ"�v&���e���Ků�1�'H�L���Aіe���!���*�?��>caY�P�5��
��׮�}�VV���2�Uix)w�I4vf,����q�'����ZH� 񔛸7�ZS�������<���m�z��Uh�7�Wt��������H������:)�A�k�K���R��~zբ;��չSzg7$r�2�_�Fʏ�"�\���3%�}�f��<��4Ҹ���ܞ��E��彜�a�r��^ ��<�k�3��:�L���]��@�Ti�YI�|� �����g��l��E�S��<�{�p�A��%�3'�Д�NM��`���5�4����F5*Q?*sW$�)cCo6H�U+�6�3!*�� \~?�n����#�M	F��oXz+�i
>�����ͿnT��x�޻��O9�>&ꧾ;��c=�2�����(�qtz�� w�%$|d���4| /H��0,t��=Id�1�6@K������5U+ɺ.|����+��>t
��D�fy�2���S��RP�����k3�M�v�Un{sY[����i�Z����������P��<A�u��`+L-T8��x��4��g�@��u��q�oo2�#@ ��7��0����1���]��=�;�%�dm�5/�q�i�#4�@�#�\�*�� A�
i�(RؒF�s����!��:oYꗚ0(xB�Ɋ������+Y�*�'G���H��F���:�����8H�R�{��Z��a@	�=�z�G	,���/�u�Æ�It�;���v+ށ6��0��&���e�a^}������GXN�q�6�(puUX�����P�*��� ���R<�¥N�=���\
8
ց ��P�J�(n��f�AΟ@�R/iDD@�Q�ZNi����|�����B�5�(B�QlR�W����./�N�_Д����"�H�^���~n=�	�y��h��}������տ(^t�cNBux��wd�#t�쫑���񚁄����#�`�d��d���  YO����U�,��A�'e�/��`P�%g��l1kg:���n������_D*F@'�jF/{F���f[���^�_P}7���ݑ�0`���S�$B�±6Od��&^�r"���!V��@^6�<k���z�`/�!���0\��9aa�l�����S�=��Z%��s>�ZN9ż�4E�Ф��C����I^B.W�P-�q�J�8w��3�A���Gl�O{$��^��Fh������9���ϯk�b� *W�bj}��ʽx��h�w}e��]�>T�IZJ����H�9!����moG#w��v�f���b�!�����J&�Zz�8�L���:��
�a����]��ㅧ?��h�q%�r�`�T��,q����Z��ib�Rڤ*���V���s���433��,�b���Ȑ}�w�i�~3����eU���h0fp�X�M2B��6h?�Rpon����iV�O��h�6������r��~�tY���ݧTn���;2��z�e7_��D;v��3}�:e���������˟�Cp#B�43��`X��2�u;�	O�ʣ�#��M��X�-�>���i�0�Ks쒒`�J=��.xx̆��*�"[N�_��.Z<B-��[1f|�DM���j!�(�RM�	Uh�Ӫ����'�5�~�Fw�R&�D��Z\����N6l�Ulk�|����f�qE��HT�� �b�fW�	Z�%@�w�I������h�Ѕ]��=?��'��V�u|��D���єЙ�]��Y��u��P���c�����aE$2	�pvZ��� �K``ɢq���V!��uO�cT��\A�ϛ1!�����F��O�re�eXH�#���j��d�7�� P��|�Hb����!t�q9y�fP�o��vXR\w��ޘ��T���Y��Άcu�%]��7S�'�l��$��;�z��R�B�����|��a�;�N�Vx�S:���,3�CKT��G�9��s�������p��-�*�s}�B:�:^�/�v�!�K|p��&'�K�-Z�@i�Lh�ˋ��M�h�q���*�[Mv�l�-_[#(�x3�4���
]�o^	�ް�����J�F��P�I�����`E'؞��Ubor���}�������T�W��t�4t@�?E�&v��[�H�I۩L߫�T�Hɑ�˓ZWXF���̿�4Ы`��*e�oє��T� /��24�ۼ���Rb]�{�|\)f��^�#x4��-�JD�wu&�v�H6ap���ޏ"�7�K'y#ߘ��Pa54qqQS��l�"��@$viij�ظr���r�0�I�}����d�0�m��g�P����O�S�����v�j��Hw5������ �b�ώn%������}����W64k`��ܵ����l�>Rq�.�b���O��UL�0f���Z�ζ��)�I=�3+����tg���a�J�>
���cC×�"��g�<'�I74��n�?�K��or�x�XZ���!P�1�����k���zv�t'���޾�"H��M� 䩣���G����@lhm0�Y-Q	N{3C6O��J}\���E0����ڪ�)8U��Li5eU��	�ds��7m����5$)�I宔��'�96@I&׵W7��;�A�T~�c�D�"�\�@p�:��k�]�F���,���j�Z��.t����Y���%M��T���~…���*"K!��m�I O:לe.:�Zr��n&d@���2��Z�S�FKm����DQ�z��,�|&9RyJ����9O�!����,ؼ0��\�A
�J�w
�bsI{ ��_;���7�1S����=�#R�;�2����"�/���.��Pڻ�W��:�㐛���q�"97��Ϗ��G⍤�S��?2+�V���;J�#�Wt�����6��f��36���hl�(VP ��Z�t��&\^SG���<qOܢÃ-a.�p{A��A'�C��gc6�u+,>� �~��9Οp@X�n��(���n[:0$Ɩ���NՅ��$��yuG�s��࠯4B��"��:��u�=e�,Z��9_��*% �?0aG:�E��+[�yq
)`*�Bʹ�1�ۗ���rz���Z"�߷�NE�4�:�':|��o�_�K�Sv�f�P+����t��NбB��w.eBI?��h�Y����n�}�:\|��HV�����ht���C4x%�p'?2Y!'|f�q;�^�H�<�O+�?����g���ޜǶP��b� ��a��넣��[�̠������u<�G��'<j�VK��|��M�s�;���IO�m�x����EPr_���Q�X}�m��b߂�S�
��:��f���f�1K~� d��9_�3:�r>�'L��&n_t���a�e�ŽC j�5성�n �r����.}�c�����+,�Wbf�D#(b�7ϧ�v�~�9#���[x��X��J�3J��S���a),�������(����c����G��O%x����V�g�A��/�GS�są{C�c0��e�M����"��oM�(������+X�\>�_�0�T[0�/��Ŧ>���l��ĒN=yD��{�0��{N�����]3�F�!*��F���w�&} ~�DWH�v�?wҸA�Q�'��7�Krf?r�U�d�ݿ�i����d,6Y�a+��Sp�E=n�����&+�5��i�{�B��?d-���^���=�s�{B{�e]�TM�����gb�*���0ٱ'������#ml�w��3J'�4�BX����I�#�AD�@�����e���j��Y�A>{	+PČ��+Ul������P1L	:d�2���]E&�l��Fe���� �l��>%�:hSX"L��,9AlP���#pO⶛�3�cI�!q<����T�X5�{l܍����N O:��S)<<�:������{Y��~�����l�xSbӣ�F	W��e��Y�-�z�w�3�PX-��Mz�b��?�},��c��x5�~�Be�o�cT�Z�$I�]}�ɇ�{��v?��^&Vy��߷���Z�*�9��2W��̷x.�Đak�`�Z�z%Ǻ	�����³�uaBPׯ: �L���'@�q��u#��QWb�+�l�N*�+�
	������nE���¸���Uk��:穱�4*3���,�;�pa]��-%?kZ�6�3�+q7���Ŭ�<N!���ؒ�|A�f'�@֕�����2d?r����F�@�Y�������TfH���O��P��i~`V����ծ��^�x��Aժ#uX�7��~��Q���������<�h=/x$y\ҿG�,����nV�;jx拝@Ι��3��n�d���֛��M<d���iZ�0R��]�z�Od2���&k�����\����8�Ի=�ݷ_C���d�u��m�j"�����K�]Xk��PU�M#��<��p�{3b�B1:�����?1=N+T3��m����#L�ԍ�ٷ�U��+��{P�wҫ�G�'�׺�z]i���g��,$��}38��Ns���Ѡ�j���(M�(���� ����?�.i��́OL������	*Jك^�:T�+X� s@4�];�Hq�a��z��O�n���W���}*���OC��PH$)v�=�٫#4��>��7�p��tr�x|D��y�����(Y�^�
[z/���ހ
�ETލZD3�C:}ҹ����ɏ��;�t1̈́����P�&���y��B� �U븼��_�q]�U�l�ljFh_�ꇹ()�&��3W��'�Cs��SJ���$ ��XW���|�j#C������I*�#9qh�_�L{�>ѐ�B\��#}f�*�p��m55h��9[�����	������a�QCe�33b�ȸ�-`K�m=�օ��R��ciUXA�gͽ`+a�Н+�a��j���[ixr P�a{�x�t�~�(��^5�bY����ky;BNA�M:�Fp�d<�;�.��>g/#�((�d�8\�_4����2/�&pv�d��p ���g�C�ȷ�U�gY�J�bڥC�B�G�*w��9�3�!�x���p�����޳���Rh�Cp�����^�l�ڜ&���0�W�����W?!Vi�K����R�|�+��&3#��~8g�S <�EC0�؋4c���0��L���>ZP7��������N5 '��{m�0jR�02_5���j狰�����8����zW��kzJY!O��OS�b����~|�Ԯ\}�񨫎L��
���)�����a
=�&��d�i��4_l���R������AsoZ�Ж$�g��+�[�%j�*���`��I=O��l~�ݞ�ɧ4�MB���`k�1���0sun_���z֌�l���7���v� r+AhT�1өP���C���3��i:n8��C�i=�-`�R�Gz�\+�H'Z�+/Bj-Im����	�|x�����B\�"������j�_@��x
"fu-1C$�rZ�%�y������ܢ̋(��ɢZ�Ѿ�����:K�<6�m\�0��Jܭ:�9�2��^��g�uL���e��jn��<��f�%���\�k~��0���4��sY���U=���.tPݺ4@��6�_p�n�6Ra��!t���V���h1����6��ΰ0��W��<�uQF�sl Ru�#A���e���4&v��ͩ������>:���Qd�ڱ��K�܊��������ܐY[Lǚ<Gk)�r)��L�`���1X�Va�C�f���I�Z"e���!6)��<���Sշ�U�O-?_���,_��f�8�"�ѡe�^)U*
R�{����ϝ�;qc�S��
h�a�9�
����ģj��9`�*[�4i�b/4��:l���]E���*B�@�~�y]�'�~��V|��u��|!V��h�6��S�K�}���_D��M��_	��L|t�/ˣA1B�9��5pP�F*�}�ܳhָ1�E�ս�d�ʻ�A1��(2s��a,���Ԇ6�4|��󕲛��e�������>��e��-�)IÊ.e3= ���������y%��"o ��o+���\Mzщ��#�WPN����\:+���n�"��=�]�"�t1m��ŝo����aa8j�R��vڒ|"✰DcVE����Z�å:�^�|�<#�>�-"�a�O5��=J:y�Ά���kv��j���YF��T��LsG+y��%���[��b8Es`F��1D�Ϊ
r���sn���[V`4�J��q#�D6w� @��� s�?�@0�j������_7���-���cF���$	4{ڼ{�d�hq< �D���-��P���z��!.�+ND�׺�ֳ���X2:�z�^QS�@@oP�V�tG,�3�>����y���Db%^�Z�ʥ�w'��dj�����VT_6}p��6|JZ��}hv,��޴����Eŵ�r��!C׸�D�/u�|�s^�H���rg��בy(')@�$P܌b�"6��\cd���T� 2I����y3@�<
il�,r[`��¼�ܛr[W���n?O��օ�\�!��H-fG��]P�����AbX��\~e��y�W��6g�#�0�I���j�>a��%�ܐX�j�?kaΌ��>����%��� x| !���~��&!�Jo��ܵ$�
���h���m�[�O��g⃳;�ѿh5�88�Φ��O����ѽ�!��&`	(&�
���sxB�
�+9Ut�w�����j�8���-w�J�n�i�7v�-e'���Çx������ީ�a��a�E��t�)Y^��c[ղ�{zaH��-�ّEd�8pq��/�4}�&kq���(ƫI*,do%җ�V�9b�(��:f�Th~"�<�/�[��4}�w��v[��W+t��Vo���/��5󕢦W�-`�/�"<�j^b'E�K�:�`ٔin��R^ZyV��:�e��mARf�Ɓg��R������/���0��G�DB�ҒKᱦQ�g���K����.��2����� o��^x(
r���Nn稇6l�����!!��!��Q��#Hٲ]!����0RG�V�i:e"	'���&��W��`���,�_���"e?�����[�� ��F���myͽ��8M�D�,�ЮR��X���?��� p!�snA�`_[���%fy��$��Ei��x�\�|�Ȑl�-�_�n�xĸP?��ozj����<G��9&i�eƖ%�fs��6��¦QѤ������-NF�|�$�NkG8H]CG��f��I���d>��d6�A贷(�,O�ze6�%�*��zhok?�X#���!�2����l2c�r�\�u�\�a\�,���/�T��d(�C��W���/�.7`. ��N�{:��/��l.&q���9dL�K�~h���z�s�FL&���:�$��"�߅)�p�K<c��;�8v^��oD����ș4F!?�M�x�Oҿ��q��P�`��c�E��X�\�;6���Alos$L3����_�e
N���ǂ��I��g�'}q��N�)/l�O��,":N�}�s)������;y'mJ��>�ې��r~u�]8���G��:�:�=���I��F5�n,&��*�1ue�B����Z�X\�4���5`���z�N���fD����Q]I�z"/^-@҆$�u�x[E ���p��v�G��Ϥ;s�k)>W�/2�8	V�v�k�RTxR��� �f������ gl�"*غ�V�F.Ld�}z{(S���y����z�1����,��P����j�A~���굡*BM��U���I��)Ʊ��nW����u���������j �|�����bϽ��+:6�e.�BQ��B�>0����bt���TN���0���ٸ-��b��\�G���Q�)�����p��5v"Jґg��c�Zt��"���yIw�ׂe/���t�T���s�6��L�
q�����!F@cV٭�&��D�>��ˆ�y~*H�42V���=?�M#����!���J�q
���o�*M�T�X��=^�jr=�Fݽ�$�*b:1�C��.ޤ"��B0�s�}`��u>�J�
�
�N�hΰ�"+� E*��u\��cKv�5&S�F��	�	G�5���10���3}�H�/C�H.i�?j��22_�:\mH�� �ý�L�Ύ{\D����$!S�ؘ|�E���F�T��Ĉ7Z��`&,�D�ż#���)��4@���f�[m����'j≗%�D9�큩�ʢi��/q~�m(VL։Wf�[��&�ڲk�j���W�����a9�֎D4"�A[��cJtaO����Ѭ���̹��]Ǧ�NƱJg��n=\I��J��q�s��P�D�a�"�)L�ֲMl�5�?�5�+�M�L�gm��v���pF���yQ��NKs�=trp��Z�ɫ�*�b���f��@EzZѝ��`���D[� U"���JM;�a��5
���\EY��Q���������í�F� �3?�p����8]۫o^�|I�sX��ߘw�XMjJƙ��H��s�M�)��١�Jk��JЪ��uϡ5z�Ʃگ?�;[(& ,�&r牖�u/O�Z����N��e+3;_{EfK��h��.&6T��(3?x��5Xf���x��]��k�~���)�(L�`�V �1,it~�t��;�w�0�e%L�/�ز����fE>������h ��%�ܙ]ӺD���~��5\�>#��iy�Z�s�.Ƈ	���3��
nH��gUc��V��*^eo&@&�aQ�>em���=�p��B�E��?}	�zx����}��77}�Yh���Ѱm��ED���б�֢iX��oV�d��Ix��;��w���ԭ�G�aϧ���L�m��6��5�ž��o�D��0���68ח�#}��tq���۫����R�p�M=#���?zz�8�=+�T!��,�<���s�G!qIɖ��V����?�2Z���|��u��1׏fkd|*��}~]w�����b�hZj����Oc�p8SQ���|��}戼\/��iy�4�U�S�?!�u�/��*|�mA�	��J��[T��^7��M[�`�,��]I�{%u1l�ev�ߌ�=I��t� ���������t��J~/�>Vv�]Ro�u;��jo�a���c�ʶ��B�����g׹>����ʓ�����IG������`�r�NI A��ė)r�,�^}hn�e<�\4�=D!Eja�b� ^PƳNn.��s�X$��� �K��|�H7�*n�
��!�1�vU�h���:Q<���������1]��<P�DR���=� �FL:���]���XV�q�	`۞FV	`��8��F}$Y���`�\� &ǅ����59��o���^��U��HU!�����������(������I����gr��F�n�B�=��\Y�P�P��"G.�2�;M��~�ZB�Qc�Z�fG���i��bx+�@±�
�1g/;7�zڌ�⡑���Y�:���<��"������qQ�e��K�s!! ��Y�*����M��4S#/��~��u_mY�Jw�	6�ÿaZkf�'=9�˳���E��]Ҙ�AQQE����B��%��r��Sj�Y�c�?0�ٽ�]��٣�[�*�e���.kI�sH:�D����m�0Dx�X9Qs ��P�=6�*��Ev5�k�a�� kۃ��W^����#�KR�R����*��aF�2�s�.���g1p�ʚo�W0dp�On���-\D� �֙��/�1��k���8j ��a�5[K��O�DK �o��>���#=�p0�����H���U*��=Z_�:���Ze��H����z#��f�3�<V]Ә��d��*)�	��V�0o�<G��i-�����F�t������[��~�`�n����*ba,�
�ސG��*���P�ɹ~��W��%���j.��t�C]R<N&��h��.>��`p��ס��O�18'LWK��}�HL��A ���Fi.]�g[�D�n�w�l�ay�NkHۗf���'�	�]5��8�Il�z�TY���'3��� �v�}���^���w�����6�O�?+�9��8Y�����o\5����y��n�F}ֿ%�����Ÿ�����4�ڑb��.�}�̶S.T�:6��g��5�|�� ��H��1��W樱��H��*�(�;���\�YyB5S:ͩU�AKz���������'K,nJ�uU�b�������Mm�K�`afX4��	S2�R�)M>
�J�E��Ǫ
*R�ࢨ��:�(V�}_��e����G�q_X��+�Ӧ`�����;��`�V� �t�*�&`�5G������1�~_�����a;�X@��{R�\b-�Vk���Ճ9����#SՈ��'w1�I0«���-ଭ?]�?�H:^���L#c܇%-9 ������>t [U�'Xk9��+f�*L����ܐ�(���X�U��O���F�k�gb������SR�#(�pI(o��{$K����`��IٯEy�w�v���¥(P"|Aed����,�s��m0x�ٷL�/%�Y�l���H=]q	�h�5�G��'�A�]�����W�����봉�.��1ZMl����	��c���.�+�D��ہ�%+t7��VB%m=�" �9�B�B���2c��x���[�~�x0�:x�0-c�J�J��/\���$��F8�;�r���{��c=��>� �GƮ�-��@��~�46"]V`��OI�����,�D�\���]�`��6>]�G��V\�su[YG1���1C�ز,_�D�H����[ޘ���=l��`���齏��o�{{��e�o�P'_��3[�.eP+���߸d8�Yf��|�Ry(�J^�҅L�S]�M�����UX���22�	��m�dm���f�e"t���M�̈�!
��#��\&�LPԨ��JjR&>X��9���:Z�x,P�t�_����g��_]��*	r�:4��Ӹ�q�B���m���f�윷 6Z�F�iØ�t	�0D�NhMX ����c�����bH�t�0�b�����rQf{&�H���_X��A�_~9�o�ȗA?$A荅��\#�K�	�K-�/�����X��"%Q�sp ��+�K�C@8�B'~��j��P���Y^�]�Z�lHw��xj�L�biެWGk$����;SM�$$�9�����m�����Bټ^�O��eN֬�$QwaX�$��X��&�e=�"�x$\��3{�p@ p`(*�Q@dg-T��F6�Ϟ+Z��G����\���V�j�U�	�as
�޾��j�{X�E��궞R�}����	r�Ք�����4L��\��I��K��>0�7�Ѧ8����F�N�3X�SO�ʢ �`chmz���h�� {M��骄;�eP��B���HK�ڣV@��S4����jS�dE��_H� a�H��TX���$���J�����.��ϋ����F]� ��������Z��	��,Ej�@-e�0?G�yY�*rJ`�)O4���Z\���`E���SN���ާ����Ћ����w��2�&x���_cbaW��y�}^�λ%5��_@�Ϥ��{
a�[��O��d�N��ߪj�tH�3Ŝ�-�k ���	�ӓmĐ����菬</t8<��Y��#�#^�Y}�gZ_8��4y�!Bc ��"`�M�F���VY�}"��_��k/#������֌���If0M���`�?��ع�Y����#��*�q���q4���Q9�:ty�Z��J�b�� Kf������C�}��Mn �	�(��Z�c:'6=c����lE`7Y��
�SeV�"��٣��@�u=����8�[�_uY�M)-D��16c�G�E��1�'�h_��⸟�B8�N_Vk_"��C�|���\lT�y�6T���v3$�.�U}����?�8`4a��Ց�ZM�a�״��
F���r���Ip����nc�c<�k�b����U�njVrK�Ǖ���>+�L�j���z�mU&Y��H��ͭ�w���o�WA�d�՚��'J8'��_-���4��XN+��7
����So���}kT�R�pYM�i"�{T���|��Ҷ#0&s,S�֖��:�+��=.b�ni۽�(,2�� �4��wO���E"c�}rB��+GD*-@L%���o�ehgT�8��ўf#o��q>k��X�q�2�(�9y�RȻ�",��Y
��97��hL������Ǹ�o����v�q$�wtSU�5p^0�Y\��aʑX(��u���P�<���nѼn��t��$Ň���-��2��>w ����k��O�'���@�└�Z��f޷L�S�=Q��;�mP��D�Ar��J���^��8{a�q����oG�<_���#��9,l��3Y��I��5`f��/�!q=�:���k8&�~m�z�G��f�߽Xi�Iwn�$���'1t���@���[7�&�!<S�E�|�阦i>-�8O�Ŋ˵�˻�:k�B�$1u��9�A�,����i�s�E����D�X�E(�K�����������������,M s�kBn�Y8��aCҐg�ߊA�,�Tc���/ww%\L�{~A/@ b�
x���tu���}����X�-�fI��w��l�:es��.$-�����>m~�hopn(.B��N��L���3�3@H�%TyIx��)q�B�1����]�OeK�N�0��ms�.#�f;"ub�w6�?JR�s<�;nE��c~��p�(��0x�"����gQ�Ҋ��͸�pNF��J�(�L����
�̒͸�o���*%����ƕԃk��b:O~�KE�x<t�.l�Q�ܗ���d����:BoZ�5�w'�b����a�w
jHc��*o��i�:Vp��T�Ē��%��J��Z���_�[�1}��_z�ʯ�_cW��;�����a���oKQ\;o�
�z���ƔibJ������9w��1w^% ��iD��xq8�d�K�w�ݿ"���m}`3C�Y,f^v�8D4��u[�7��	��ʃe�z(�z���lD��3�[��q��N՟������=	r-#�٢�>1Ϯ�D �y��u�+E�99��'X��d��eI�cmDG�G�IЂ/�7Bɣ�H$!lw�Gy�3�{�$��Ya	cV!ID5u�������K�*��Ro���
��Ֆ�9��M��Q�_�6G]���_"�#��n��ֿ)�֘�%�rJxS*U�%���gDS�m<��@t0�F���x��y� ���B)�й����>
�%/��z!#���n�TX�˕�x�W���鍳��x�O��ȺF=[r�K�^Q=0n�A󘚠<̰F��� �����l�F� n�U� o�U�l+��Y�15�>��T�h���Gw&�!U�H�1b!@�$#� b1�b�T�-C���ش���!U4�Re?(�f!�xH*+0=m�,��NrTݻ�Y�{c/���AN��oDa^�:�r'�����B�{RH�p��ԧ���&5��X||Q>˞d@ �e��Q|`��(�� j�b0}�;�3��E�<0��F�~��%UWxӜ {��SD��C������XrϓrfHT�u�gi����`Q�4~�(B^`'��5���u��7i�U�c#�%��F�K�_3�,��J����ߥ��z����,3�Q��#@�l	�yR㯋�^���e�2_aj��S ��`I�e�qhȤɩ��k��Qb��hHRN�Ą�Nݙ-��ˬ�Sk(-�+d1o\1[�w�%=���'L%��;n�F�*{N�����>�´89���TƺNVUV0�c�/U�Py?,��J�g�]N����/��Q��h/�ʤ�n�'.UzRd�/.Z�*:X(E�C�Ί#9(�גb�9%�tIx�H�����}���:�k#���m��Xi1����6�/�5\4��77(]'�G��DႬ/���sl�Zt�k:��*/��Z��:�Cج	��,~C*�P��T����nB{CW��k�c���W�8�:_j�е~�񠩃��ܗ{7$!:=����?��wF���$�����}�;�}ǧ�o�U�5ĴҖ����*���b,>.��F}{��A���f�� 
���D󎏫A{pW����)l�*����C�P��Y0:,��¢��ӍQ���0�K���eˁc�÷�b�B��Z�[�*	����Dy���  j��K��q����q���P,\����NY�Ag͂�p�,��O�Q���e�N�	0=hN���F1^�7��}FG%xl&Z:t���mp���:�V��Q�p�<����p��Ț.9tP[��<zL �Wj̺�>�P}/��Ψ�e�sPl)���F��e�Em V���jh/�Q-s��{����T��\��� nӅBB�.�*�C�^�%�K\ɋ5]Ab� cU�o��rC�%5?#�/��a�<o�|�5�&���xP�c����L�*^����s���}����Ͽ��;��"�&�M�v��
Go@A�&��]><pp��7�������W�W���������h���+o�-�G�����{ϱ��DSA��!�ā!�v���8��\?g�pC�bP�i(�Y��"�j�N���Z� Ҽi~��.1��_"�D��c���@�H2a�wP��s�$f������.�`�����"*�$�!�*4f��/}`G�p�+IT��k_��r�k�À�M����{U��*�$�3�F>�)�ڝ�˷ �c0U�B��櫟c"���ִw�f{�K�J��bxq�����HY�����&u�i�Q���j'��i����|�_��Y��ڗ���>�o�yL����H�&���	�8Z���YZ� ���G.d��+ͺ����\_�D���Hsյ�~��F�\��,M6����*p�@�U��ZB>�v~Kqa(z4�/�Ģ��COI�p���{<������S�ys���HfW�ѪS8+�y1�,"$J�"����Q��7�_Ԗ�5C�bgaK���D�ˈn	��B���SB�p�v�co���m���2� "�,~�r~��B���9-�C��0߷|FK��3]y�"�c�85!����F�o8��(ar����s�Sl�	|^�F�|�毵ďJ�Ʀ������Ydf%��,�;Z�EQ�����Ep�s&܄�o)vMR��'�^i �	t�vR6H��E�4bϮ��HLgnB`�h�Sܵ/գZ9�������k:Y��Э��X3�������Y��MGP�T��*t��-k6*�\N���CA(:��.�
N�d�6ힾ���`nlc�X���.r�� �2(��B+"U�6{B $e{�c8�:��SF��u���:61{�J������j���mS���;�S�s�Yĺ�[H_.���e���!����H���P��F����^�ΌW��!k�.�����LD.c�7L5/������ˮ�>�D$/$%�#t�����
^����a�aD/�ܒb�aŦ͚M�����dR�m�	l����b�"�MR��-����ľ+� ��P��K��[E��~������t�����R]|�5C� �v�5�b��
�o����"?���94�Z4n���L�T;�೴��Ȿ�5�1�T��3h��5�Q�ipd�W�7�W������J~.X�3�^hM�,�=U��=�O�{_ЬA��ǹF��1����m��x�@������aS�	F����CLc����Ln�o�8��b��7-{�T�{���WS�ےXS9��%�@���������t	�]�%ܵ��7�?���w9�f��Qߩ~�h̣2Jia�~�{�yT_E.�W�]�L�]�� ��[���wH.j9���c),)V�2�:��z1~��vV��vr�	/��Jd#I��0�T~`�d�Q�
��m��	Z} �P�&_Kl8xX���B��(���\v7�]"^D,3���#��h�ᩈ���r�z�*�E��~?K��8e7	;ǘr���>c!x��_(	}4���W���@�%n�b~1a�:$�ԑڧC�꤀pzqg
�%J"�j��IT�T7G��7<q���b{P�w�m��U�3�͟"�7!��n�_�����xT�*\<J��3���W���Ű�Nw0;�r�;��)!(�il�ɟ	"X�'���/�
�!�4���%fJ M_�����D�"���/���6�8�n9�M��qo�g6��C��F6���T	ܣ��DAT�C�G�K����<x^Bk�r]E�_LHK�<�Tw��I'1o,X�$��؞��?��I�g|X��M�X��}���Ϳ g�mK8YR������ �	@�秤HE�]�:2�rJ~%����?�� ��I���yCl{�Kwǌ�������]q��AQ�mt}S�)KU�3�!�&Q)����4��Ν�OF���N1�Y JN�E1��4���`���e��avQ�Yyӌ�I���NAP�h�@�?�m� o	Z�����#=05�xh�3���$�?�[��9k�
��eC|Wfum氄���n^�tLsx����Cm&ܯ�B=���lO��l�r�j��WW���K*C��C��Ӫ�H)ޘB>Y+R��H�p��)ϗ�,E�į-X��.��2Yy(����fN������5Unw�|L'��U}��v�t�Ł��9uD��3ҏ�[��u���3��V��@�g����锥���ެH�,��k���] *�M��ۘM7��;����[9d.�A/���t�c*�X�Mr%�M�������n�����A��y��f�X㊨g8��{Or��7���>X^�GyG;�Bf\~~�k� l��@�
18\�b9P�n����U�eX%K��,�*h"���C[RX���{��Af��i�Ȩ�"�лJ��e/+W��&Lwnqh~k�"�k8�w��-ݲ�1������N[P�,��A����L`�'s�6
 �A���kv�ksrx�%��*�^c	��"�%��)�G��A�|ۨL 2�bP���|���C�i�h�U�.�Q�o�u[w�/,d�y���P�ϻ䘶ڴ�qN��w�oF��W��h%:�H���F����V�#"[�o�U\�b�Wߒ;�,�<�'v~�6��e��z��˿����dI�@�+(-�XRVu�^��F_�����P�������-_"���I]�-��kh�!��G������'H�.����T�į��r�[t򹕑_��:P:�r����g�Џ�zD��>�,�Tj��
�����ЪB�Mˊ���@���ek=4M�QV`Q:MM)ʕ0�s��@!����_Ƀ���~bB����P�wK"Sޏ.�O�P��Lq���\�ѿ�^�ݤ�LSP�e{���%���yܮ��*�@���igg�^�V�T���bL�fT��z�f#��|�IZͽ���:�G�Pz���lmj��<,�����g����6��ܬ6�ݪR)�Q�H��񿻻��jTw��݄���yd)������<Y��q��N�+��2��ּ��^�5��b�$(���ocV�mͿ��<7�^��XAR��z�"bV 6������Jí���
>�-�_��h�^�h2�eQ�?��5�hR�����0X6�̳���$�K����mj�Sjq�̍W�\xl�AH�-�9'8c�N����MQ�/��KN4	���#�r5�{8Do` w��d�ͥ95��ciY���Y� ��^�լ�p �=���E7p�gxt���N8Ϊ��?��F�6,�s��$R~~�ԚN떌�	S
 Q)eY)�_�}"�)O����a��
�9��E|C�'�2��e�4iX�U��DL"�q��iR���-`V�l��(�0���/\qmDnI-R�/%<�$��*�2<���@b�.VKw�a b�<m`���d�����>%�FT�:��H�?c��zADY?�6_,���}[}2��+`�%��0��Z������1L0Y_$;�P�%��#�`��%I���������z�݀$K����փ@�ް&M��k��^A���NKf|�t' ,�����d`�Æ��/�0�#t���lm*\rQ�Oxp" ����̈́?�G��VM�@\�*�u�÷��
YYbT觡��G ���|�]N�X:}�PMAG�۬[���:�9f��)|�r��8-���P�R<���$W�
�%��D�'�}�!uK�`TTzzc�Q��I��6}�j��Mxoˤ�g�XT9j4H���iob��d��._�eg�"D���i/>�q�hm��s�k$�ǡ��{����0L@L,i�M>�..|E�\DƦ�M�Ň�]�ǥ;����m��	^�ѻ\P�����3�b��DG�(��Ѣ k4��OЗ�ط��O�ߢ�;�
����~�?�]�H��i-f��,�ɞ��Wkf��f��փ�\{��A��q��4Q{�ǉ�����ڍơ��cЖ�)��m�[�A�Ya��ԥ	�4lk II��]�H�ƅ+f��9�x����Y8��������`�;��Dԍ,5�vH[v�7�y��2Q�׳[gƎ�&i�Q�O�ҾY9I:K�vW(HR��z��xM����IH��5"��:�Wi�f�Jhc�6��y�i���q�im����ċq�:d��k��O:���
X�G��%L�U�� q�o���}�W*9$R�<��u3}Ƒ��ӓ��-��[R�5��H=ߊ��q<(27Ek�(� �����B1�5h-�ٗ��ܜ9���q�.���CWZ������6��7^`_}�/��&k� W���W�_��ڱ%U9-Y I��qQ���F��V�]��*l���}>�O�E�d�	�.eb���w�¢��C�A���^�8�aVg�ժ���5��^r�xT7��ғ�M^�X����]o5��zZ�E,Q�x,�r�;�����_�7ңL����zM�[��+����L����O6
�SV�ޑ��=�O�mx(,�ם�4U���O�C)ntm��]��o9���ژ��%�dMhjiᩜ>+���6�K���ݥO+���c e)8\L�>J[H.����̈B�gB�KY����{>�9�GY��4�a~/�|v�m�2����sg'}*�=�G�y�@��i�.����b�z�T)�`��ʍ@�)�^����߇�hC]8�7�$��ڃ?�r|�JP�fA��!z'fXt&L����h�����(��<^X�P�+hs`k
Է�nN��Uo�7�'��?��/�#�1`Ā��b��:�P���i5���/�7I�ίl�@�w�,�adX�[�����N?{6 ��Y�5�! �r������]��,�¯���=�2��P�އeu��*4�Lc_ٵ�"�_����E��!��0-�������*�K�'�؈�tux@G�b������ȋ��y�W����[j*�U�#�R@�$�?��B�Q�!�w�E)0�S5y����!P:��\�m�QY��R�U;@��9�N�8 m�`����y�c*���H2.�����!,� i�u`G9�%CS����NY���Z6t�R��}��:M;�u(�?q"B9�$�a��R�[�"',��b���҇��5�T�S@��p����]���I٫�gBZ�'��,E�Į3���ם�L�0���W�2Z�ip70�h���n��"�$'��ftQŷ��ջ|=��|�b�J�_��N��;����a�!|�� \����d�8��@=&�7�	���k�l�����2���y�c�WU�X睘��#!t�ъM�b��ڼ�i���-Y3�-IY��
^pεR�������\�+(��N�f8�č�=�^�2	�@��3���_ă�yƵEe��l�B������u�
+ŉ#�<e� �Gz}z��x�b�j�kR�kd�s��lB�(:�Ɗ�=���(TF���3�|dx��5Mf�A��E�>��(�-��M���j�$j.����#�Ftvb�u�q�_�_����s�L�y��^�Q��D?7�*f�-@��K����N��&��FZ���y�+C����O�m�C�,6�	�6}x���D��kc1�����?�vG���n�(��Z� &PH>
A>6�����&�Zj�܌��o��������s�����🏿wU=�(%'%	?1�n.ox����4�RC�|%��I~Jaiv�VY�� ����ѠW��R�ʃ�v�m�4v�����(o��ʘ��N�{*X`I�(��9�U1�9�*E��@�$�&���Q/����ւ��/ `WS���+m���V�ŽzH�� xÊjn�ve�e����)��H�D�Kn,�o�NI�޺$��"��h۩��Y���;�Rqá�c�c(�qT�1Bqt��GK,ƬTra��dĄ;�������òд����=)��ũgVS��
��^�]�Q�h�h��� � ������-n�TWy�K�^�@���%-L��`s�
��|k�bv�'ue��+����cJ�¸�}R��:�.)�7Mճ.�O�.K���[|�ڊ�ʻ+���'�P���O����\���0���Y���F��%��HT�3�}�7K�/��'�ɡR[�VRl�B�R!2iB����nS,Ϛ��u��!m� Y�X���5XβE�9���B�/&^>Ǡ]���yኢ���=�d�&�*g�����A��t?"��|I����h_xPX*\�̯p��8d�QV�3v�z�X5���U oJ�k��@�US�������U���çxg������T��XgK�=�e���^q����:02<R���Sn�F��������*igM���mwwknJ�Ւ�����W�Y֪�"�4�B�1|���Z����!!��3��o=	�����+-L���pw��;�}K1����p}�;�d��]pE��d��9�_M������٧"|+_Kh�Uįq'>st�~�m�-'�{')`��[�e� 3XJ�������d|�:�g���s�,��j���(�A1��ro��b]�r��x�N0g^	V/
>'bzC���F������D(r�q���*/Lx❫�����8?����
h˄h�%#�kă���ĀC����7U�n�MKM*�$�w���u.8�f��NP:�GȀ`5����_V�_�i�I8ֵ�*M K*e�ofܻ����B4j0��"��Yo��������:��%�5��8Q��/��uc��s�c�HQ�Ia��b�n$V�[�CR=C���<���8�K}�肚r�Ф �Uq�8Ug��zo�C�O�Q���QfX�@`�����b=���9�;�2���8�YKQ&/��|�>�Y������ \�<s(6�ʝ
D������3�V}��J�#���y�DIGZJL\��.�*n�3��rb4�fw�Bb���0Q A��l0M�I�q�~@ppЁ�i��t2f��G�IuѾH��5G9b��hB}�E��ƪL���8����AR���_�����@@x�
a�"VH|�3��V���B�ʕ|�v��A�ퟷ5�ެtXU����Rn,̤|ehڢ�&�Y��5/�^;7֧a��^�xb3oK$�*#mЎ8'�r7�9��P%sHX���1�\������If'{�1�w{TFYA@&Y�����a�]�l+n�j_��^K� 	
��ܩ�3�U�w!�L���8�0terj�l+���ݤTà?ˌ��OYw���,؄f���O&&���,�C�M���m:�&���ń�ܕ*���z��m��/���a�m�=�!F����R=Y�O���|=��SWy2Ij ����]F��N�5��,�d	�A��?�u�ߵ��3�$g��;m��J
.�g0y�X|��x�^u�"ql�]G�Pu�2�*7q��&��y�*�)b�����Z�Y��}v��G�����Ϻ�z<��7�C\�ʥ���fc�X�Sn��P�ԶA�#;:��x��ᾺG#$h��{"��d�?9F:�p.���T���Hh��ղ(3�=٨��Q!<��]aBv2���77����az���iD�i��y�}��q�[g��d�QM�d�ѱF��ߟ 0���ڱ�����"��,<�i-�/d&m�rm�OH�����;�'����_xje������ۃ���C��T���Of�4�m�y �Cݞtv|r�Qw��;�����s�����8/D"q�&����aɔ������ l�̒�K��MU��Mj]sX�%X'�	[��V �ā���	ػ�Oڀ6���8�k]����Q�"ؙ���g��K&c@���*�Z�/�[n$���c��c\\�֧{#3|� zoC#���<�4x`m����{]�M�j��#\Qu��Z,��c���ƛ�Cs���R���X�Eq���Q;����VB�t��*ͪ�`O�ѣ�f�Ȋ�@�\]}��D�����B)L5��%���I����2lں��P�f�(7�oN���f�T5�Q���re<PG��h4�*!�D(7ɳ��/����n�D��j�.ٛ��C�sS �Z�d��g��!Y����9�[9㰅B^/x�
d�2f3���Lcp��ȜN�t�Q{"�V�9yD�ha��Y��N��g�p8��)(x=��~�dG{wT Z	��F8�0B����G+�fؤ���Qn+�,��Ї7�Gһ�AE�<���	�F�8�Pr�����$�z���wT�~!��j��`��&J�����r�8�W0׸a���/��:��Gy/�k���:~T�7�u'�+���S��|םQ��s��~�i�X�$�r��_¬��{���&V\;47��#g�Ą�D����sWhYI,/�i�@�'��[�Bf����6e{��	Ю�E�Cf5)�x��
:�5Rχjc�����fv	���f��c�(���d�'-��5 �v6,���Gz|~���r�/����v��h�pw��RUQ;���K�78K��(���+��ϛ�����zw����E-���)i-��PZ���^�7�9r�j�3_��C�Z!��
����w��j�.��D
rzvj3L�x��j�&�[Rs��3�*0FZFs*���7�@B�b7����T��Q<(���V�&��'iu�ԏ���;}�`c
���؉=pj�)��\�"I�άr�%~5Jt��*��O���)���u�2C��G�{P�M |�<⺫��Zͣ�5�G�e�b5��`}��s�m���#��.	�)�C��7歎
&��	�;A	���3�1�D�a�9W�Kr�)����vw�KJv�O�.T��تp5�V��e��~�������G'����sgY8�D��B�t�$��u�cB��pL��q��i�5w�c��l[��䊐�V,p���ɶ���8���j��*>��WQ�>�$�c��Fg���j��s�S�"�F��~U*�8v3���v��%�5�ڸ�Rǔ0�`!���^��9@I���� h=��
���Uh`�+�	و�
eIM���Jv�q�����s���u������ M�P`��="6��&�	�Iʦ���z�}k��8)'����ɛa���}�ؓ���.�����"O�X�Jر����s?�
h�|�L�P���D������"��N���0<�5��m��Z�Q�15�eo)�W��ƚbI�ɀq��Gky��Dm�z��O�:ayi���}�l N�|b��v�R��ԽQ���X�ES���K1��C�j�7>�딟=n{�����_w���� ��>��N��;�����42�x�-��G�`��@MB$��ƞX��/V�_hc!��w<Wun�Ad}o�:�*-日��@Д9�Гy�M����2F�Ѹh��Z�I�@=�-6�xHn?_w��[��!,%�-sn� 3'ߍ5�4�k�xٙ `C4��U/	����3����T�L�c���`����K����jM�� �P3�2 ���n����i��d�'n?L�+������ꭖ���I���SyC~�I J�_-v %�
�}��M��m#�%��^H :���ɪKt�t�ɸ��Q��a#z�ߺ�_���G�E�� d�������$Y<�����xy�:/fn�R�*�X�M���+OYz'�skh���>��^>g�C�?+D����h!�@/n�pW�,}=��%�-����
��o�7W��#5֜$@'Sh~"<��e^�彶�G-$��K�AR>���0l��/�gP�f�=���P�%���%�1P������F�_��t�4�
B�Um���e(�X���M.I��Z�&�S�U&���x�g��i�|I�� I�ͬ���ݻa��S7�ϗ_����w���4��\ﭜ�Ӳ���pB7p��BI��{�ߴ��R�[�)RH$9{��{=���$��}�����+9�ԁ����%��LE��i���n�����.��/ݾt��!W�@��+�����o���\��5��W��MM���tG�V.̜���)><����a]ϙs=�'}�o�q�
��q)P��Î��h�SL(�Æ�3�eŁ�����`�k����d��V��K���#63��&.�՟-+����Z���4�U�ʌ��\��E}�;A�FO�Y#Ѱ�z,dJ��+��6�e���K��(Q7��9�s��JC�{��R¾0����d�-Te��S��X�{���y��د�qq˓��֑��uY�vt�Ud����g����񇗅 Ob��e> �B@�WӣI��fXҎ8:�G��~�����`��@ �-2�Z[	�Zr?�����	�v��o��R�֭���""]s����߈H�~�Nf�iyݲ&=�`��¿f��ͳBLj_�W7���CŊ@�&�};53���Y���=/�i%Ӹ�<�$���]���#}[Ђ�9���?b�4d�Y��_m�RK(�c�&W�%���S�O��@M��J��}��ѱj��	�T�|�8��g������ѻ�DF�Z�H�D�v���r���x��NeȘ|�#8N#�y�|�'��I��3��mv��Ҙ����S�]]�%5�Fv^��C��DJ�3p�����k�O�
b�sh0����ws�d���P+�7�O+J8M��a�OE�述��Y��"�?�a�����sw��B)���:����Y��L �'��c���e�&�N4H�d�qV,x��Bi*Z?w��X��;��0}i�5K?65r��=�!������Y�\${������Z1=�f7�dgS��Sj��_H�Op��<��qkB��G3C̟����Y*�@ ���K#�
a�#yk�X��������I�����#�0�����/ʲ!�j�13���PPR�~�T1lukQ��	@�9�C`^\b���#������ �`�x����+���[�>}�X@��k~��1��kA�5�B�2w;J���E}++5�Wv��>c����}s�e�[Z���Ά9�����b�j^�� �^}ke_�Q��5�{ g�e&�����5��-���=:#\��t������I�V��-��me�2&���l�<c�m�6�Vf�""7B�T��f�[���Y��/q��+A)����8m�?�?�q��wb��ȥ��]��,��E�t�qr����-�,�#:���5��N/iE�nt��K��O_Pmb)|@E�b�,�p��L��+���$X1��s���;��m'��s��L<fs��Y���U����k�ũ�KO�e��"K�=p_n�J��6j�ǉ<��	 w�����hM�d9��=�r��ޜ���o���^��+�-�:���ǳ�#ߥg��H��X���[�<�ǧ��H4׋a��eB��A�F�� ܈�F�����%�-��P )9�2�^�iN�Ǣ�
"�% C�#��LTe�i�&�{�S�tkvگ�c� N�۩���U)�+Vj1)�&����-�W~1��0�#�7�RVMJ����`��[��_��g���_U��Y]�W��d�.fݲ�v�؁͓E�'��Eh�Y���[�k�G;�&zdbx7话N���=�#>��E0�ƶ�V�+Sg��mw�٦a��1*����a���*<�u���=�9�y} ����"x�R-d){��fh��j@���}�w��N���?����F!��V3�#�RUb�0G���ӫ�F�L8���Ι�o�:��&#\ݕy���*�J	l���\�eYp+.�#��\%8y����b~�L� %����7~4�A�[א��v*9�?��˖�f_�/=�:�㢐(5���+��FY#q�'W>A���P���H�b���e'k�g&-k���W*�+�c�im�V��D�|8�ۧ&��o�Үs�����@�\l�|9���&�G���F]V�y1����@0�
���/��I��3Cf������2��Q�W�!Tt����]
�����W`ķP�&"e\��� x�ﳕ�0�搬�=G^�qW{�.�[P��DT:�x��M��z���g�O���7�%�����!��^���S4�ޟʘ��.�{�Ė�b��L;~��8d�ijڟ�ggr=h���|�&&�r��$��H�} ��x����`��f�Ri_Ϊ�qڨ`q��\ЫI|y�u��p�B0<[�v3[b�S�A�Xu{���K���l�;K8]�����5I��Z�v*�<4(��7䰁Y�E�X`����RV�����,��J\��n��k�I7$��dV�D�A4ަ���[���NrL�X5x���@�M1/�+n
!�J]�R��?��$�S��U!-���I�έ���7�����g�,�h6q I����"�Α���A�J�Z(�cszk�8ˀ��