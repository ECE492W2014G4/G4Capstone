��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�"��F9s�`&���a�oq���F�g�O�]�<ݲ����eCL��D���{�5��8̝DFI��Zp\m|Q��
�}�6C���UnF:<�jΈ�2�����<����sf�k��,jڙ�����2��X��Ss�HL��	�������+g?���N�Ż�����|�v7�{M��VNB
��Rs�゙�Ld\��X�'��R :�J���^�����kMkx�Q���3!P}�e���Z�Y?.�U{�RP	�)��lI{tI(S
7ZF���	G����j%F}lI0DzG��������u�u���n\�pX�2PV.x����x;�ʯ֗k�����a*d�X�"�Aj\ϧ���r��$S�a-�������8U���W�Oq�(	&��J=�+^��M�ڙVba�آ���b\���T��h�Ng5���uN�k���	*C��VN�v7T�uGv�̝���?��뾓������]��}��q��Y������r�qѵ�2Yơ�\�i�vr``9]�*ս�X�D �=������o-������
��!� Z����+�����a��>�aN�غW]XV���0'�a�H�ohm^�ѬL��+ۣM�����A�c�ܼ�/g����O��/��Ƽ(e��={��VwS�2XR�$yn�y]^�9�mbu������d5�H�l����{��?/x�к����&�Sr�m���42I�u|��k~w�qR�`�a���C���pskK���`˅�[q�KҦ�*e�\��@w�<�XV��l��B���hlnf��/�׌3�T�E=Gj�@����������x=؞��J2m��!�/8B�"��%mn�{3�":!?͡�,�0e�[���bo��
{ðs�o䬦��L����2ǋ��Z�x0T��e�0��7O�ɐ�'5G�s�V&�塕+)&N���=�g#�y|��ffNĝ)�$	�f�
<�4���U�!k�ʇ�j1"�o�V����R�7?� �KUk��ڀ����y�x�O��N8��'piZ�ː�J,��IH
�	�&��;4�\@Z��١q= �-fw��f�<γ�ߕN�s�3��趿���#j����u�L�J�����4���5r��Em�]��^^�]����|2�OJm������K���\��M�V9�t���E��!
�aFJ�@�t�C����z��g�[KnH���KS�є�5 W�G�=b+�]�r>s�s���ϠA�������Ʌ�-iR|��|ʤ�dg�v��x��5r�m�.��[4Bٵ�-q��-��{��u�2�7�%�)�S�}y�r8@t^J���\Y�ZE����4$M�[{C�Ⓙ:�������}��s~k 8�b�L2M[���B��i_���z��^��e��j�Լ��gEҲ�=vmk()1��*�@ơ��/!_�*� v��� ^�	|hԼ��k! �I+)6�#:k����Mv�O�����р����/��,��)Bӥ�~����X�����h!F�\K�a�d���\WG�n?�.{�M���R�'N;rR��U�8u����d�n(��>n�)�p;}��u�"�]9�&_�8Z �r���8���<�}�����5��H^��W���=Z�:�Z�1J厬	>x��-%M}�|"�~�5q�tB�C(+�]m�&K7d#�>��A4���E^�cn�h���rᚙUu�+�0�X���E��m�ZtuN�75�5�76&W��w�����Ę���2rW�C���Ԫ�^.v ��ʶ��B����^�������e��Ѿ�2	>�h;͂��H#Y��ϔF }�Z��<�|p��֋������K��vY���K�'m����Z�o>㞁��[E7Y(� a���@ͱ/�}t-��F�w�7������h/�5�a��9���ͨ��e���������2�,
���a4A��W^����׎}٬r�$�A��i��6���kF�����	����:��g��`֔�|<�Rsb�p���5��]}�0K���y)����(|�۶�0vU�k��Q���J:ʩNǅ�r�Ɗ�~@�q�[�d.|Q��p��9��5�OHP�esX5�+���Qu.K��쏖�R���-o��6�\�ԟ�Z���������ڳ��U=�k���|׻��o��>kk	ޘ����U�g����ӫm�8��ϕQ������;@�Mӟ�c�oH�3�zb���X��u��+@Bө�!��	�����2�4�����$>�L�
��*E&u��^�(�l��i����u@�
���WuO��K��*X��<d2.����D0eM^���n��M�)��D��9��5fp�=ċz~�����n2X(�KTP*~-e��&>�sS����+��J��x�Xz�<잢�Mvgݛ�xuO��A�F⥗�����';$���~�ʫ��B= \��ԏIa�ލ�Zb�"3Ͼ@Xn�NF�J�
�����kDɍ�)��K�xq/P1��.�;$������� �b�U�]b�%��l����#�����m=����-��[����S���Sc�,�p*g�J��@A�8H0��Ty����gZ%�#���?�"�� �,�u�+nS����Ȓ���I6�f��ܤI� �f�!0@��չ�Rٯc��'�7��٨>+9G�2+ٟyL���ag�_]��[ +~���p��5���2B|�`A��΋�}$�1������1(fM؎*,4;�A��|��q�;.֝�aP�)20n.� G\OGbx]��!����;�$n�͝�����m�#1��vv�$�E�Lٍّ��j��Ti=ښ.'O�r!M����{5z)岰����(��$��{ ��5md��C> $���=:3�����ԙ�b�����v�âM�Gb�.C����!�`��5z�A�qw���l/��}����S����s$��m�a`@��U{0����	�-��� �]�^��G���2� ֭�<�Ӈx�Pzaϳ��{C`��j�,$��W�'tN���|=a����Hq����U���{q� ��ч�x$�*��bdN+D�-��º�9�{}>SY�E�+	)e�jk��1Ǟ�l(~���q��	6��h�3��fz:�R�|�}v��K���˖_��������l�
7�#P�Ӱ��4l4w}՟�ϩ���Iz(��ȸ���Ѥ���vts�̙w>�ı�T䯙�$j���YÁ��ge=q�Ѫ�O��).�Y�:�Q�3Ϲ1��;�*���x�Y(�[�`�A �(w��$��o�Γ,h�@,i��P87Rmt�y-2�C�B�KB��@`�����>�[s����_�b\1��}�_��SљY~/��i�ޢ
�T<���E�N.�2I�2s������2O~I�]#��#�Ͽ�Z�&lC�_�Q�v��x��%5u�;;� 0�,z�!ݿkV�K�fF���N& 	�겤���?2�^��B�OZ���s�q�Kj��ɷ(X�2EX?���ecF�Z�H����JS���F���q�q�cBeV���$��G��b˧�#���X�K��>��A|ɇ���A�s��5hB佚�jf(�����?3o��mP(9��&���������\Mѡo3.ьq 
���T�3�Q"���0�C�����Y���|6�c��J
/r\\���u9�V���S?�JN��Kmda�''������^�x����d?��Yk�b��] �n��ub�:��~�k���F�EU��ޓ?��W����2Lj�A��������"F���b��X	���.I�͛����ޏLMu��iE�m�Mdz&d� �z��{�C����F�ic>�o����⣘!w���{m����9$�d�ٙ�~�@�Fg�o�"sr�W�90���H��� ���"�B�o��ףç�����_�p���5=
`>FV����e(\��*1��8���r�2)�ήW5��������������������#��"�,ӽ?,��c�+O�D���qx�Ϯ��D�<��@��?H����ր@rM"��7%ml����Rx>��s\k,PVO���4 (,p����/#7Ky���m�ʦ&�V���uD���|��X�[�5�>�>ڳ�)Ŵ
�O�>54��gqr�
��[M6��m+�D�+�m��{�N=Iʹ&G�-hz�1���Shx5?��c�7  �=?*H�ƴ�*]w�ik������4�Q�&m��=��ҁ*$�a�,��6*o<ɛ�@}G�(F����	e��N�vBS@B����z����8��:��WHm�"�3_Ԣ�'�/�U4'H�r����Q��3a3#�i Q%k�����������ba��_�G*�������W��Ё��m$7.��c���3��a2DGf��C�5u�vX�f�+�p8!����r���1nf�3���5����ߙ3Tp�̈́ϑB����z�� !��x�Ζ���D�;u����b����>~tI~(��D���Qy*��x^p�u��o:�6��Բ2����_��Q�7��ռ�,�>���R�9 ���Y!v]l���!S=�M�!YlI�kh#���Jb�OK�[�z�,J��t�j�ݐ�y��ivE�\���#�$ d�3/7�}���N������=|Gݯ���1�!��/��i�S԰`�P�;Np㚈�*�"�sg��|e�w�~�����M�~Y��Sm_9N��U��b��3��~�����_!~�����ܔfګ@�ԕR^X�D��Ȥ�	0������̹6g>�����o�U�>��v��.l����U��2x*�t|-�n(r �PG�],�_;ؽը
l��A0����ĔǾ[�2�ާp��=1(>
mYJ|(T���+{�ًƇ!z�8Lv��h5mVq�¨/��1Y�7��|�^�'R�+�k�ǆ��#Y�p����́�����(sŠ��s�9v�nVɨ���E�]?�6�����]x��&
c-�p�d��dIr�_O�nP�Őh�--у�����al����,�洽a������|ߊ����0ӳ`�#'|F[(�N�l��j�,�N�*^��Y;[ח��^
�=骙������ %��X�����ͣ��ʄ�&��
��c���䧥<Q���*��<k4P�	1(��<�&���l[�^�󿵑�Y�]D]�92��ɵ5�*��[�X	�`z�MFc}\ �9��T�-<�1�B��*�υ&_�ļϖ��h�!�2��cp��z$ep��g�X�8!�|ol���Kp���8H��Q����[+� ��G.�Ԍ�i6��
� �=��Il&v��ݛHE�cP�R�.p���&���|Ϝ���qc�l�@)�6t�7��J4x�6`.ؿ���Լa��=�D*�����x&W�?R�]Fz������)���6�F��%��y��;�3	����t��47*�N[κ�A����c��ކ��0�����M�f�LS��!���>)��Ė�I�{��ve�7���bu�=Nq'��S�x6��g7]T����Et|�D��Fʝė��f@��R#�U#7�N����� �o�]�c�[�F.�ޑj�g�$� ﶮ�W�|J��k��$G%:�/G���h�Nu�QQY3^;�R�U�w1���e���c�$g��:�.-}.3��@��1�χ�Jr�D�xh����r��oC�k[L�.�H��r��5��bw�F����&�5b�"�M��/�^�bj��pr����܄ ����x�?�!��r]MxCC�}�BG��ۚW5KG��!"�;�'���텚�"�^s0��+�lku�&�9S��)�0�>���~vh�|EA6���h4;^-LZd���+��k�)�Wj���c�5O��
i�R��n}�X�����Xq6��y�����"̖n?�V�l^�K��?��Bܲ���z����VK?Zh|�qw�r��z�ַV]=G�PSa3�:���n�x`�f��/�12J �[	فL̷5������_8���Y�/�,e���9�Yˢx;]p&cs'�a`�Ke�b ĥHS#�!��w���qءp�������4�"Y�C���eX7(��*���'�@|����w4�sH���P�@Z; ɿh���5{�՜�i[E���?B	;vB��uUF���7�;��@#,^*Fk�cl��*a���Qq����7h�b�6
k����;���~��p&&C�+�e�9u繎��LH�.*km�p�;k��4�2k�qJ�o��2�w�t��1�u�q~2�<���v��c��.Y���\�@�{奍����ʔ�t�P�b���o�>�����1}]��ѕ�֠+�l�y��~d^�������t&1������ƚ�9���c���~,�5��-1P�7!k�-N�|H�[�Q�g�Z�%b����'�)yl�y*���i�0��"\P�����{(��ro$�O�V�����-\�V�'pkJ����s�vI�X��F{�A*��5��h�	h��g@`B|3��$�5Qt��x�|;��_�kL��:��}�g�	��w	�Wĕ��� ��� �Z/����xE��4�t�D��T7�w����!_l�Ftae2������$�5У��gj�/r����m���r��/�!Ze�͗���"��5Ƿ�^꺶����K�-����'5��!��}�My����j��?Xt�m�czݼ��'�����[�[����wR�U�ʔ I~`��� Q:��_�W�g��-�&�ĕ�RH���5{�Hk0�_o�Dmçz��O��n����F8���KSCRr�A�F�B���k��ٚ���l�����B��c�FS�*۾�YxQ����Q�HE\ט�G��>�%��k��C� ���U5� ��u1�*%����`G���olR�A#�|���D�%����2���������?F�+�V9��2����[]��b��q��lssϵ7q��hL����_�{�E8ΆRy�����l�Ip��)��A�*@�sb4`���/��*����iEBʲK�?�m��!�}��θ7�yq��ﶒ+�{�1�.����,�ɯ���G��Tؠ�9�{�`~���˰����~p�軂;�r�'�bYLz�����y�ݵ���l4@�!��s���~�<�_���Z�Ya+DE�s������2t/�g�T�g!��?��LO��{뾏ef~���:��~/�k�@\C�H��E-�c����>��Qޙ�㶧� ݳl���D����렺rrh&I�p}|���d�y�E�)Ժ�oVx>�ȎJ�w���b�U�3�݇���A��\Bo�vh�ф��$E�m�X87��>B��`w4��3>��l܉���ts��B�Gv�W���j$�#o]��`Xt�i e�Lh����?�� R���)A1b~�ċ<(:?QؐK�p�a�~b&�a��^�o����o�;}��_���Yyo"�8n��MH��a��:s�.\�H6�V�c!gTǘ��<]ۿ�����N��<��m��Ϡ��%�=�,�B�XQ�JK ��;5ɍ�[�)��XY4�܋��*����>���b	�+|0���]�q8^Ɛ�V����O8���YU�����^�wk��}�����.�����<��e�S���*�UX���
4I�����x!���>�e�����X�_��Y!5�p�P&���m-O�:(�>Ы����;�mY©��v~}��f15[��O'c,"�9��
��9v��i#�o�TP��΄������;�2��
{G3ck`�h��|��y�Qx_�@�*�4�����+'O����2��U3�x}�~UD�ֱ/J�6l���#q��4����G��n��ؕg��:�k�A��+�z9×P&y|45����-'#:!�*�I}����X8��i;� ��y��ÖBh{lNܝB-��%	#��a=N� ��r���������P�AҰ�\���� �k����j{�i���m�θHK�u���<;��μ^K�M��[���࣑�u���E�{`.KY���ɔ�S>5�����C�F���J���z�q�,8����S�=��1�3�_�:��\�6ʱ.f���T�o��-�-x��*��[C��.S���p�&�?��	۽�d�D����w����u��Ո�@	�� ���b�:�R�վ�X��4P@9Ȟ��P*�۞���4�u䟱�R�I%J�NY��o}��9�;�,�y��������=C������/��~�n9o��L��۲�J%Tl�Pu��J���%s����j�0c��l��I�H۵�:
(7��ͅ%�P�7�M닐��u��k�����	��DG���MJ������vi��(ؤG��.;��̮���JϞdv�Pb{\{K," ��E�%�٧��+�e�ʾ�A�����=���r���x���۵�8raQ��m�,F������N�˳�X$�&�4��dC%!g汷+��S�U��K���
�jH�r)�%-��A�2�����Ig"���zc���4L�{y�%r��e!�$Ml�1�\'�߾��	�7Y� [�_3DM�#�p�!#��b��o[�+��}mc��N�3���������s�D�����^W���!�k9��n(M���ezZj�ӡN�M`�*�I.�gau�Y�H�Q{
o�x�w'�Z7���v�iN�0�ni�	��?7���s���_3�B�x��!�D�'��Q�i���P�:��x��(y/uh=��QO,~�_�JkYу�I ~ W���
OϒI1�T���?zn�r��h$�Tq�Q�-�����D"@�8�s�+�,�t�݈��Q���*[�u�JQ��T����ህ��l��R��ڻ�p�1l��N���&�|�%χv���c�W�{c��7�=~·��v`�6����3�J����8�@�\�^^`Z\S��$��Q�	Km���O��nG�tE��l"z�I�I�o��?�����Bu�∠Sx0pr~��KS��w¼5�3�>BTo�&}P��WE��~��Or_!���s&���~�fF�c�K��Y��i�ְl�����q�N�x���{<�;�M��$�s�ضu$j�3jρ��3u�-� Fr��D~{�h��81�~��D���~�fb�]�I�NJ�3�UQ�m�����P)U:��[���4� ����ϖ!4׏,.���"۳?�b�P�!+Gt�M�i���~ɩM����wpO�w���� 
^���P2I��@�ް*�؇��]�mK��=�>LQu�o���,��I�أ��?�:D�m?}c�I
��Hy�>_��V@D�9���� �2����\l�4�����K�^�P��p�d����0���xA�����,��"��%��J�������D�I��=�Ժ�g����$h��!vT\
�GX9��s��'���z��2}��7놯�LВ��n�~�W�n��T>�GY���r�/�X��ͯrB���%�uӳ�fX��k$/t����L�S��-�V$�Uy=����A2iᅴ�G�\u\"�&�c�A���/�O�ۉL�% �_������ l� /��OM!�2r~e�;(��
�J!�Aw��0�9�ь�y0f��/�5;X@�x��)�*F�/cc�.���u2�v��-�QX����+S�D�R.x\�c0�� �Ȼ��̇n�0r�+������a�d9?�IB�;��mͩ�C0I_���9�l�fd�G�АČS��=8�ƍ����j����V����m�2(���+H!������j�p���,y�0�+�s�:�ͺ��@_W;��$��n����	�G�8�m5~���NV����Vz2�;�~틃k�%d̑>���<H�x�Є��\R�3�Sh�2�/%R���5��J߳jj����GSq�u�o�,���:O��5R�x��$s��$xQ�) ��E�C{z����!�=�Ԛt4i�G-�aO������l��r�A:��VS3��0�9�BmV��K��D,e�;iP�+Xp<X�N�b��L�L�d7�&$�p��H�y{d��!��0�'\�7.5ҷ �*��:����D�/�Ľ����'"yi��x�g$=$���{�0��rL:�x;�d�����%�?-	P�m9��p���y-�Guo��:��5��iaN�$.���#�i�]e�}k�ZJ�z�"@��g��^��9#3j#%���ii^+NhS�Gf����]�ȧ2�C#�ĉ^����}(��Q�̩`Ⱦ�P��U5��f&3�� ��;/�ֵ&ʤU~ҵ��*2XݥpB�Cz)��F8�=��_�'A�Ψ2��z� �K���c��3���-�V�a�W~�NHwFƒL��j0=\H{:�|��;h��="�����B6���j~݊��p.�w�9S�������%����O�e�
_�0����u�J4��߀��,U�+r��*�Tv�3�F�۶��4�=O�X�fu�fpN�f�G[B<��ww���*�f]Rng[d+W��!~ɲko��4��)���x�X���ۓ���7��9&˫��%PI�̱Aǰ�90�T�埮��M�!�������s�F,��A�HK�\1���@'���%
��pSZf��7o���-��L_�}��Vhe�r��`di�h"v���:lg�f�J��ň��|'��t{���v���E��	�i�׬��)����Af`%Z�3T��9r�Gp84r�T��� �wĖG�I�Z:��M�'���#j��)4�b9)L�����<�a;�OP��߂�CfG��N�7����%J+�͋��[)P�=�Yp ��B*�4�Z�^1���u�4�j�@t�4����/���[K��&�04�
��=K�8�׏%�ʛ�`.�f9��vv{ɞ��b�|�Xzڼ	�^`�d[��0[/�s��Z���M}���Ul��@6���a�ݚ�y���|ؓ,�Ӎp�
�*�	s��.�8� sh�^��l�v�����R.�yɪ
/bƶ<l}�t��n�u�7��B�=A��>���g���T0�)Y�o�����s,�n�=V��E��E������&�9���9\I��=�n��E�*�$�D�Sfh�S#
��*۵(`{�E$Bs_<c������T B�2�b��
bh�>Y����jt�/�8i[�w:!FY%�h�����Bx?(V��a����y�i6�,O�&���4;X�<�j���Ԇ����#���^���jS'�KFU,d�|A�OD�=��$.nv��DG�SM��y��mD�̕��/ #��L�#����oL�%x��U�7)XN�����<\��:�?��c�H#���(�n�v�Oq� ���c��D�.Ys�����״;��,���!�iY"J��_R�0=�7˸���W7F�cj�g����P���������s��"�_@�{Gjg(�J�}U���Jl����A1����}z�p��~����ɓ�-����TI٣����?Ե� �W�
�F@̬B�h�������o
�D�i��g�"�+01%�|���8d�b��(�&��w��e�ʴ�'��mw�-#�Q@��օ`0�\��;��JN�muu�0���ȒуrE
��-�'�v1*�1U-p��H)�P�>R� ����B��a�i�/��P�)W������1���^��>w�{?��%�F�5�\�Nw��5�H��7u�������y�&]צ���w����9��8!I_^�D�c#��F+.��F���Z�f;#��i9}ׅq�f����)���֏��6]���eVC�h���mӰC*����6�^�&�����b\��K�l��o�w�pb�Eˠ��e��,w�'�Se�(OZ=��Cuih�W�������Ex��lnׯ�v���5�k��Q�n�͎+�(��4k$�7��f�Ֆ��X A�L ��/��zV;R7_#�ܕ�[��=?G�^�<[ʱ%L����=8��|3��Pt��>����{��7t�({�lݼS��|7i/!�^��_	�g&!6V�i]���h������qo�����=|�Z��LY`���(��!�s8s�kKIO'���;�Zbl0���GaOB��Wj)=����R�f�)"ͧwP��Ґ����y` 1lM�;�p�w?B�\�SORL��A1��<u׬��)��Xќ�7����K!�D����)Z�l�����Ү��g�x����#"!���Ŕ�d�x��cǚ�N��5�eP�0J��P�Ú;U�Ik^rbq��3�%y(�EP�y��
�L�Ppz� m^�d:�o�,W�!"�(������l��~SsQ��O[�ѱxY��i�|��Y�_������'��^A7`I|�����g�(bN�,�V{�W!��HM�;��R2���
 �z3�(w��Uh�T��y�QP���jpJ��5 �l��M��47J�saa�$Z��/W��?}=��'�����u��F��9���<<�*��h���̼,0�{����?6��Z^�A�������	t�{��;���_l�i���a��M	Vn��	��$���KH��|����~�;W�b��(��M����8����W�<�m�[pDL�{�(�J�)�Ko��Ǎ�, 4�!�˂Fl���/�Y8I*d�5x���a�ĳ�]m
�LS�4�k^k�7�V��)Ö&^z�<��>�e��M!�
(�G�ﶫ�b#����y&�u�,���8��82��?�Sr@�e�q�v���D���ߗ��8�r�*�f��jN\X�g%�9Ѫ�@�,i��=��Y(��R��'=��dbz��ҽ#	���xP<~�N_b���(�W������@(��KBpU$�Gb���ԍ����@�����gXc0���ŀ��5�N�m�è�5t��-����w��$[�I�:ۜjXʜo����k���_Uiܴ[.c�5\� R_I�-*��mk�u3:�u Ϩ��+7��M)����J���� �?���G�,�`�\�D�]���zC��a���P/1tz̟��[b��L�ZƐz�bC�JmxF�o�
UH�2]�p�9w�?�=z���1|ȼ�M�M�ULؾ��&���h�d+2�b���I�$��e�ʱ�ZaR���&��~e���IR�S~ɣ�P�Z��II �3�o.��M{ؖ��i�QZ4�O͜�"��F���/U��Hu'�W�BC��� K�p���r[�R�C�pJ�߲�D�trm��6��8�����J����4�e�\{��)��M����4�<̵�����$����M��$1GS�����@s��%e]�"��??YU~B/"��o����Y<��T*�j�w��]�=�jt]I#ݚw��b��� �1e��#��1�_$��^o�f�=R��o g�-yl���Ɂa1�<[J��e�a�l�8�s06��x������ߋ���w�o��u��L�Њ�Zs�gڶ+�ԔP�۷C(!��f?j�����1W��*����!<Q	�������\܃�&~���_�2�p�W0�U�L*#Iu�.��d�N���ȣ-dMޣ_U�����-%� ȧ$
q0��2Մ������s�u"
��X��r�ل��R%��[,1���ڥ���9�醪��i	�]���y�������/��D_��ކ�.���0����Cu�?k�M�@~�q���v�+l�F�ݎv1�!oq�	���Q�P��Au[�"��)��RI��DeI�����]�|�]yz�ͪ�<	�U6 H�5I|�k$#�^�]�ӨF֒`/u������͓�+��m��%�f���UW�h�d}{'i�nN��_ۼp`�L&�L�\�z5����+��?a_ ��W�ߦ��^8�7����w+1l(����}2��'�y6���DB9�B�J��b�ZV���3���Ŵٍ�>Tr��o>Lأܣ�+bt?|J�َl�F�q~v�F��0���l�2�b�H��԰X鳮���YK�*W'a���%rp6x�2�J�U���YyF���S���#�&�0�|<��f�ˢ��5qLWԕ�gAhJ�$�v������D���qr a���iBZ@:�{p�:����$i��P�1��d=aZ�V
 $����B��}�P��B����P�dh����F��л���W�R������,%�i� 2|2�>߬�:f�l�0F=����5�[;5�|�nH�6����ּ&�%Q�X�T�����
�h���C0$�\HlYQ�{�N�@r�������w����}�U{.��*��*�;�(�{�~���0l�����cAHk�-j�T�>ОR�q�-�;�
]�lĉ@���U$�n�Lp�����諺���}o����n�%�IYeӒ>����q������W���uF*����}%�3j�/����Kb�b�f<㧡��U��	wŨj�B����]?r��y��ÃA>۽��AhE=%#�8��1�td[BI?�dX fr}jP�r���S�P�ҽ�����rh�4����a��g3�qI+H�loqK��C�d��+�m�U��0t�
[!6�R����Y��OK��%�I!���F��,�+$���K����Т.r�4n�h�+���ג���������W������aD�ni�����k�ا.K�1�뾄�x��b|9� I��}��29�/��A*���֝c�17 ����
68�]C~4��[v�s�Wc����Y����;�_���D;�F��4��2�
�o�>��{����Lq�$�)�rS�%*!O=A],������n}0)=�����3㎾j�='�>����2W�=���R�}i�2��7�G��Þ��~Z��>�˛���m��X��q���35�(�a�^���>��DmH���� �An�����:˴E-�i�V(Q�0WP��,Q��cT����^d`ߑ���p(�6���2%�q�@��1۾vB�n�ȱ�pu�s=� �5kX��%�-�j,ޑ�(q�2]e���R����D��᩿+�!�:�
�l��|}EѮ!Otϻ�@�	≽8CE�m��!RR6���"����۳u��;݁ԛ�w�� �wD.�� x]�H�����F�w�u��I9|{�TU��}s)�����"��z��?��MP��5',�A�g�ۣ��s��v��Ȏn�2j@f��I=$xva)t_z���iq������8�rm���r���Δ<�i���W'�l�}�n��Π"Y�x5�=����}|w^ݩ�OZ�܊d��iI��rJ�RUS�M~5}$�1
;�1���ڳ���'H�Hfm-�W�(J�N��#r�ѡH��6ٹ�2Ⱦ����M�ҙ���!dإlzx��O�^��3�m��*:R��ur����M�	�}Up̓��X�)�^٧�r�.}����)n�>�W�V�>�C�W�q)�����Z��ۂ�KAҋ�F!��n�K��&��#����1i�mvm	�V�݈���i���jT�� Ͼ_1;&��.3{��
b��Q�8}��2�:��	jߏݼ�'eI���+�����{T.Ё���i���p擼6.�k�'��Y�I���'�$i��2tz��Ѵ�*jX��w�,�oĳ�YK��L���v��qj��O���^�Bv�qc8������_�"�*f�d��,#�t;���`FjB���+�u�$ϓ`r�v��F����Y,ku���r�B'�0��y����Q�Z�5�*��t�n5�|R��r��E�Et�-0��x�4��!���n*i��k�͛�C�6�[���?X�s��B�1rZWn>k�o���%������ �Y�p<�P����w�(=v��#����RW[���G��y�=��&�)u�޵�sH�Jȑأ�փ	�PfĎ�ں�G�5�MP�U֔�����D�VCG��J�Z>X�ܰ��%C/�a<�����h���p0�j�X��E~w�B8��Y�C��a��g/+�3\��(����vFf*��0BS�E`�5�RBW�Z2C��Q�����aΑ�RZ�+���J�u�0,�Y���d ぞ�z~��d���;Ǣʊz�����.o��F7���A�S%�dKkƯ�~��h�L^{M ��8��>�ү�g��Y��M	�j�ࠔD"�������N�TRLp�w}�R|@�e,;E���[�h�߰!�B	�5F%�|��,�B[DPN��v?�X mM�Q���U�O�Z��.�WOJ�T��k��ϛ\�CE��r���FX�/�2�u�ExY*�8����p���=ؾ_jP����{�	$�+����'��EѢ���������̪˛�x�k��&5�������i��|�?�̧(!>�f���H�����nD���"�gsx���I�S��J��ɧ�Д�N��:w�	;�֭>���B�O�袮cƈ�>��c����7�X�܆DhfPӓ�[Yg"��e+����q����A�wr/g(���m0Bs�Zk��$)}��y�L<bE���@'k�Ӯ�.L���9�/S���]ak,g�Цț�?�^w�Ӻ�Ǟܳ#�я���C�#(A__e3q� ��M���Qop"��zl�E�G��T�Rd�ⴀS�ᾔ,��J��Ż��_rM_��ޮ��PP�]�+[h�fNn�T5cY̝����5�B�u9ވ�%$2_�v�0&��wJ�3b){�hgs�@����=��E�w��f�eq�M�lۈD�h��)/� G=��)Na]�`��i���y��iT|��0ק��d<�SSG���V�6�AQF]�0�?;r�����#���y��GJ4j����3�%	E�ov��Dܴ%�)&K ���>�!XsH��xh���$j��-���s��q��<A�e�Z'��q�3����26Q�O�����3p�Xxo�F+�I���L�]usO����1���&&��Z(\���닃ȍ<r��20Mu۠g��M�ME�Sİ
�d�z��0!�i)��t��O��z��t�$G�Ys�Ӑ�I($Z�bfk�1��LP�0�^�+���(	V�R���>F��B��?V@���- �@,�'�  �Ҟ��JE�wF���r|�v�PH�c��*x�x0�|��R]�ϡ�&�B��$}�ԫ(��cO7Z==T01aQk��u%���j�8���61?���<�j�W�W%Ԇ������|����g�6)�Xc����NP?\�n���v*s;���	S��(�N��b��w���r�FQ�6��?5���3�X�,H�Q)eǎ.�e���Ay#�7��'���vg���Mt�u�j�S�kj��j�L��O!�<���h�2�BU	���� M'4�?�%>���������] T��[��e6Z�0��l�c��W �P̾�Ž�f���$��zHB(7L�OVv�&��)�b����=�S:�L5�G��g�����$\2H�\���2N��v ��Ǭ�-N���
�D��r����bw�������SGL�-ht�_.QTx��3�h�=5�T$�L�.7�F��tsx�!��<+��+)��j��F��BB��K��{}�v��5bǙꋴL�"���2��J:6>U�_�)a���.�z��a }�T!vb@���8"�fɺ��0�dY��9*>Ȁ�2$C-ϙLA�p>|���}X�_8�g�T3�?�H�.�����j�,�UXQJs���m�*eQP�S��N2P�o0i�`M�^pF���빇�~2�)��=HV�F_�˿B_X�Zk����iC�t���Z��d�-ͳ(���BZM3��	�)��ӧ�j.�i��@>���rj��1{/�FA�%U�[F���2=��+ jx5+Ɯ�iVF�9p?�孬�߾��':����H� ��Ղ1Kt��@�]|�@l`��S��\�[�ySUt���Չ⫄�b5��1*�7~��~��E�B�pr�즖�0�o��!�W��2Ca���]�Q�R~��NQ4��&᭚8l��׷�L�4�C�&j����+��ո��cx,�J�S�K��%�m������rU[[p����V�X^:�n�D}�O8��l�rxRR�l�6Y���;�hX�#]��U
�x�b}��iґ�*���ӑ
H7�u+#��E�ӈ���rYw]`hVZLW�z֑m�>3���I�{.����o��\j<:m�+�S�k�$	�+�(2�89��������J�����k�{C$���"���	�%3���-*�h��K� �9�Gg���ٶ���S$̜�A-��;d-r�6��7P`2hq8����	��m��f��χ�\�C�-p�t�����t�G���5�ԅ�B�`�QX������U�>2f������KcՠϦݎ|9�~�v�,��&8���*���JC_�p�Ud�x�Y�t�(�4���7��������3B^��-{Z|z����υ8�z���(h�Ԃ��Nݔ�	�H�֤��iw�[�LiH�Z,hCaӵ��_t���w�_��O:݉N� �)]�W_Pǉ�CY�i�cgi�,s�#8KTo8:6�)�(�d��>�?kI�9��9й�h�}-6� b�a ��9�&u���4�fpZǮ����"j*��Jl�`��y��f�R��]�/0B�g�� Ώ0�at�=�N8X����oU��Vh,�J�[���^������D�F>��{�����n�T-z��n��XI`������|7tW(/��4�)�cdv���;�RT �g-?��Ѓ��q����K.P�{^��n����9wuN��8����0�(��C�"�8-p9::�~l^����ޥ��`�TM&g��~�=(��J�+X�n�]��r��������$�֓��f�j�1*�똨���ib�z='q@"03p��_�m��D�Z�=@��5�6��K�%���J�5���(��m��1���e��F�?�Q �c��dVU"�~ߤgEI���$B��}�|-�9r�	(�s��&�.�?���dBhHu%|H�^ۦ��w �� ��h�g�rq3v���%�D7X��-��G�;fF��p@7�CY��"�N��8�CW�9��W�R�xR0�D�»Jri���	2Gځ���?"K����CbmR�_��o�����K���g�WW�P��d*�Q��̟�}��*����= ���X�<'Bs|)����AC��6�-�͉{	ise�,j���nÅ��0�?�p�5��a��J<�w��[C+�� �@���<�uuĎ�L�s�e�W�b�Wd�\�=IW;F��_�BC+E(R�,�3E�^Acf�?}#P��{�2E1-�7{cZW�KH��j�Z9ǬoG� ���/����HZRC��CT�I����o:����z=y��A�˥@t��������$AEl��qb#޻��R�]�ܳ�m�'IX&m�1�xf�]GTPɢ����B��N���D�~��	|���Z�'�k�ˢ�:��	1mR�	���` f�V���ū�������� J�e���L�'R����)P�f��=�*S�=�6fi>��Q��/q¤]t����Ěږ+���7�f/�s6��(7��:2��X��<}m"W*�%��\Q�W�N��$=I*Y�[6Y�<��V�:Sj��^�\��f��E(���5d}!������h�'T[��7d÷����I\ !!�s�$K�vS�X�٫{���t���5�;k�o#f�qp�N؅���IK,���G�����=d��Np|F}n�8��+�K'Q�DgL��%a�o���p=�s:){fb�Y�f�����f�.S��{_8�Y����@�����v����VY�#�Ws�9�'x���k��X���&t��kD�j=+M�v4�
�=R�ٳ����#d����r��Y��ayZ)�A�I16 �<��͑F~��t��1�10���*�C�M�޼�Hg�'ӆ����e�Z��0ޟ��H��d�j���Z� ͱ��$����4w<.���
}!{�ɴ�����<<��f�=�4, E��yr��#w�ng�L@2��{]Q��
��G�|n4��չ��O�bvO��1Ea%#8'��^ts�ȝ����Jނ�S;/�����SE�-��$b����#e�!��!ҶL�Ei�y�I]�ϗ����f�����a�D�~/�o��v�sw�,L���=_	iӦr��ප��R�:&���Ϧ�Ȱ�l0(���j��1��j��o�v�b�PF�v-QƳ&)��L���X�b?�[w��.C�=f������5wF׹��u���H�n��^��e>WueJ�v�VǗ����2��8��LJkG�f�A�e�B �@�\3h�����?���p6u��#�M�8K�3|���$��{<+O�o��Q�����f?�_kFv�6�O�����G�h�v�+ٷ�>�!��B�y����K*��G
��&3Hi����i=�OhIH>���9��ɲ���*����.^կ#��z�L�Pf
CM�tP;�Aus�<yz��� ��O�����C�WK�(��` �_&}a�ԁ�dAKIý�{H� ����O��ܑ���w��˄���$��$�rM�]� ?_�j�3�b����o������>)#R���A�1m�ί���������5VR͸�#O��
1�/
:�F��.TE��>aMS%��ۻ;��c�����Ó�/��r �|[#K+2��ib ��0��z� ���^O|lbJ��J��39f�r| �x������rvAboO�P��DW>B�r^�ǱƸ�Ny�0~�޻�6`Q�{��a΀\�_���2��h:��_�a�鏒˴`U���ֈ�h+V7�=� 7�,Q���[i�"�2��w+��Fy���f����\��o&�b�U�+�
V`��5�:��y��R��s�*��4�O���DNW`�hF��H8�C!�MU9�"�C'�ou��w�)��R�Ն&�� 1.��#2��N�$���� ���u!���5P=�>w���WR�=S(���z�RX��(��T��Q���!/`���c������Ѹ���Q��)�E8���D!Ί��&}����q?��	��'O�0՗�Hl�J�t�p��_ewؐ�<��KLJ�TM$���e1����k���XN� u\��=#���vls b̷��ks��k4��2؛�f�:�џ�#`�E�RlXǴ���o��М\e-2�RE 4G���I���*�*��6�W�Sl0Uω~/鋻�+�S�"�Ӣ���D�i��c˄�FNęWPT�����Zo���(����s�E���z喀�M�v>P6����R6VgI^�Qq*�a X�됺�^���*�,�P�_��*�����o �\SJt0{����bܤń�䍱+�w>�S������tB;�P�~����6V�f�%Mtp`l��v�'��=Ch�:j7O��Z>[��U4CO5y�ԛ:D�BRf��ف#8���Q/sW��Ǖe�jRt�J�.�����$/��4�@k=�{k:� h/T��U�������Zݼ%�u�� 0�>�(}C�V=Jtd�}� ��(��͎��~so~��`4q�Tev�%):P�*{2��_A=T	r��؟�*	�2���ıl;[J�0q��V����D	8ϓ{��\�VIe�(;�۰�
C!
�g ��0�2V�9b�ы�5C��B���e@�YkP'��̢Ao����%�Y?���#�����u襭�c�^C���[�S����hQ��<�n�
�k��T08f⒱�"L��s��Ɩ���C<+��3�S�2�_P �����A���d�ςm����\e5��rq�,E'V�f�)� N��%�2!{�,�[�B�<�gܝ�i�aMZ���J��0j������B-�0��V����ek������XW#D@������tj�R4������I��~BfHw�Zʃ` ���nb��\3͒�
hQ0c>�ɳ{�����T��g����b�
����E!Y"2���������#TB��l�E��Su��K/�,��=�\g��Bt��I�0uu���D�kV(������b��^,�� T�z�X�һ.�/K�Ni7�(����{�{l�S�~�����q}�"���ZIG����/�9݅B�	 '2ٚ�3FpG�99���=��	ˮ�b�,�U���d��O)�r�)���Bw��P3XOG�A�K���LYO-X!�IA�Usڀ�T: �hh��蕜�eO�&�?i ��a������d�g_�>4�]�h�۞�u�v��I�=�`�̙]ٻ����jA�����&�d�y.�9�U�Խ�Y�|��Mw�wJ��)�<�`��L�-�W�s��f+�	J�����������'(�}��~Mh��0W9i4]���Ϸ�ۖ���ᶵm$��c�`�Z�.+䠫�O��66(<m���_8����^-�}w�b��S�����!Fo�d82����s��*���m�7n��M٭�����0����]H娀�ĩ�͏`r�H��Ȭ.#���AA�E�pAU�.��l�sk:�A��v��	�6���.;�l%�鱰���%D�wE��os�F��R$JF��a�}w~��ن�N�3.��" �j�o����g����T�0��^�*�Ǖ�H���M�B�E�j�}�z�Y�1��&߁���a�L[η�P�,��N-( .yѴi#d8.�k_�O�^+ƨ��ثfD@�E�
X�[衲�Ku��gp$��7΃9r�!�7y���}h7=Ό�
�D �������;IոI�A��N[X:c3 �p5���%H���1p�k�`�tmې�7zF���T �Ď���}�߅�!��e���&Bd���&}�Q:�(�b�y�$N�Ha�X6~���F�V�s0"��U�.Z?��'=��������2rf�o+�X)R�k����s|w��<����P��=��0}#cX~���W�1�պ~n�]o'�=�Y0��v��$�B�!����0O���?���0��x����5ڼFA�%��rm��2?���=�����g��!wmB�x1�K���`y��ո�Ï�@���_�`�*�_Lu��-,���CA�Rz����x&�B�04�X�D���é������A�I1�I��-:w���Z�����'� zߧ���Z����y��!�? О┖,15 ��8 �62��0�"���@w��T�<&H��J�������soF�c5sr��Q:��(%����[$���'�T{����,�, ԃ<]�*4��B3�r����9SD��_��Ř��P�8{��������H����fl��+� ��m� s-���)N�,��KR�1�hb��c՚�h�g��r�_�Y:��7�k͗rc��h�ԅG]tx$�T7��I5����7�_�Ka�z�l��iwl�	�O�g�Q8_�d|J�[��j�*K�=�ήX	���o�¹�!hv�� 9����U=�54זy`�|bK����H,���FK��F��oE�h,� ��}O�D2��� H�z�#��g�a��L	�K�1�x�����p~Z��#O�P{lHα����"��;2p$��.&�}�i��~�^Z���M������0�Rq�)��+�Ӂ���Խ?A���"Y����g�+&3�&��)�;�E,t����7���<��ܳ����E9��*�Lc�sq��KR������� Ig6ť�c����^6��x �G1(Ɇ���#E����d�Hs(
�J�ma��^?B�^߅������-�U`o>�e�����Hb�H��7�"r{�w]� q��{Z.�v��'*{)'�8���S�%Nֈت~�8&�7�`��P��RN
i��4fe�x���#r�'��5E"��_`������E��?y�7���`F�8=�$1P>�4o�fq��ekU��=?b��|�1�B����jQ�����F�Q����#a�5�2ʽ�TF<�)�H,0k�fLτ1c�é��؁N�sE��t��`ʪI"t?���1ݢ�e��X/Ek|�w�H�$���^h�'��MJ�������9� �
A<�W���D�����a�S��&POn���\��
X�uv������V�9%*�x,J��/���{��7pST$~ҩ:��y�ۀ����;%�T43ڌU�aL��P����U����U�!��8S�lU�Jk��4�60B�F0Z�=�s��!���4�} 1�~
��)&hOA'9�i�◠�d����� ��0@�Č�� �@�=�k���w(����Z|����P�Fx[���nj�O:�\�܏�Z٥�o�<��V���S�hz�=�1�ja�>&n:��LY]�4�i�%�P^�X����&C�oF������f��xR$��;��, �g���OF^�Mm�i#�Gw�:��y�^�Wh�bJ�}G�k�^o���gZ�C�-�w����U����BZ�)��D��E��Ī�P�"����fH��Ih����!k����܃X�cC-}�;S���T P��/�J{֓a��d�a�sܽ�:'D;�f������&*�>Oi�و��1�@s����6�P�/��7_)j	#�r�~�����A�&ৢ)v)�K}�o��R���ɠ:̈́f@ͥ�>��e<�w�C@���Rj�7�ma���	C�0��ǝ�F:I��C)?*\Qbϔ� /��,��4�'���l��>��&��P㾂Ck[��y�pGk���#�:a��f�����dы�܏��S�"��Ύ渨�f
@�֓��}�]������-�僇G~��qc��xߺB|�S⏆֤�����QB�%x�	*��׏�� BG���npϥ���V��p�&k$����du(��KcpX|r�����z�k�!�d�Mr�J|��yc��������� �Q(6���mB=탇����Nua�k&���˰�_�P5���=sҾи8���(�&v�w�<ED
�`�Z"�܏D���|�T�����/�W��;D����Eu�QAB�S`�	���MK�/�?�̈́̍����4U��I䞓�	���{Xoz�UM&���|�b2�H�A^f�ł�z(�V\&!PxN?��ߍ�c�
�p�;)p��Fc��i���:C1x�ӑ&�w��� �/�`a��o�x�|/�j�;UNW��[ˈ�uPT�4P��l&?��@h*�:�B����r�7P�N-�W=aGF��,��|�e,���z�沣$��w��f*�¦b"Ԏ3�;� �r��w��M������͂)(�,���V�F�W�k<E�?g0a:X����/���
�w�y�/y�1}0�v�_vH��{AE/��
�}e1�T��1�Fn�=�0���o��A�r&�����q����M;N]9'������EZA�-�����w�/��X�Pe�؝�}���U�H�O]���� �Z	�z��
��%��u6u �̛ٞ��JrX�{� z{��*���JTaS���_��K�}�n��Z�?�k����_n"�m,��@��c⴮�ڥ	�ym �$�����F8���QԴk
���I�W)p��>��T��˂hM�z�ڙ�S)�CO�vq���^�}~e�GcS�$�v2�n_�`���J�$�FYeܗ�3��굳Hե6'�=��{�e��DFg����	���R�P���`��r�&������~@=��@��O硏K���/�����+5����Iͪ.oP1!l��r(n���Ł���C

)�$^:��Hk_sř�ۺp�������%
�@ͳ$/�}��X���3ż�������s��u�+3�Զ�e;�3M
6zr���WpO�l%G+���ra��,�O�����s0I4�
�zS��I��P�����>]4X��ͱ�m�Ɗ:�ho禛�j�J����d[��M4�����A��(].�,ђ?���O��y����+�^x�XE�1�A�)�x�
@Ei��	�H�TY�%�W�g�X���T`4��V��m��-������k�y�ǵ//<9g���nOS���l:����u��[�J���T��k��n`�Za8��e�) g�欰	������{X��XQq�F���E�%I:�R#�́u"��Pq�+/پ��������a������n��	턥Q�G�3���\��6��8��#9g[���A���=�$�����T#�a���|�[�$õoH��e�b�Ј2bwG�@�H��([��U|n�ݞl%�q�H<��M�CX�ᒷ�\�ol�G�o8��|h2�_o�v���Y
�<�B?j�B����<9�^!ٻF��5R�a �*���ڏ���t�^�Y�w��C1��������ׅ�?�� �^k	�k�%;Z��|��T������N�p�қ��[��yCW�ʴj>牞5��F���5:�YA+V���w;�
i���~�B�^�ݳ&_K�ƅ�e~�W@Zv�[`��5��m{��Ī�1�v�z��UO���e�7h���	4���h��#ﰆ>�t��Kp�<�Z��s�@,%��;V=��Q%F]Rb�	#�?V<BP�A`�RaG#��oKݛ���=a��Y�N�	g@�����	��Q�CC묅��ƹ�	[�΅[�g� �WD
�����4�W�JR|?�*���x��ԝ:9Ġ	�AM�p#�;��?�K�}z(�DmEVRYI� ���N/���{�2+�aGŋ����@kp�r�����-|�N���)���.����mE{�0��z��7�kr�!Ƹ�ueb@c��Z�`�+����g�W n��w�Y�� w�W�$v=�#g^u�)��x�'κS��hg�W�2V@����{��P��T�fh����'���K#�Iƍ��v��C}nz庉"���V����Q��t��� V���k�@tD���_�h��+����u"�1���G����e�݉�ы6�������e�̂p�����4��3��Bn����|5�1ix���نI�g��*R�ۆ�5q�j� <�=rO&�^:bH��QWߍ�<�f���\Q�CBr�!,T�"Ԛ>$h��*] ��B�����ƶ"�W��$ڋ�}8��
C[�.5��z��&��x�"}_2[���|�4�Yǋ*�.�gH�מ��$t�װ��,��b���b�Z�,�߆�)�#^�A�Vs�@���c������8�����d�+�^�^V_�/�>��W#�aU7a`d{k�O*�-/v�&\gdj�(��%���${1�ָ_���#egU�p��ߥ�#���(�{��0v>2��|32ϔ��T�t[x,�	�,���/���;_��3�[�;���#I�F�d�1�Պ���}����Pm�b�^ 	��d�?₏����,��"J�*u��
�5��
$�Z���e�b��D����67X�Q��*+kp����g6��zw���x�.<"�a�n	���fڍK�a�O`&�11�3� �>�����ף��q}�iC��F�ҼϞ�����Q�o	�4��e�� ��-�x;�Z�%(��QH����鷉GR�X�{�#J2W+��=��3#��|����&��O�x����>���<EBv��p=ţ��w.ۉV״��c7V�Pԡ��;!�����]fT��K.�0�n�$�T�
A5�6��L������nDY��y����p̉�TVl��<م�ms�)A�-��jC[z�;�ɛ���Z��d�%�����.kz��P����S�>����f2���g�mm`�q�E���~���G�CD�X���7�esD>��cKM�h��̂Џkn𢱩o۵�72�K�cm���?�߯�w�q<g�y)�f�p4�^v0����`�D�#۰��6oS�ʔ-j'$Z�y�F`�!h������� ��2̨8t���Qܤ��mv�B��!� �a(158�{_�� B�6��/���3J�R!Pk�!��7�
ݗ�c�X�-}>mM�kG��%W���|^!�rL��P$pd�������?�����=���/+��\׃�"�%����EVnz��w���%Fhs$��[E�g4��@������IEl��)��#�~h��"�?0(f/b�s;1y��1F�+�*3�z	JR��!Sf��G�B�1?؂اsu�1����"��w�mv0���/�uTG^=��n��S�������F�9�3�	FR*uM8�?��Yh���|?���o�q+h�2')�b�Lv+;Y���a=hU�q��m��ik���9��]��q |�h2 �	���Y�`��ȓϚ�Ӡ-��|:��	�;�����i[�銐�@��~���|E��㣀�y��"�Y���k��7k.Ic'fߘ�x#�۳�ϙ��ښ�~��tO�Hq��gE�~?Pl��v� t�w���J=O���&Lg��|��x
��~WN~L,:�SB��[���Ց�z�l�P�*����TG� ������z��&�}�O�ĉo.�h��l��Yg���׉���\��2ӈL���~�Z��o��� �����H.W4��ۗg�}b��s�;��x�h�:V�����m5��� Bc�b:��.s��e��E�Hpm�/�T-�z��KME=Y�p��(߭(����,�U�cf��!7U������[��(DZ�J�B%�y�������l�V���~�5Ҕ��b=C;��[6�!�E]��d(E�w��C{�식I�
���u|���D/p��f���fRn���P�v�e��`C�GwS^w���>����,��`�H���p���H������yH#�y��w�l/�_����_;�yq�:��NV;N��Y���f�*T�S��Fљk�/�0��S ����:#�n�
m�NO)H�TD1����a9ߓ#��}"�Bsc�=3� ~�t �T�I#)�C�ǰx&�q�1�k�R����(���#�x=�;:�ֶ7�Pn�
�I���Ԛ{�9����4x��y�hH��H�uJ4�4�H�G�z4�#�^�Ve��UMwy�H��jvr�A�ʍ+6
�J�]�	��l�d��M�]��]-On��)P�|)�$2Ae��.�ޜ��WRkui`)ޚ�����;���b��?�#dC�[�D�z��l���b �����dv�J��|��=��b� ��a�+%�2]�+R�Y�Ex�v�g�_hÙk
BthA��1�������p��e�y!�uu��)pL9������.�XW���:sA�������l��3�0V Τ�r��	T8��9C�Q.5#��{i�sS����(3���s�s�U5�vsi�K�XINY��Ĥ�����EY���#�;nV�ʤu�$4�K�@e��`�׬p�׫�\��S�S��� �KhH�v���}��-�AߜFFCs�G��r���T��e�v#��|��Uk��HB�Y����>�}���� ��H�)�cy؊?�N��=�U��-����g���";ث�dK\����Ym�ө9o^��O��ޅq�0W���:����[�[���謞a���{r�CUF7�ͻ��-I�ߝ)H� k����x�\�\
2m�"�m;�P.*���I�02U�7�wAe���w�&��]����D����ݏ�):�fGGz~���[ߚ��E��W�D���mUx�b; x�O�!e��ۈ�h��z��۬��cG9+�dϨ������e�XU��7�"�!����˷s���6�'cE�����0�'B��P0Ar��-So���Qk��i͖ζK��5��(�:�Mr�w	�g�9tfD#��r � �#���4�BHDܸ)��u#�yv_1�ǋD	���ɀ,�~k^uU��K���7��1ΑBI���W`sf2��
@��ˋz� o#���s���m��gp7_��������3U]$f�;غ��:���BQ���_���Vp���e>���H��>U^�$췩N��9��K[����[3�κ��=u���P&��!��:}=�S�������Fuy��R�j��v;��8���쳗��̜�cϑ�xfu��v�빻 fC�e��Cƴ=�G�Y������3��;�A
>5��g���ݕ$�[�WX:��_�q{��W�7D$E�%�dbIXd���n�wc�"5Ot���[l*��iW��C�A�zj+Kš�nv�#�,��by	S�Kd�ǟ:���@x�g
��;F`3��1�N{0sb!%�/S�n�P�ִZ8���a@�� E�VǦ����"�g56'Bq�e�H,>�qa��ޢ曁h�'�ϸ�����ZK�9��+q�tjg�z���0�����