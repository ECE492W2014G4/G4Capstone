��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P��v�"<ߞ��&'��k%P碶�R�ӣ�sĞ������FY&���P�%�YS��8�T
M��z\���0���@����Q����դr��:�� ���ʥ�}���D�3L�_^ �����Fz]��ȧ-+�`�9�HM3�q����<DO�T��|���Ndd����>�|bW�hs����02q`m��U�s^�-|�M!���$f��U�d�H�u��K��)Bp�r؏L�P��)B�i�@vQ��C�c�i�3^|�
�����/���Lh���g<r|��Ǉ��i�9�������.����W�{���~Ш������J.X��;��d���S�(�M���7�������{'������3T���s^��(D����W���<��Q&I=9:Q5��H��b =P�@�o���B�f��H�>Q+}^C�=m��6���T:���"~-���7�;;x�FuJq�%�k��^\��Y���Ϥ�!F�o��d\�&��e�'��[�}|ŅsA���5.�eY��0����G��㋾�X�dc�/�ydK����N��G.l|�!���.�;��~Ƣ)�-���WR�"�����@�oZ��Wr�C����Aa�Է�����|���LBT�q{%Z�����o���K�8x�ٵ5��t��]��k4�E��6]�h{4^"�HdD.�Z�V����}���g���8=�����t�)\I��8�X���:f���sp�sZ;�đ.I� ��	1�����^ᔑ�=�f2���L�XS�� Ɠack���Dt�(��48w��4̘p�w[H��Dl�����DpB�o��_�<�Ϟ_V[�D8�RU���z�ϺW�͒>�.��N"�:��䏓57�G���U�Q�]D	�/�n(I<�r����3�� ۧ���P.#��R��G<�h�F��� $���J]��
Ji��A��J��?���Ju.���Q#��:R���)��b&�<�Gg��Y���>��щ�E:~j(|�H��Y> ���.CImG����~БN��7���meEy ࢮ�b v���_
˯���e����\�u� �/2��?���L��yU��=f8!ȩ<i7�d_��[�.�M���T)3`Fv����� ��~�\bȉ%�}4��{�9�t?,�ճҊ�b]U��h�k��UO[��&�v#`����α[�\XƲ2Ȓ���e���Ĵ��TE���iז�nb�Օ)�@��T�U��n��M�_��׀fDںFU�|���z��y1�������o0�ֺ5���[����գ�t1�=�ӂPt�<��G�"ï���F���%tz?��I��i��4�p�(
�
6�;�	�)��(�K��2�'� �*��_�ޠȆ���sٹBґלI�e/�Jr�_�j�qv��}��V�i�A���,�4hơ'��6�/@�RW�@m;3�c*׈�]�X��K��ۏ�Ч,�d���=C �*[��t�G1�4*݅��0�3#F]�&*�cD(�pk�d����fn�ǩ�&��/�>ʮ��2D�Y�������Sˌo켂�RG�ܝ����T�`��=��]�d�&�Q}f�nz<�x���"�?�@)w��D��~�Y�A��d�ۙ�^�hƂt��p��a0_v����#�H�ϳ�y�Mh���T�'�>�e�س���Yx&o�}u�3A"&�?8��&s�}/~�e}Q՝���2d�vq]`���xQ�<TO6��(�RJ<$���M��(���,����੐���*����z���:J��f�wn*m[]�Hb�����_�) yՍ�Hh�j��A�t~�F"#cK�Jy���xK�����v1{0��L��/!�bB�Z���<n���EO�%H�7��Ih�3�ې�Yl��#Ь�1���I���ͱ���u�5��ʅ1�gr.�ix^a��ji�:�������jℷ�%S�麻�A*�q%ؐL :U��{�����1��/t������gy�Y9������,Qi.����-����"���J�eB��3
@�z'��w.M/����L�Թ�/ �3�[��^��D[g��������+t�P�D iT�������\0%\�G��H�����C[s>��t [k�
ĭ끫C����TG�k�*O��������
55��M���'�D{EL`�+�J��h�ޑn��W6!����ܞ��Z��uJO-t��镱9D�DН���O�O�����)ΰ10�U��Q�A�ʽZ*��	������Ї�s��N�6Ƒ縲6�s	��H&g52(���1��72��g�=����awv���s�yeم ���k�H�1h+~B�g�hM��P��ȃ����>�U�ɕ�'��nO�<5{-�!2J,�@Y'~5ؓ��X���O
�$?�kg��n�~j�}:|�+bi7��2�i��Y^�f��_5{"q���0@,!:ӣ'��BQ��7!�I46�JWޓhOFX@"�N@ٔC*~������/��";Ej��N����Q}�ۻ��J�!��bN�D�~�U_c>!pn��i���~8�Rk5,��q�h��'��<N�p����?�6Q���sa���a��W����[P�*[���
/�֓�R{} ]���&:{����C�ѷ� ��4�2v�4Meh~������ޤ�]$S�W�JET��C��R5L;���R�yC%؂~�4_�Br��?�%�v�P2�4���9nk��`
�`��l��ʧfu�s⨠I���}�7���#^��p�[�C
��\&��69���_.n\ه
O�t��M����*�;��!�h�VW�:���b�J��S�݊dB�ٖ�+���T'���T�e�����(��)t��y���'�=J�S���T���+����s��p����Z�!�/�WM}�������`C$ۈ��Z��E�:ԕP(��?��p(?8�w ��<)��H�čBq�0
�쮚�JO9�C #'�(��q�R�gf�f ��*����ab��S�Z�A-����R ��ڲ�=+�!8+�Z��n}�?��L
aK�!��:������L��s.6ؾ;6_��7>����t��"i jי�m� �g(;T�1Q� �O��v��Sh�h���I�]�semp�6#�������(K�56~�����h8]w�n]E�F���邻�WSDR���nX����~�.]D��ǅ����P׸�ƬQ�	]�����x&� l潵�sL(�Ρ�)E�a�ݬ򿅦	��I�tzcs�r�3%��UA�	~#��tf��&I��s�w޳�����-�=:��n�b��>&۹N��x�(�vQp�P�c��4A9�}���\M�AQ+��׽����̞ZC��P��03>��i��"c���ф�o2:/�R�{3C	Z���r�:�'T���|������!uMR�u�\�\��/0j>!��-S�yx��l�\�@�"��$Uٖ�5N)zXIL�ς�%���\����ʕq���O&b`�_Un��V!���RP�|��6Y���M+-[�m�D&�Ӣ\�Ԕ��B����� x�黊K��%R�)0T�p���N�6�V�HGבũ�&o;�w�@��K�H�Ds���hx>�5��=4�Y���5�=L/�~>����*�}�C���ҽ6�"��[��&pjy�G���
)���Ǡ}�`���8�@G નщ��t�U[X}�3�8?c/,#��{&���PHc�7֚K��oє���U;��Y��zS5�=�s��
aA�����_��H!��r���e	�*�
����r!��ީw_N�k��k
j��w����װ��ʹ"��*������#Ʈ5��az�����~v1�����pd<`�)��:9��V�F�������Q�﹫q���ތc� b�jH82�����Zͩ� 'k-洙���
�Y�Oq\���%U)Գ0���r�`3RG��NL8�}�s͙�� �p���՟�2�?��Zֱ�����9��w�=�bt�U�@�7�t�	`klYszF��=�.�ԬP����>~�ћ�!����c���1��ն#H�)i��6����6�f9̞a�Ɇob�cJxcSs͚&����6�8��6s�����;����w1P{c���i?;<b�2���H�`�����t�6w���٢C͙����qN�W�I���h	B�D�7[��j��GG�A�e� �T��
��T�z�-'oHI��g�������u�+�6�]'�������$�&�Tܳ�̪ZZ;  M�1�O�`�!ɇ�=Q����}�3Dũ�*����"�0�A��^Z���}E4Z�j}�]H��,8�:�>uKܤ�1���clG���,�a�IB���$��@\SJ�j�g ���`2� ��o`�t�,��͋��, �؃jc"l��ѷ�5�T�j,���s��������a	���Va�fN�k@d[ԔA�t�F�Y�!�/i���n�t�Y�}���Bs��"Zyō�i)C�s��E��#;���*`(���8_8�4�B��Y�l��=3�� ����)�Դ��S��Qf=.��T؎���/a(
)�-;bؙ[A��`��m�U#$��\��]�g��SA��-�����e��phZY��~�i��W��ګ���ۣY��I//v�~[o��18/D4�L#h�O���R��П�XH��ӽ��θ�J�hD`���iʑ d���<�K�iJ�54 F�\�	�	)�OU&�3����%�"*�_{�w����S�W#���w��Y�᫭������ ���]��
{`�rl7��B�L��=b�Fv[��Rg�V���}��G�K!��m�pn�l�U؏�ϰ�ֳ$CCds����M���8�l��Ҳʡf7rz����!�\<�A[S�3�hc�	���?�Y�K,�O Y��ξɪ�f�Zs�{"ZQҶ��]��z��0�vآ_���G�g���G��-���v����v�a:/oeك��9����I3��59N��Jgm��Q�z�.��B�͉�	�@�c9[�H����tb�tf��6�X��8�:v��N�/E�K��P�i�<�.]R!�B[����]+�u�Oe)�2��%���@�ܭg���m�W�zUg��˫�9��LB����F(ƾau���	��=�H��r(:,Y�HG��<\��y��Ӵ},��<Σ ���\C�'��y�ZW��7-T �5rӑ�>�є��膓���b�JjZ�m���|^�I�7�& B�P:�`@y1O�L�Z!�{�������V�j)c
&Z�s���հ�p�t ��������F�����E� �~��^>�BV�
���W��D�̈���ǔ*�^��-�W/]�����=��,<���q��N�C�d �����jmzѸ�0���@��8�j����5�H5I�3t��R	3����������s�TG�j��g��YUF���*�Uu4�!��d�T�)P�ʁ���!��፹���A}'��<��藟������&�/5Q{��N[��������������h��X�7!|�C�u�&�EM!ɖP�����
*�*T
�7���h��! .$%Fj��`Q�iu���E���2f���U;=�����Q����*BT7yg�,���s��­�<kc�V��lnǫ�d� �۪�!�]7������O��A.���{dJh'�d;�����!:j������ӭ22�v~)!u�o���W�:Y��e�r)Z�T�*�ͥ�Z�g����}n�Q5��
6O�q�L]7�\��4���9=�{jwg���%/�쩖b�
cU�.ζ�Zja'xj��ɨא�\�zZ��3��D̫҄t�7�-�a��.���6��bR��@��wE���W�9�	�	y�9�uZ�~c��;��R����͏��j����|���y�_!�b~��ג��4,�G�iHتpʵ:�"#��@�^�j��8��D]}�`��8!�'E�?�Q?^]鮱;_xrS2�LM�?˳��`*��+q�ܔAƙ:m�A �L��y�>��8Vy�7,�� (���-�O�A*�+�SH�
.���!�������)�'����Sd��1 �A������xK�(�Ȭ�-��	Eu��\�ʍ�,mNo{���U��/i�p���kPxO��]0���9X��/��|uc���3���	�����B�{�w�W��=Z2�$x��y��r�9�£�!��/T�kp���7��G!]�� �$R� �� ��2hE�|�q����x(�����}�M߾���.�
��3l��T�hԝ�L�Y�Ok~�y�|����)�WQ��+����N3�@���|��� �	`-=2�!E�Hd��*vЖ�*JY�����N*�����/2f>���ON�$_�AZ������¬����"���?�b�ٿ�|t[B\�ҷ�F,we��"�O�a��r灋I�Z�v�~?�x�(]����]>���'�3���9�yٯ��x�\�?kP�I�`�Y=��Ѓp�K����
�j%�%=&�N��d�KA܍�7��7�	0�]��Gx��}���h�صnr��dLLBe��B�9z>N<��!ϓa��܉ �/?�����xe`��vP�O3�wă�?�-9�6:؋��J]�lIX����S7��z���,|\�_I3�0]��v^}L�î�`:���(ԫ�|,=��Z���$_���CM+���������x7�Y�<��E��_���~=<U�_�F���%�����o��.�"���lA��.���:�e�b�}���f��&�⶯�{6@7 �	����{\�{��.����R~����Q;�_���Z�9�X�g�D���ĸ�J�*�SҽV��Q]5����dg!��!D��b³<z���>��`��s#�4��j����~K�Wؒ�<Z�+�z �����C���dEk�=��a&((�kX�t��d�Q�����=��B�O&�����1(�Q�5���u�qX݆$ su)�"��f�[�5�����LX̚Ս��nP� S�U���SU�/���������K���:�=�	�����L�)�$nzb�(D�?�~ߗ��c&8�3-d�{�tV��<,��R�$�$-�P�xx�(����/����-͵^�ԙ�]TlƏ�yҝˁ<}G�=	JI�%�{kէ�����]Gs}�]�=�H��`�:3����`�7�#a� H*��_>���-�Q7c~f��A�`F�Z1��C���c����Z'31@ΐ��r�!�TWQ���g��/��,`ע�4I[ a;{P/�֋��x���� 8bs�8j�;�>u �6���3��^��B��_)�� X\�r4O9v���b�ID��BU<xs-z�hPW� �˫uQ+�n]⾫f�B'o�!9����("��爡<%3Wɬub;&x6\�h9i�t��Xht�����TH`vo�!l����v�nQ ?����Q�xE�Y��]܇ť��	��(b����EFq�?e%YT�j�`�O�fh!��7n����ι��o��BL����<�e3z!�q�f��71i#_�Y����_�L܁�_z	��g�M�Q�֏��7d���m��F�p��X�����af]tV�"1u��4�n�!�#C����)t|H���`(���l5N6e/2B`�u��3m�'z���<z86���uZ�QP[J��Wm��������˪�C1"4���B���{ ٿ0:�����V�o�Q���eP���]J��������+��{H܍o���=���ó	�I��w~�M�{�H�:���䟫d$����ɾ��у,h�1� ���2�U�3��+�gC&�����]-�崾/�}k�X�����*�/�YĆ��s.J1����V�.��ʅ�ǘ8)�6J�������'Aԏ�JGk�y�K����뱱9[��K��8F,>2J^��Q��P�v�����-AF���i�D�5ŷ�������Hl��/������Y
�U3DK՞g/9�٪��Q�~J=`mmFq��gz3$���B�X���ٴajJ��b�u7������cE=��i ��M�v��{@��;D)1���sB��,� �����Q�!���_��\���f>�{E��M�MZ����qx߭JH_��������у5׉�n?ݷF��Y����t[����bt�9uA�<6�N-HMG��#jF*�y"��2�7O$�KC����$ՔXF�?,;eR:��6���i��JrPڬ���p�aׅ��V_��o<\�^�{kHu�\������WgE�A5n:����ae��C�u��~�X��N.��U�<an!O��}�Bv�}��4�?�t�i��iD�>䛀��5 U���x�gp��#�E��S���h�o�~�2���j{Ƣc2��Z,����!ߞ�i���=�a��	l>���l�.�	 W��+�{���z42x�_M|&aݶ13��92�)>��Y��N>Tԕ{A{��+��$�Xjn5�������q�S$%��F�e�y6�W�5b��k���uZ_Tu5�x��V_��>�\�Iǀ�Q*S�{�ؘ&�:�ۍ;�W6�[�?�H4�,�O�@��,5k(M4�o�gJ�X��d[�&�SB]j1��?�.J�a�82[o�X�a�c3�_8&�G*L��5��C�f5�,8p�&{]�1��'t`��w �>X�W{��ڑ�D-%nHT`���XdR�N@�#d�8��|FM����w&�g����+cM�x��qxG�6�5�)%;�E�[}�q|����J�J�<�Zs��Iu�׷�2vX�44� u�AR��ь:hi>�c!�` ��Zh ��ʴ������g+Њ��0�95��u5�(B4��G���9�ϣS��x������lu��7zSx{��(]+G���-m���K@�K�VB=,���]�~\�T��~��cP.��&�f��'+5]V5�'Z>�{)���&q�D~Z�٨�R���(�>��h�AV���/����#�A�2yDg�lhQZ�r�=������*#��ì!ǖ�d�A�Bt�?L\IE��6������
yq�
�"��ɹ�]U���~CKXG���iܘ��_�=��`h1�5�@���PǝH]��yJ��}￡��>ٛ��a�{!��5��8��^/�!�$���K+poA��3Sӥ�������U�m��<i3C�!�U�ѻp���!3���u��N�r��J��9V��\��5̓R�__�8&&:{ɟ ^1}q���%�Fc!1��'Yޥq�؆/|�MQ��I���J��i�u�6aJTB�ܻ@t!K��ˬc�o�ۺ=!��[��J�?ı��H���_{��j��.7v��ڭ'�!�¸?9׎�kxFv#!`=� ҽ~�t,� ��l�i�td`��Ҕ���v9�I��]���7���\���!7l8ׯ$�~���^��v���:Ș��Om%�d
�W�|��������dOJ�A ����r��P�S�HT��Z-M�Ѿ���as�wٛe��?{��8T�c#Wʿzw�Y	�IT��ȶ�Փ����f��l�,SxHvS�nb���l�x�J��Q ��2�t��ꤿ�#�2]�.y{�dDˉ�>TA�d��X�~<����|�<*���u��61���AO�9D	L e��b ��#���o�~/e�g���_/ƻ����5?(�� �A��xF5���dt�r�Q�J�)��gG���P�H3����f���/#u-���,�t����wH�fˡ����<�h|rZ`����z�e6�=��
�\QA��s����#��W�6���)�x>�p�� }&I�0e0�~H�E$���qB}�rD�`Bq� �)�}e�酙"���p����̥�HeiU�6��l��0$�����"߸Vp�R�����ß4��gW�?����42���zn������XB�u���jul�Hz-�V܌�%�7��W�0fc��O\-��	���:�r�6����������HT���Q�?f��� WMzBk[�?�qt����z�# jp#b�7���S�C�s��&�
gE�>rF1Lv�g~<�7r���=�|[�:��W����9�~O��ؒq�.�.ĳ�Z,4;[�\D-��f���Wn'k����ǭgݿ&��
?5j ���bWmA�'�'��'>���p���_p��d$�zE������g����_�f �?w����A,�]���w����)�ъEhwG�k#��ac�	�yD���m��d=�/�Ѫǃg����S������4<k/[�̣�Ƀ���{��m�u>m���_���q�'�T���e0�xy�R�'F7���ȼ����o�L^<"�Nn:��|��?�C!Ą�bt�l3�1gJ/�r�`"[�:8M��J,��.`C�u�:�cV;�nv�`��%�����Œ>��5[�ZNT֮����,Fy��sՊ	�Co�y���-e���4j��:ѩ��S2b�e�q�����1��&������x����\2U��N?ٴ�/�ʓdX����`��r�H��Md�����+�E�����H\���.ö��փ�j�5���!�7��l{�vz��'��K��_���3�
���5�큸Y�]é~�ų@<�?�$�6UP� oX����aڡ�g2BdeM���Hߏ��M�A��YwZ�5�/�M6Y��؏�'��Π�)�����g��K�kb��*��@�X�hYS�\r����ř�ޞ�:�DA�̌�����m���.���n����Ʒ��^E�JK�Nq�d����/�Ywwf��ݕ����c��@C���Ir��� ������JS��\qV��i�7w�Zb7�v`-�ͥ��@�}�K���q}���w����]��r۾�-��b̊诼��Bݭg�ܾNf�������f��] c��O1A�Z`0���I�!�EA:k2ǉDg�>���R�`M��ho$jWt O`A���](�E���,��̄��f�~�Џ��Z+�>��O��hQq	|�/�+�eo����,	�;(JE$���B����d���6��Q�8�v��D�D�؛�_ubK��<�V��VD�b�}t�Zf�^�|Xe���%����_1���mذ�΍��b�M�����j]�~�Pұh�}PK���V���d�]Y"C��B�*qd6�[�5�^�+��0C����v�H�aH{�Eg��D�`D�cx���j�7�ǡU�w
C8^꟠�t��-b��p�ՇR�. U\�i/�Y[�<�N�\����,~t�mfp뢢SW~@���1��`�!1��-��Ԉ��m]�+bM$cԴ�K�'f��:��ː?0�^ݾ�*I8�	%�D���ɉR���4af��,[1�l2���J���	v��x��L.�_�b�B���
�)�d-�k7��q����/qޣi�:Su�31<�禄�/���/r��)�*�F*��Ӊ��c�f�4�dK���|9Du(��'�p���g�V���C<
�%g��j퀪Onh[��A@=Ey������e�M����:��L��E~:�z�/1��s�
�)9�dNگ�S��iJ?nIg��{���<�ۂHg�LndS�o0��bg!hh��8o�z�/aȨp$hs8�Z�~�S��d"|��N�EP��V�1���OV��Wx�d���z�L�Vn��+>��f�(�\����ULr[�A�<w5��
������V�t�n����O6\��MAr��0�((���S]-JF���f���F`@��yf��&J���v�����5��Z�՛V��1�k�_�����R��V�Mr5\���Vu��~���;�2�xb�����ԭ>P�D{�,ߏo.�B(�ZF�S��tD��:D�=tr����.R_98Qs�J�z-��I�D"	�H�X��	?������C�J�tv�@�.��#x*�)�R��BYJ��ع��/�����	��cч�k�ZM���dq5���n !y� �lIuާ�����ގ��O]OB*,�$�i���Ȼ��o���q�eB�z�;�<�6��y��E��^' 7w���
��?f�e(~�	��<���_~��lRx�{=�D�d�PՂ��������E$��~N�&Q0�k9i�V� =�#�44�����Ѳ��4��������w�N���zc�W�A= D~��.؎��|àzi,4�@,l˳,�L�c�=����C'��*5tY���������6�t���|��8��'bTݲy�S��VcuYp���|G�A�A� lhf(-�ʹ�q\���_�DBv>�_�X͑�
ѮD����Xg���`�D/�F�MG�//kX_���Z
ꇨ�F���B\�N{�����vF�kRw�rf�$���覛�oo��-�J��"7�ɬ� r��H|Y8
�2$i`vZ��:��GWحiYp��
΋���Ur�����2����WP 7j��5.ғ!HK?��Y�QH����)ӷ�{����R%�L8M���4��;���,O�R��u�F������:}gYӀC�G� P3�[u7����)��=���w	�H�q�Q���~ݲ/�!�=9� /4L3N4�G��=�xL�g�s˱SL��[Ɖa��r��N��1ı�u�OFuO�A���9��J�0���=ݰ��X�ʀ�;HG�.���	]�U�z�}���� JӇ�Ց��a��u�W�
��/M��9d�3Q�6$8U���)R�h�7Y�.�m���)���W��ď��aئl�{����q%h����l@1mh^˶2c�2z��K��@���#*�?���h9�`�8ek	$[��[��z�/+C�3D�+hP���H���R8�T�F���n<��z����GP6Q����Y'SC�D�=��L�@��Aő���b�*ng��M �����jZ�?�X�z�	v������jy(<%��=��7+�6����"n	�����Fg�/a��h���s����0t� 	ַ�+��*X	�RN�\�"c��b�!�L��_��Ȑg�"�M��aM�,2p%A[B9wa�-lz��Uׯ�äP~�L%,Z��>M08�J����׼>غN��1�-E��ް�3�9�q$��6��}Y��1g3�q���Q���