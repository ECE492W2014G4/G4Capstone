��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|��V�^�Z�4���%�ڢ�kU�j2��.��n�{VoR�.���g��ɡ��80EFj��ƕѻ���vBͿA���CeŢH�y��?Gɻ�+��aFqB��X�ذX����D6�y6�� ���Ȼ�o�+ܚ �'�J���ڜK�]?�]�ك;!�Uۍ�j����Zk�b�fE���c�;��m����;]T{�i��v�QN�x'����j�B��-b�V��{Z���zS�uOV"�E�B�l���i����6 ���$�N��ۉ��&?����ؤ�1��*;�L&h��aD��l�4V1%��3�����i����'��O�a�:��n�n�*��B�P��q\�m��^��^5����H4>e���R3?�с��b�"��5f��Lz-Z���"꿚#_�~��\ZY���N��_ݏ���(��h�{`D����rO׺�=�<���C���Ԍ���,�#�:}:�]�/ԙ���Q�%/9&�\ۨva�'��v��+Ϥ!<^���Ыm��
S��t�B��g־��i��T>$�o%K��F�`qd2���Z�W��+�&�x��7Z�X*�A��
j{/K��cx�M�$��F��� '�|I<��-�Z4"�z�s-1�\R�!���YZpJ��{�C1=��&�|1��(_n"�YO�r4k��G@ܧ�Q�ՅX�����oI2����{���X�i�+]i����l����ۚw�G*�>SCɮ�󽭯���zI��ƍל^�@CP���X�|��2Gmq��S:>0��!sB��d����b+K��A�yU:^q[��NNo�ޯ^�V}��HS���d�NNU@��t=8 �؟�ZQ1��~�$�b\W�A<s�����/���T��E�OOy�y�l23�(�o��ٗ|�_r�g�׍_��iIC�v8�e�w� =�����-{��W�o����������O)��k��$^�xI(Fe���|�Ä�؛��L-�Vx��q���N4I��zd��4�qEE؋a]R3�T�#�պ�1��q=e��3l��􌌰�+�ԟTV��×,�S-/S�S���.,�����Z�&�by��~�G��r�7�,��TF�D�Ta�-k_��m'�N��L��!�r�ۘ尡��kf��3������Xl�c�{�y���A3�V8<S���U$�hh)��ӖN�:�Z����ݘ��Q���]14�*�1XJ��B����ĩ��{�t-6���q�P����C]�h�N�lq�84���_X��l��Y�l����ϫ��FlK�e�:�N%45rIQ���w�<��|��S5-6D����ܸ	��_���Q��R�F�!ǔυ���3dy��|�n�c�ԁz�����hV�7�I��D���~�1�p���.ׯ�9�t�K�L�;4���oB���{��B�#Qmv70���,�x1�?�Tу��L����nGR7��z��i"�ެY.��G.KOGn�)�I�����vM��8�����`S���73|]�[�c��B�Ղ[����X��r�s�UCp�>�DH����̈�w>�&�^�\eq\��C`�V��idp�jn��=��	����B��	���Ss�"���oEZFު��)��>Z�T��e�����K���+=�
n�z��q�@�ա�<���a���w�jU=�?�=�kQ~搴(%Π�i�~r�U{#�w@a?@d{�D�s+�*܈жNk߿|ܚ#m�}��U�1M�����p�Q��Hu'�tT��'����Ct�T[=��+M�8�S}��</a���<��x�|ϝLiC�<��S�
 n�uV�1����;
^3D�\[U
&�]�1m�	�I�4�l������5i� +���;C�����?�}柦���Eeϸ�R!.]���T5:K��u���}����t֔)�� ����-h����]^�l�]���f~E�GB��+b���(Lb���9�._�!������5�����TU�n�,��I�$F6�sI�%	2��IKH� ��'��0����\������B'Q�Ẋ���e�͂�C�:/*F�Zi������h��xl��f�2د+��3��t��=�[+0RqB[��yI��N�	`�
��wL���_7Z0��<
}��5ǸHa5�=��5�1������z�}QؾR�=W~��m�U�}�Q<�aq�9����CB(�u�[w̏g`bg�)��W�	f�*r?a�g�N�P)	l��D8]�4�0�1z-��W����[�_<�J����g;��[��7��>Y	�=8Y/s��¤�ۿ��&Z�9���^��c�nN�!���+f�6:�ԑ�(0���ZB�d���x꿠LT5&��-k�tQ��=.�e"���T�J@}����,ȟPȨ��1��y�]�b�&ف�m���椘�����Y�n<ў/�?D.��O=�촤��s��X��e�������~P�s�ϣ��jf��}���a�]|���4�?̗D�d@'fl�9����ys9��߼�6'�Omo�=�p�q`{���|В7�m����c���_�Tv=6��1�U,ٕ`�����m�Œ:}q~���{�ڇ����H䋽OߣY�!_[8O�M��ȷ϶'�z�N٨ S��o��D�����'�f@���R/��K� �����cQ.��f���}��^��;��:s$@��+ч�1Zu�os�7z�F�]�4��}T ��#���M)9���>�#\4���Kur֍(ׅN�l5V�G!��z�G����.IKU�;�v	�w7�$$m�sZ��[��k�ZY���"�PU'�J|�B� }\ݐ/���Z�;g���ټ�!d��i _����25�K���j�j@�Kf����O�w��tR%���E�y&ޜ�t�.�K�hP���}]�H
��ƒ�=jt}C�.j~�� ȃ��;�n/Y�LĻý1׺f�o2�������;���e_Jn!�ڃ�5!���R%�׉޵�l�
.�s4�ͱ��b'��-,i�0�?�밳�������zm�@�@T��@VNQ��&��s���sX�%�.l�/T�a2YR��ѥ.7sό{"l{[�b'�8BtV�b�$v�+}$�7�.`M5�Mhp�G:A�`amf&^M�=jj�\���v,"�cI&lZE�g,Jr�!���,�&S}��5���-8L��C+cQ��'v	�|�bmdvU�'U#�x���.���ؒr�4�@.�z>��>=O��5��?\�]�gT�8��!,�vBD�G�&��-�Sm�#�e�#�R�4� X�ȏ�9y��������ʹ�F�E�l`�Qh%a���\֏�[��R���@&3Z��N�1��|�玚��"3��*�9	��[�_�ˊ	:`}tH�ǁZ�0_*c��BG���C���I�n= ���ߍ�I�TS�8��Ub���Cj���^K5n�U��#*��)g��n�>vp�����rV�l��֭�����j��y��&|��e��hv߂%Vmk,�s"@��`6eF�F�W�v[К�������&[���F�=�N��h�N�_{�Ǝp���Ĵ��t�����Pz��Ǳ	�R��ޣ��nG�8t��բ�4�a�	����`%����Q����?�+�xv���f�ȝ�EO7Tl�p�Yܪ�暯���ZeY o����\C��v�EMC}�ϧ��1��!������<�g@0%�<S��=�,��y�Ι�#����{�.z:�J#9Ŗ6�el��j�b���5�A��ڋ����I�_1Z
���JZ���/`c�5$���y��K�})Js�큿��@ȃ�N�T�~��	����=��Sq���Ә��	>���5{�ɢ�1�C,X��p�ce� 6Z�j����k��z�قj�&7pA�O�g�����Z�x|W^l�����N)�s�����WUՔ�A��N�p�����8���0��JZ�T��e�|lZ�Zuj$
�7���+C�W$3b�v��:�P=���`K/��N��p��s�0h_�V*b�� ";lA_	���Yz��NZ���<g[S��&{����4V�H}k;c��15�:PH�Z��l1��z1�W�Ab�i��A�bd��q4u�h��i�3�8�f�Dɯ�7CL�k�)��z�WZ����L�A��g�_;08|A�8��x+(n���Hhy.ӳ�bze� Ov�ciVq��G
0�)�d��L�4����
 k��H��sY�Y�3�݊����7�B�Lޤ���-W��6�XM�A�����֗��š� DGEF�-*��q�z���z�.rq^���4"���b�(�����y���X�3�r�>�!+��Z�_-w�s���?4�)��d��3�\ͧr��k.�e�F���*�j>�&>�źuK��6\�9ˣ\=��WW������u��/�ț ��eՙ�91�c@�M �'�h_&k�������w2:?���K:<�̎�Q M��y�{�DE�nO�b:t�GΑ3��Mm⾶Qf����Q��
�]�&3j#XrV�Y�z'H)���x�r�7�O�&��}8ۮ4�����2�E0Ǡ���B�Cr�\�שZ�R������]/W8�?����<����a����0���hk��`	;'ra=3��3~]脴�kN�" 	\���4l,Sl����:^܁~L�8�� ��T���5~+elX-[�j�4�SӐ
�X}�x@ۮ��jv>�*}�w�4��W���&�*�#e�&"����wt����z7&�5D1{�x��t,F��n~�A沙o�)��Kg�"�Y��Ϊ���đi��J�!5�+/(hK� ��q�%Ih�?1�<K���*vQ�FQ;C���c�%���yQ��T���B�	�B�|��k( �9�����h&y��d܋3��#A.B����Հ�f�"p&i�~��`Q��H"��+�����H�U�����^Qj�M'/dW0m>5��1��>�鏟�E5a%:��W_�M'=��J�.�$k.�A��_H�Q�"�@1.��"�#xn����H2�ig*2�d�A�*(�����>xi�[�M�5�HoZ�9zM���f!,��p��+}B� II�5�/�h�;��
��c�N*]�c�����芡�dx� H�0ʢɨ=��њ�O�� *x�6?�	��Q�pԫ�Y����l���f�b�;^�1��rm+˥T�X���ʠ$������w	T����OS��\-�a��e-��N��i�]|�1ن�R�y�iv�(Ê
��Y���K�B�Jo$-WOz�?������s$!x��:;}�~��V���ejP1�����]�A\�D��O�A⡕1��{¿F��0�r���U'^��KMܲ�u}�l��Uk�nC��{�H"��c�OHp�v�e��n"ٯ	�4����sT�������$��m�~9�#5�[/��p�]�?D<���s�g<a�o+��;LD@62������b*�����=�ZʒNjlG����S\s1�m#�.5���M�Ά��K9Rr���JkIU����I}���������RI � �n�V�C�,�~�Ŀ���97�]�ta�^a��㴧g�7FZaw2!�	�p*g\iobmu���:���%�`������G���]K��x���ǚ{�s8��3:�t�v>a���,���5r���
�V�W���\`���٠R�����a{�B>�Ou�s�{��95G�oO6c����lW��=��y
H��j��`���T������=:�}�
ut���E<�픺�\�ؕ�s$��s�yv��H�D�����$rO�8Crb�����팍�ѷ?�*�G�f����K	y\�B��|V�R�Q$�ffT��b�/�3�i�o��w����aފ��ܑ�=��}į��=���k��������	�E�XtNluO�_ �x��XT�T�Ǉ^dH�6�k��
�����=�M�N��^�cc>9ػ��tȆ���%�~�t���%�7�ԽF)�<�8�E�{GWL���;6Z�������H����O�ƱU�=̆j�؊!{&�V�M`�weK�c�Ef�W��\&1����=��8Q��U!���)��z�&S/�/���-`�,�13�j��,!���������D{���5��<���
28�:��3�S����w�F���n�U�8קڽ�K����#�p�|�]=d�ޓ��Ń�h��i��9�� z՗;�ՂI���B3�qڴ��ZU]#�G�ɏ	5f,���$���4���i�)0Ԓu���"��P������.M����S�+7,���ӇJ��?��kC=��������CX�;L�����nwZo��F�g��t*����An]^��;h�cʷ)F����"0�{��M���OK]c�_A�9đ\e1^���Ż{����hX'j@�d�կԐɰ�;��zd����7�mg#��Cq9)#Mxؒ�*J�뭭[:��-�O�6�?�n�z8�R���TX�)Z�����§S1/As�@���҂M�}?.��ܓ� D�^OU�L��V��1����r��F�f$����X��ѭ��Z�)Ǔ����k�_(럅���d����Qܠ'�ZLE�X|'b���\V�J!]0�!��5s�ͼz5��������ɗ�����嫾���S�ޥP�d��B�5H����Z 8�	�%v�1O���s�w��l�/ȑq�c�yۀ��ux���E7���DK7+o"��4��v��ꄔ 2��Iv{frNN<<	��L���:�X�CQ! �u;[$���V'7ʒN#=� �m��X؉@�h�[��9��S�٢���=�x�`UrG+��|��}l߉��J��6�M��߁�`Ŧ�E�*4s�)Q��^Z�1~Y�0o��`�R_t�?������VҦ��$g+�}�S׶��mb�4ԟ���~���7�p�s��0�.��� {w^����h�5�l��Z����г�4Ke���oΎ���d�nU�lo�*Hg�ۆ�%�C��!J�W������+�,aC��.X�<�CR��q�ť=��*(�~�8�i��k�7�����ܛϭ�yC1;ȋ>��Џ��cMҌ"�L�Z��c����K|��V��
���'BDX�G0���F�k���ȴ|�xف���FD���1��E�Q��7���"�o^K~_�B�E���lH��.ا��]�Bߔa�d��\n&�w���8�~��"�x諴Wk������<�s�z�ʐ�|���μnu��9�apWt|���NP�T��d3˓��/Jܰ�;bkj��@B?j^}��Y��ny����F���M��S��;j�c,6U=�z���@�ǝH�{p�V����4���I�z���(�A��1�����h[r1�o��	#�Tߥ�xC�zi��(3Gh�x���	ٌ���Yv�"�(�9H��#9��C����l\�-�}{�lڌf����>�N�k;#�3"��2e3ymn��Ʌ�j�k<2Vv����^�Q$u7��铭���iZ�/Զfܻ�(9�� �`Y<�0�H�ɥ�$f~>"&��)ō!���R=X ��A|8&|(�~3.���89���k�)�@l�K-�Ĥz�_ #�u������o�7��-��;5���Q�`
��2qؒ��WP