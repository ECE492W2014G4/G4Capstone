��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|����z=+���v�����p��6f�z�3��w��g��ķ�H7P�\Νg*�.�%F>�vg�Ԣ`͙Қ�y��&�L<��Đm}x��(�di��N'�K�π�wգ&��ݎ�30,pŉ�$[�1�5� ��_.G/4�w ��Yʖ���(�E�T�OH��cN�w۫��@�oQ1,q�8a�R�j%��j�O�=�29���`���X�!�m�}ͮ�E�L��Btr0�V�[t�c�� �I���"�U�I~��I�u������m&�1�؇�5#&<\+�7Xi�9H@�y�^�n�1(,�{����Aǧ�C�vP�l�AÅ���(����RĿz���:)�v(̃j�'o!(�/�y ޹���7�#aߤΕ[�[����|��'�����,/b��I-K�1$b�ĭH'���� �*�'Y��7(k�sy�����R�=
���Ӵ�w?e��9:�w�K��-��+znzau9�fQ�� ֿP�>��ykf���˪���1��@�R\2�$�*3L��+�?�zo�fB� C����r��Q��54���� ɨT(�3L�V��9�Dݍ)K��6�"�,��~i ���x@�-�A6����������/�߆�岱j�8�90��o���tH�#�J�cW���2-��"��͠�"���@^�O	�N�+�Gt0��4[��[������5� u[�Y�I5�{�V���)E�C�e� w���9�7�s�Kl�h�=�$2z��D%^]����3s*�O/�(��Q=yAj�H@H�ƪ���tkÚM��3�}H,��)w	,Ji�&so���̖*����`�@jE�#�.�C����[���A�Q=F��x��k.��Rf�e���������T`T#÷�@�K%i�൩��-#�E�r���_���'탚�SQ�^������of�����:�%�ܭ-��ڦ�='���0�G�C]�K�`h��#Ufw��b��b�f�ܙ=�qH�T��2�G��wQ�fYFi7v���C$t�;p��&^h�ϩs���{>è*��;�j}�)�]�"�Z��%T���z1�Ն�}�$*)�o�x6j.���zH�4׹rtoh��q��i_��R����"Vj��� �'�)+2�Q��J��4�cv}Џ��w��)	Ŭ�ܬ\=�!bu�u]�*�_gV����y]cn�=u����?�\1 x'&i_��M�����C��̛�. �Z�Y!�\
�c�?_�(�4����F�F$m�(͌Nzu�g@.�u�m�ݳC������S{g:��s�F[r��K������(o��hl
+�yMq�.7ad0��Rx*W�'S��V��h��_J]��A����Pn��*`(^�1�(*��3�ګ����(�΀%C��#�"��H3`OJ���j3��m�����LUȰ�T��%�yvvx�<1�/ߤ)�Nݕ�ڎ����ct�$o`_�O�7�)i�u�ѓg�m��0�n��a>��(�X6����L ��U	���P����Z��c�B�u�q%���k�JPՅf(Ⱥ���s�؊��|o	�/�d�	�&�j�Ի�
�����E\]�������[)��Z>��Т���UTs~Q�mK�Z�'�H:�Qd_�P�77�%�uJ������:�����<7?ɏh����nh�0�@��_��)�Nn��a���7�H*��;fKW�m�c��u$�bg��#�3���9>Eot��K]r�lrB�5�m�}9G����6 ��L8A3��'�P5a{�=:K$@FcE[���W�71c���j8v�侎� ��<�	k��,�v����9�eR러>�>>���b��C^�q��%���4t���������V����p�C���S(���X��ȯί{ /q	\V�W�y��RC�ac  ��v�F=��<��IJ����5������`���C�͇(ݻd��oN����}Y��5�w�k9�쥦�h�f��SC3�`)*��r��/�8����Y=d,GuB7\�(}�%5�*�sO�#w*��<G����Yc��P���A�t�a�z�=��B�w��\?��B"���Y�H����Ԙ��`dQ7D�4��q�RHy��
ʗ�{�d2�X���a�v=[�(t۽���t��x`_�U3���zv���A�������:�s�XE�n�|]h,P:�&���+ّ�F0�J=_�v�2�si��!e�>=�NH:�^�ͳN��+��f�ܺ��M���{c#�"�5�a�]���@�>��ԥ�<3C�ͪ��De_�N؃�#gL�Ϝ�R�>�""�ړ˿x[f�*K2���^���Hߢ����l�C@)��hG�H�%��5�y�nB'����"�sf>s��D�����
bX�D��\(/�X�zu�%��U�l�`H����l�� C:A�'"����m�Π��?bM#�z������,��g>5����nZ�,_�����D�e����L ��ܰ��Y��#��L�4 ��Ѝ���܋�'2I�<X"~z�;d���D����[�J9�"��t�"G��1�۸0ka��;����
����.�&���p
܏L���^�<Z�X����u�,�xd���%�B�^&B�A�\��m��2��] ��M�c�׭��ؽ�w���F	��T*=��{�{Ak+e�Uq��@�JK��(~�����1F0��(��?!�C�NR��4�:���tin
{Y��iȸ��f����r}��#�>#p�`@_?az�/�@t	���[���� B�9j5���%�e/^#��}2Zu�-�+�H�8-�Mи՝.��,+�2M1Oc��PΪ�ݐ�� 9,����WA�^���vמ���YX��p'dN�$����	�$jȡ���;����b�N�6,P�R���qF�D�e���G��sC��v��6�
Os"GbXW	��^n�y��
�R��C=ݨX��|���6H.i�sQ(?v'2S��Q@��nJ_F���)�]eϙ �
�*�]U1���eց�(��9uX�h� I.�)U�Z\�]<��>��k�+�)�N���99�JsT�dLd���f��E��߳��Ь�e��x���vp�մܛ��25�#UW����PpޡTd�ɋ�$���ٿ�KalK���ә����Sjj(�?�1�ר[�/�g��-��IyPg����qz�5�li�uӷ�9S�84�z_A�4T�D�pB��N����ǋԸAeNS`|Ǳ�B���QC��j4F��3%����@��-�������/K�n	z���%w�5Ɩ�p-J��o�5?�2�C�>���I��Dy�e ���l0���<P�3v���	!1�ܞyz�)��&�H��7��!U�X7�^���'鱪�ڭF����7�*(y����%f��,N�Ymґ�F';��)��*U~&��B��iJ�ox;szO!��)yED��k�hF*Z�������?DR�HQ�$`2�*��7����j�Oʱ�̎�~���ҋ~����q��������^�6:��Y�RB%mܧK'�.�o��e�^�;