��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��/��Q�w���a5P��B�~�/�'̙���S{���^�qѝz��'�hřD~dVr�F�!5�=��[�\�bYzy��d�(5���*���D#����=�6�c�p�GCE�N��+�xh�Eaa�Ƭ�z�5>��>s(�oƤx]C��F�i�TϚo�2���E���W�۠N	Rw��#fa�E����ǁ'�iM�$r����?�W���aݒ�3��L��'�ފ�q��p��FU����vJ�k�~���l���wFpe [�29��Zq���)Rq�� �CPu�)�;��/�V�2��'cu�*�Q��펊(�Ľ�|�3ڟ����<�0�D�>,�n�i�63�'�҂M�N9���Eʖ�P��5��bG��̆�~��ܒ�sH_͔8H�e�\7rt�9ΝM�O����0Uh4s�{�qog�J-;�+&��G�h�-2Dro�Z�}=�r�WL�K�\c4�]��v�\�i������K^�nr)��d{F1,	bw�h��H���H�tU�f,AF��_Ct	I'§�y�����Dz�H�QVsw�X4!�b؍�,��9��r|�B���p\h4���%�K�������_TH��^g�e]K�i��U��v��ķ�]�b��.� ���`��&+����*ɹخ,�5Œ�?�r
���!���5��~zVKrH��D�o��n�Q�z�e��`�i������D���ފ��
��~�(��>E�(1��㕚�(KE?(�K�����TC�δ
�w����A֔������ڲ����s>H���� +d�h��"Ő�-h���S�ώ��.��`�t�j���ݱ���<� ��wd���5�f��ۨ�4�Vl�Pao+.�kװ+��fF<��NuPȻ<�î>- ��D82�Jj�48�T:(�b���EO0�Ǌ��������J�`���Pp�Le���K5��F[��J>�����}a?��B��?K���0Ki��a�|~�ڑ��P����^�w���}�yjƐ���X�ge�����}�N&�����. ?u��?.w6I�Z���M#H=�kq�[�,��P&#=,��U��I����ii�`����8�a5x�W�XA����v��p���Dz��x�$����ť�{I!h�6t��A�x�b<��.���QB�ň�n��
�h���<��>��3��%��ؖ⒄A�a�m��2��sq�,,�m��g��y`��B8��;F.��f��.q�|�Ҟ���u�2S�_��>3AL��H| UHk��:ad#=����i��91�j���Ȇ�kG�hJ�Ze��{��r�DIۙkD@��I9��:?��Qge
�p�&�l����A4gWpr7��@��Iz��c���-M��zgo�"]�&�D�k�^�q���I(���	�[(���,�ll6����5���L�b.o��&Ň�E���:ǝo����͂��)s��?�f��=����ɦ#������)���ę(�x�zȮ^XU���fNY�ė䏓Tx|��-A�v�� W�ggs��wK������� Z���]X����>����n�36��eMz�渨C�j�� !)Q!q&�g��ȉz�cBv$�$���󵏛�o���ٿ�"}�i9f.n�*�6?N���Y5<��Dj���A���%6�QU���,��ܺ���֢W��Z�'YF��"���T�j����O;�4�Y��!�A��9��k�wKo��ǵF+u#��AM��;ڭ'"�H�\co@8��ى��֒�fڭ`���T埪���x�+4��F��3��$k�F���?��5��hQ�1�%:��[~���p�#�!��Lߝ�����ƸY2ʵ���,7��ǥ�]�E|���=`�]Xx�/�^LK�TZ��z�ѕ
�����v�;K*���j}>��C+H��+�G-����#&�&jFɿk�5A�α\I��!�����]1�bX�(�[��	=F��EJ��?~n�������n+cG���$s_��鮩�����*<�h�Ūtp�VD�Ww	�BmfR�Nı9��锌s��ocR�����cU�Xbodq�Hz��lw�I�\�!�F�}�?{zk>����?�Ų����Ҩ��u�����u�� �#��fn0J�AIc@)y��������v�gv�Hr��"h���^�H�Z�"�9s<M��ү5�i��)|������`��Eˊ�d�h�<���1�j~B���K���gd��r�~�O_�]���mұx�#�*��֪*?�&#�o���.� ~�S��p\��Q�س����w��R�L3*���eLr��'�|,:۝��GO¹=��
��@�Z�P����-d�:j;`�Jb�$��_�(�G���[�ɷNdM!�x,��5;єG�1��7w��/�4�Bs��!�f���:am���Ey/�p�n �  û�#H@��s����rV����{�lw&�D�bh��\��9ZgoӵU���7��8t��Lz���J�e���b
����j��	P8��]U/�&R�8UH���D� 6p�G�a+���E����1'L�n-i5*�Y@�T�5C�%0?L6D��4A����/+�l�
��ǒ�����gx�������T0S^��k-z5���5Q�g5rR�"� Sf7(�=v ��ꥀC����߄��/\��xz��,��Ug�i����;II�C�y�ǽ(w�iV�#�������B=��	ASL��	Cg���CNX�l�O�w�s/S����I�'�UɐA �w	b�u֖$ڻT�!�P�닢�Ms����>He��"������5�!c��vROz����?��z�k�gnc6�n��J���2�
��/=}%�s{���30�t������ыcq�����x���K�jX��pdr���ƒ@J`�Gx����J�S�m����ot=�w#�u�i+�d|�Y;�}�a�

`��C&����̔��;y����Ƙ�E}������<������V�g����nԖ#fwit�/|V���=�&f���폿?%�
kAf3;��2�m��i�]�
7�(��ċ����{��)�gKӏK�~�:����O���7f�ȵ�Ԇ����6�'����\^�p)���>���Ez���'G�N<��'�捕�̻p; ���/ȱͺ� أ��=����3dQ�)�zD�x�¸�.���-���Ϙ �g�;EZݬ���_�̱�����9=���~4��1�
����%��x���K�fG���z��i�l�݀�4Ny`'h��}R��&�딶�$w;?�$~ƈ�	��Y�.�#e�K�x
g;��D;�x�ʊ�.I�z�{���}k�mS�9U�!�y� �}�l)����3ˡ[�'#��\WTM�7�*�K�j�9��/��MӖa3XA8�7P�̿�n�߄�ē�\��kv;I���n�`?��dnK|vd�ڑ�m�پs�@'�:�ih�]���VS�W$��&-ё�UD�]�k�C�8�O(������$�Q"^����I;!��l�i�7��f�`gS�a���C�YWd��0�WX��DƗ�}�2 �cw� �����s%PH`�j׌w��#yK�t��iD\Y�<s���;f�S1
C/4z�/j�ci{4������Հ���wkB�C'�9Nh�E�j�uG���{�5�.
�9�X��\�˝��=����Q]t��m@���Q�����S@�]�J+�!'0xMx����q#��Y/Z�Dw6���m.���^>�1z�:�9����O`�UT��;�^G�7�?;�$g//	�(���ӛ��^�B�P��=�̺�\�?�\��bME*���*���K����9	��pp�y�~�uMdu�M��� {Mj@���1�q��@w̽ȬZ�W�uG"�p�b��N>�^k���b�����{�1�*2?��� �v�Z�6��b%z7�� �z�'�4�'7�d$k��0p� ��%�CS�H�����Φ.o�:`.uA�>p�l4TU�8;ځ��j�Q��n����1���>Am iG�v���wDڟ�s\o�4l�OW"�ܥۗ��y�F�ǚB
R ���1��������G�h�"��+��P�~2H���õg�2�8�K����r��K��Bض��Q1���=���[�!����&����@�P2��)S[T��x߼~��E�*�Ea�q��3�c��.¥q��ϸ:�0�7N�!�U�.|&�x]�CO3v"�a��os~ZJ�s4,q��,a���FV����S=���U�v7&�j�i{�v�E���_�v���
�6sI��[��n<@��-�����*��Hې�h�@IW��Ju>� \�9���J@MV=2p����`����~1���kU��9Z&��V��)D���l�)�����VCDS>��. �.��ݮ>I��6yf�R%����5�-7n�ٞ��9#���~����'����"��$	s�;!��,��U'�u	x&y2e>I!.��phg�X��ϭ����V�h)��po���Ŝ�{�j{�\c[q��QR��3�}Q\{�~�0���(��+�۷}"�\m�'[X�^4���m�*�R>�
EB!�?��3B�����#?��B}r3���9+RV��Q�u���Zb%��~��Q�LkE�������O�4s@��.�@����0o�tg�Oy\�+p������!��|0�ۊ�ǈ=1$#�D�b �S�]\�3s�=s�ZM�A�c�c�qf3�Y��Ժɳ$.y,1���R__u}��N�D!��pX��^�1O6�{��x0-�7 �X���*�#+��
��ޅ=�t��q� w'
��R`aH!Sf�p'�k�N��� :��cT�Z��QhA�_*��F-h��H�h�ҋ�v��Y}	�σeE~��E�P��A�7!��d��W�09��c8ڝ�T�q��w�l�۳x���W
n���KB���+�
E���򌮪��4g�HrĎA��V����4e�ρ���8f�kΉ��Xe�w�����Q+��$��j? h��ٕ�:���ƧF��c<hy�?U�!���F@^�ă��?�w�
.Y9�o�ړ�pU��Ǡ-8�L�IDV!��sI���[PäڐF�O�X�*U��D��R��wpі+~��0ҷ��:h�;~�H�q8|���EB���5�òa�t��M���z|�� ���o�1)c�bo���(���U�f5e%�jc�-���u���C��Tu�G�uݽ��®b�S�A'�X]��A�Y��-�k�x��V�с��/.�;�;�}0�Pm�K�f��߱��u:���<�7�=��dw��F��nA�g�R+!�<n���~Ϲ��?��G�x-��G$�lW��f�3��\�P���D�&G��N ע��ͣ���>��rV�^���"�3�Rl���y��V�;TEKӐ�ᆗ�]��-v(�j����x(���-.��H{� Ry��>�Q<��R��[o,� �Q�ϊA���s�T�`� s�_���6�k`���Ψ���wHT�6v�@2�ޑ`�0d0Z�g��l�9�Xb�V��.J��.ҭ3x}�?*�����B�~���[�y�l�PW+=ڧd
�>c��\G��u�[�y�o�l�= �<[$	iǰ�%n%��ֵ�" Ahm�J��رH9�$�R��6����o��x`�v-�mjf^��v��cmr���H��w)v��P�0�r�酷Ͼ(
�)h�n�^��1���Z�S��}���������_��l��{W<_��p�Fgҽ�]��&��T�5F�U��3�ʚ>�S�@�Js�k  	��\�4�<8�R�+�G̍���i���|D	!�(��-G�"�j�,p�������z�}���ΠE��������~lA�b{��F7ǥ��	�f�C�#�ϤK��vhe]�c=s~����WOn��lf�@W���L��9���=���W�;��bD��e!bzEi��\Y��.[��2�P����Q5v'§�ڭ��[�U�|t�b�mő�`������d~v����>���TY_���W���1\��,�8�Z�(2�;s���E�9l)ދE�ç������Io�3nw�&r�kY����i_���7�f�4������w�D/���C�������kcJM�M�C$�"K�'@�$1��a�B|�D������5����_�3_�7A�bM�Q�[T�~,�^u�n���.)����Q*�x:4Rk�&��T�p��
n�Rb�Y묂����5���ܢ�)�2�6�઒J-�S�sS�.� }���j�PW�`&A>Bsn)�׶(���k�9�b!��w��D��63uYgo�QD\Ӻ�y����|"�2H~����~�ڣ�	���uoC٣Hkر���n7S����-��J>��h�Z_D��<�6\`�&�3�F����273/Q/T�;P�-�/�S�(+I�=d��L��g,$W����q��;���
^��#�:����x	̽�r�B��Ը���9^d��f;����ӳ�\���:<G��_܋3��D�a����i' )��[��CF�|��[���Us!>�㍀z�����t���Ys�^�Х���ͮ�����-CY]r���T���`�#�xv��{���H��T|��6���g�$϶�GG�Y������s�s��l�Qe}J5��2e:%KcΖ�P�gy(|��F�s��u6}��P���E] f\��"�������ȊC=8�-��b�2a����E������`�7�`MM�
��5�JфI������s�� �j�n�׎����	�Jo�2#�sm�_m?�Uj>%�9K����G
�Z?��@Z�y?p���Zh��x���������(q©�$*6���_�gM̞�7���o����v~��Γe_!nF�d8~���(����p_��Xu4�>�~�7Z��	E�Y�.s:1��R���������8�S�0�o�l�{I�x_ڤZ����f�/AI�!�ȃB������Ҁ����ZF�<����]���E��f@ NEċ�K��7|	�xx1�#��7R�R�t��o��K�|��;���VSkǺ�riS�uB��1dl�S��3�Ő`x||�B���M�� �e4�`*�|���o��$K�w�odu�e,�(�ƌ����(`2��a$K�����䆊^�١
�|�%U�ش�{S��+�S��z�~�x��6C2�
�5���V�n�k7�u���ILLH�g��f�CV��`�t�"��@��Ew�ʮO��;�Y��}U�{;o2�m�+cE��`ד&"ޣW��n�:�k�c�-j�H�xMSY��.�Df��?5C��^Q�p �\�E����˝�S�8�4�0=�EG��ZH�xC�]s����[e�vP�dD:"�Sg��i)���'x��&~�I\�*�+Z�x��A�.4>Q7
��bv�;��m�-����lI�0R����Z��|�[����mbiDB#�E��qg���կ��e��qbN�+A����c{?�#]�Ӗ�+ջ�U��=ϙRh�~����{-����������	�|t�8U6{���T����]:J�ڑV�y�)�Ie����sV�*D
7�(C3`
D�����']=_��	$_� "��ǟ���S�F܁���c�6εm��J�d�A>�Tr{�̊��Xd�"mKv�?F�j�-�M�טȧy�I=ǥ���]}SA�ڱ�i̼j"o�m����Nl��a<�dP�v�����w���8^�?v�#"^�g���(����m�)�7��&XD���1�5���0�ue\>����vF�HL^����@�y(.X�9�t�0
2L�n����@t�}�\v����)�L��$�+t�;F&;��J�i R����y�HA�l�.4�Ȇ��/er�Cz��<��6�0I��W\f��'�S��S.rg����^)&�JF1M���,��
���+��Qf��9t4=F�����o2