��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P��v�"<ߞ��&'��k%P碶�R�ӣ�sĞ������FY&�E�����7+������s���.�{°A�?��}K��7���`I�OU9L\�T�E: ��^�r�q2�b*K���٭�@H�z-�1�*(�ۄ��si�A�B��ui2�-��_�šu�V#f>'e �7�p�rP�"�Tv((����4e-0>V��G�Ld��陂󋺟p٘�y�6xS�����C)p:�:��2��>Ww)>P;�gY���0dʦ0��|>��ׁ�r��td�CrRh�C�����]��aQ�3�� TFF�b�^����Y4�R��f��@����E�S�2�v�`�����#�>2�hm'F�Mp���nLG�o"�MV?��?s�9�=���=��N�#����XM��3��}�6 ���sS���aZ<��~
�l�Ⰸ75��P���z�L���m�1��L+��!�,+�ը�µ}�{�^�'���q�Kc�s���t��`��F�0�`y�Wz���э��L�yL��H _0͔�v��&l�ry^
Ԟ�V����cô=�1Ţ��['|��m�~f��GMSۭ�ت#�i�u{��Pm�����.�A��~�i�q]��]�×wdE˞|�֎w�ɽx�`�A�*��y�re�%�v/0�"I;�����.����<�l��d�7E�~vv����YD����sDV��U�I�B�_��	�VW�-�-��96�G��F�B��'�D,k�Jj#9��]'	�8���l������8�G/f�z�)9��i��u{{�ϟ7X�0�.C��!�,�<`�ܲG8~Yt�(x(����53��F(8���k�Wb�=3+�z ��<_o��1Uه����-!�		���=SE�& "U�ꇑ�WJ���lw�jm�Y*@,��N���Ȁ�/�E����S48?�z�[(D7�u�@HQ���1�.��f�
(l����PZ9 ]Z}k�1���B�>9��
�Qd��`�U����7w��)�|��Oǻ�&��K:}�x�]i��KW�1�0�_��s[�:�P���/���-Oue=kSp\�M������| M; ~��[�V�8�s�`u���U���dq�`Z%�E$=Y����!���A8X�~ ��!���/��?��*���0�b UH4�/�y�`QM���e���u|#���Co�Y����G��}��`*XOoTɿ%qL�9A,�~��c>i����O�Z��vM���WmB@� ����bd�Ѐqܑs)�.4Hb
���E���.�h�yx��>sDT�d�=w(�l$�@4����c���]��ێ�[DK�D>�M����9^D�xg�����k��}q�*����	[�����f�
<Ul�.�<�ƈ𼺋d��~��5! n��/�LK�Q$g�]�zj�/��3����N�6���C���qi�i�A̂�S��c�~�k��k���,��O3<�XRKA2��F#܏7��I W䡵�E������	k��ɞ��LGŞ���Ѵ�s����= a1���Π�4�#���:�37I��ƿ�W��	��~#߳0���z.?|���A� &���a�$�W/�Z/�sO���nN�5P�@*�n�����WU�j��xq����k�n����Z�JDw����Y�1�����P��)����A1r�NU��r�dBpN����"����,IQ���;k�)�� �9E�*�a���+���J�][)�j���:x^¨d�M�EJPWH#�p[�\��(,lHK�=ߦ�S���|1L��(��NY���z�.g�D�k��]��3��# ɇ�B��e��;`�vN�9�j�ϥ�r<�n�%��V��N��R�v*EB��ǻ�f �It>�_�����d�D/��I��r�h�|��WE���L}uT�g��r�t��a��^~�ǂ����\��8T	�Z�p������h7Q���X��	6qyh쌄�+Tl�ƶw�$�} ��u���f�c���������u�1�^��[�V=cv1�%���ߴ��F]������h�\X�Ś�mdy��)�{�3�bw����,�Q�#z^/b����1nč����~� ,i��3��5�nX�ҵ�4�t��O�`S\o"'�H�l���+�Rn�D�5����� ��f����b���\��ac�.����^O;%}Լ�,�89�uH��ş�m$���Q��aY��:`�0R7����4X��� G+����;���i
T�S����fFN2��\��]�1؈촌y#�~����+F��i��(��|\Ζ����.]F�bH-9v�~SB�D�X���e6ڶ��KO�y>�{
�L�#��)�ݣ9�"IFx���蝚en��wY�Ǳ �k�����Fuxs� &=�X����#㉦�9�(��/����H{��`���N8WH�%(�IN��g����F�lSg������1����tι�%*�S�QD��Gv &��Z-��r�2xz��j�"�L
3����X�t��Z`�I�͛�2�jH�G�C�D� ��T�K9.�ڂҼEg�Ȟ����_�4�j&�Jr�*6�z�-���)f#:�#�<BY��ﱯ�Y��~���x�dL�H<�r���G��5t`�d���}4�>�";�#�ۻ��,�*�h��2)jø3g�x�l�������Q:qG�&j�A�t_bC�S?>ihd,D���$]T�e-M]��+Xr���ղ;����D�����Q'�6��ǐe�0
��RmaGJC�Ý��Z��F\��'��W��
��<��%���+���-N1H��� ����?���0�C?��q�g�JHJZ����~�G%�7�6���@n1?a����x��;)277;�kaT*
�Z^�[*�}RTH}bՅ^q�+T��u->���2ĺ���{���X�Y�G�u5����畈�T�6g��`��
	�(׳��᠉�N�L��4��%�|0��5��;�k��!��)�质��&j���k���7�x:|oD����/��x"������~�f�q¥h�K5Ϭn���.�Nynp�͊���f�D�ߘ�[�ۮ��'�wWؔ������cyub�M�'���7� ��E �{�ↈ;��v�H��r]�_�����a�T�G�o��y��G�ْ�]���7̨��o
_�7p��(���&�e�ȁ��,���ٴ�;����K��!ؒ���v=2T���y$�6+�*���~��Q���pa�X�u�4�Q�.GQH&�_��j�v�ە�|�eX�g���<�����ձj�17xk[d&F��IЋ0��oܤ����A�qk,?�vTF���5K��~�E�ei*T-3|J:��bzj�綂��?�L'�(.<�T\�c�Xs[s���^��>�9��Q�n�X����#�w��ö�z����$�rz���m���i8'9�u�7{ t�p�EC��u[5^CT�� ��k�z*,�BBv�L��j��/t ��]O��@�`|��U��8��a��S�eJ`Zsٮ��-}�{`�S
L��g�F��B�9��J���H�7��$����p|nI�n�FΡyl�dӦ7"�Ax%{��d�[BSꙂ�gƣ{�}�b{W�I����ӷM_j�h��Y�g�^RiA<��k�@j� �b�T�����\�wY6O��X_&ݮh���VY{��u����[���)a��uY� ��6��sx Tl�
"bp���̹�p��S`�ÿ^�2W���w��8��{r�Y����_u/���,��y���do��{�
n�D��cdm��c<�Uv���ƈL����ٌ��_x7�ȩ�\���� c��,�,���j�zr4�<	���1	h8s�z�)#���r��� �:���?Jѓ.w[���r���s�  �D���K�a;��F���Y<�*����L��2R����6�	�ʯ�pM�g��q�.�N�=���B����rn���h�mL�k�@���Uƶ�eF�߱��@ABҞ%Ɖ|�l�Uw<��8�9>�<�F�@���c�
Ig�VF�*$��<	�?�1�"?��N.c3�� �#[j����k��ݜ�J�B=<w�E,����'V��CB��
3�^Sh������*w����zj�@ �,��v3R����0}�,a͉�O���O(ΰ�D^��U���I�	���cH�R�CFU!rҨI�⩻=�vԪ����{8�7R��÷�ak=�֊Xs�a���j5�M�Ȋ�O�ke[�{D�v�0W��t�E��9�y����$J��p.�*���V7����n�C�@6,�
��7�z�.$�~�f�6道����U���Bx4��Wf��4�!�C.h��cX�b��n�?�U����D��\��踑d����|\��OtUL��x`c�ϬgM���rCm~�8s�_�n�y+p�dӂV�y����'w���E
�{p� M�0D�/�G�.�"mBy??*�'�3��/���i*�E�� ���Ŀ@���(+�L�C�:؁U�C^�<�H�X� �+�O�٧ ��)r_5�Z{���<�Y�l�?`�<���Yd�3���_����F�@+Qpp@h�`��E.`Q��:�u�<��%��^ Zp�6оѲ۠h��5[�@ߺ�j�{�c�e�>�hx���r�$V&`|)���\Hd�"�ge�n��^z#s��lШ����/.[����**�H(�J2	��f��;��J��z�&�Q�� {�[%�j��ǃB��4�UxofX�ӑC�r��(�-�uh
�+�U��t��|u����KU��rIE��ѿ�>_p�4�T�����f�b��HS�ƙ-�yf����HyR����!Ex��j ѯ*��Ax�b)|�k��3���{fEM��:w&}. 9�c?M��.,�� �'����o�]������-זO���չ�ɱ�r����������N���bH6��#V򀅩����^q������K:7dA�tq0+�P�Ӻ�}�O����
�]�.�l#%������Ķʎ1b]�<�c:�&yrM <ΌK �"o��S�?�;�3�|
���_�L#s3-���0�)�@��M�&&�/��t�=���M�3����{9Ck�Y��m���ia���X����k���?-�ϱqi!�q"��虘��jg���p#t�H�U��?�[)��"B�PK�p���|H?�M�����t@Yp"�m}#>Z�����U`��uZoJ��I�E���p>$U�?jia����	�8���'�Q���I[`����u?�b�kHrE��;~\W�<��m���}o��}E.�������2�{��\33���<�8c��[{�%���V��c-�ˤ�!��V��U���@T�$�k��x��=rs��\�y$�Qc�*�Lف�B�����Z'D�&��vo���V��H�(jVRz�ƺ;֘{�U�eh��δs�Tu2����~:�B�����9P����1`Y�#�ی�Q�|I������bno*|��h�XC�>f�c�$�%���˜]G�N�08�[Z���O�]�҄8��G�rf����p'TC���{(f������cTE���ԙ�����*&TwL7�z��K@� yf��L�U�T��Q��/�s��}>��Qe�5V~�����*uM�Qo�o�A��7�j��ڣ�� 9ʹI��E����V��-����B��}]w8H�����ψ�q����X{�΍sk�&g�_�c^ u�Op�
 �nM8���:}K�xG6XAX�^ 
X�%鶐:8�9L��q� 3ݥGσ�!�|V�ʩ�C�Q�#2[�����dm��툙�Kc��/�!1� ۧa�_5*��_�1�T��+�Յl;�`c`b�z��6�4��E%W�vc� ��7�ǣ�ag�/B��%�!��hz/�ʂ�k��`��*N���[]��n�VJ˹��mX.�ݕ-,���{���W�?��
��s;��#K_��t����}n�ƳT��9��s'�:��=�x}oK�G��O0�?�9��u�<�[h��Ll!#���|��ӱ��q��EP�H�4Uy9����z��?��`: �Tm׶�Y�������f��#"�v��K�}�æd#z#9��"D̑J���z�K8q��\R�dV"D]�������P�BVM�W�|I�6f�Zt�@�F1�˗�TԒ��ލ~N��4L������@9�E�ܤ9LpE�����q#H���O�s��S�~�X[����5PU4bJ�.t{������ աM��ea11��͡N����fދ��ZuQ���X�e���1�#A�$=䈐�G���'.��K�`G���v�b��k��ލe��ϼ�
T���ρ�)���=���W�eo=�x�c�R��#��|^hH�߆�ǌIc��E���.�h�X��C �����~`^���|��� 
�T��X��R-y� 2�ഫ�:��k��y��w��L�ܴ̒r������	�`���y�Ƨ��m����0U��n����-ˤ�&���5��Y	�;(�'��>B(���/���w��1ɬ}�a\-�G������gbiQ�x�;R��K�:�����Y�V_d�
fFY6��z��vu".�ٗ~:��/�S�#�G)���h�-w%��邖�`�Ry��-��S%I;f���q�<��BΙ�)�/�dt�T���8�U���y��T��L��.����C�$��wQfk���9�i��[~	��0����y�h�/Y�QY?k���Z���i]6K~�����J �k�%e�y|3��h�B`${ @v�+�'�����IY�h�X��D4k��i>���Ԛ
�-�.#(��БK�(�T=�t3 �1_ ��B���CF���L�Ŵ���݁7'[vMX���.�G�)����>�:E�f��`Af�2��?���>!jp��GÆ�Y��M">�@�Y޲�H߅����#�:���8e�f�r��w4G&��|.��On�o̫?�L�q�|k��%�.��;Mm��c���=p,�~=�4Cq{�=�	��u<��JH�l}D�e�8�Ϣ�H�yh(ޛ��y5R�ۄ�r \�~��$-n|K�l��B{@=O���<	Վ]'��F_+pı&_&�l��I��5M�C|��c�ǐ�U��Q���\�����ߘ��჆቏l�b6h!e�ޗ_�$��L=-]GͨXa�WlL�����h�PʚQc	����/N�<e��\��=h? Ūſ��w����|p3�IF@p�a@t��E���ج�f�l���|1�^�b3 4��uΕ��W.�6v�׹n�9�����
�<l��M?�T{[�d�2�YЀ��;�"�-�C4��6:o�"lwУS�CUR�·C6-y��̱���H!:�Q���A���٤ �@mqC~)��@A��W~��{[��v����e��6�E��m9�t�4B���P�증š��W\9/��
>�����Cu�QQ�+Y�7��1b�����0,�$]�nXc�2����/��K�J��L/h-6���u�
T4��䧠�BTb(ۼ
��*�Wu�X�$���A���&a=K�F=f�8}L��'�������� 6�m�_��1i��.-C�v���T,�s����c�4�uO�zܹ,4���t�U�y^�G���K��߻yU*+"C�֍E�z�*4�1���a�R�H��OqIvp+���#��p�sםuiv��XI��U�4����V��`��$U�1��0#�$s"�|J���~���|��0iC$"b;��	��lso#:<�0� �9g$3��T����l��Y�UH ���'��a�fة�n
�����Kݑ�|?������(�ᵟUb�H�7~;]-B��8�YKL��>]�m~��Vu���\��q�f"kF=���� ��c��G��µ6�OCB�Z��C^$)�+�VQ�t�~�l�θ�p��i��3����$�R��t�|��5�!@t���K�p��k��C3?�W�_ z&��vM�$H4�oF8�#k�������Fa��b��3�o�?��Z�V>�:i��u���g�W�K{¨jkL�9T��m|*?-i�f�dܮ��L�tH�ǈS<��u���<�ّE���?h~Ժz�y����b�x@0��.��3	��@�6�6��f����Ad}NR �:��!fy��$��G��T�&���7wW#��;S�X/�p�y� �>쑥��P���x2��ӎ���ܧ\.��YB5ێ�t�h��D����>b,���M嘪�;�W�e��E.��$��X�9e�*��a,s��`H���Q���wBC�o�N*�C=sp��5�*�����*q�+0ߠ�:uc,&K	��f���Y-WO���md��c�ΊHF��9'�Y��&܎��Q��|�	B^z��*�|�䵗��T�Kr �'3@c�U?`��pa��M.�LX���T5�x��$�@����ZZ�D�6���i����rD3�THY �C��FTQ��7fOe\���f�r��5���G�&p�9��������s��r�eј�����o�_��;@]!C_�Ϡs_���#�\/^ʹ�]i��f�w�=�M�L�"��N?�T��;��16q����h(o����M_8ܐ5�i����2,�A~Ͱ�	��N<ݭ�KR�|\����3�P���z��àx�{�ɷ�4��d��۷/�X���VK�/�0%Y����_�Ŗ0���8��Kڡ�y �/N�/�����h�!?���x��L�D��� ����--�~�:�v<�����H�����G�2����y���_S�+����:�h�T=��?����� �5�����$u�x�J�A%��3O����CH����oHd���Ө�A��Hi�m��Ƞy6Q�t`L^���iU^��   ��ӵ�I�&Mo`�J'^h�����Ek��M�ֵcT��h�1�9C�=S������Ud"\.0�im.�L���xD4��+rĥ@�[��b��k��Y�,�*q��枲�Fe_g`,"�]I=����N�a�S8���Ib�?�����t
�τ�\K���y�%ݿ{n�> ]"��g��!s�N����{^ʭ��N�CX�z=\��fa�'oG���ӳ�J5��u����e9���H�M��CuɃ���0Y��iT��`���\�>��b&���{.o��^e	�A�T/����µw�)�ڂ�v�ϔJ5_�_~�<?Yr�C�C�½?U��c�t���þ ��!}��)7��Ș"�l([��';�q���B�EV�#z�Q��uQ�o�0���R#���V�}xuFdxM)����\h��jQ2�*�B�t�;�tɛ�#���5�T�P�X:�/�5u%���A�{�M��~���/���9OaƮ�Qk �����Ƹ��9���:�(�CL)�HI�I�-�d5c/�K�lXU��飵1I
�����"�3a��D�"?tз�G�#�V��)A�S�nɰ�m��,=N:�DM��A#��n�3͂��ń�['`�Hr���AB���io�pa�}(�r&1~�«4���:걝�����R�io�����sE_-�e>tRʲ%���jSu!-@zb���ݐz��~a7�A�0�כ߰]�A�C�����~˧I�ѡ�a�g_B�I����f��-g�|�n�A��k�b�E	|��P��<�B?9��:V��,�����d�9���'� �-�RG:���߻�TQ�B��_�i����փ>x��"�5���ה/�݃�'C.۴}Mo��9�/�����>�ꛖ˨�t�f%�j�ю~�w�f2/gS��!��nx?��TD��p1��(�"��UHT�Vɺ?1�!�3��Hn��X�=�l�hF*���9M:����}�&�4�ZY�:��;�_5F�Di˶�t�>7��U �c������I�!�;k��!B��'�LbG$�+�)�B\�i{&g�;�i����������=>�BC?�Z{����#�x�Ձ�&���}i|q��kS�l/���v�� �<9֗���/��|���q�Ԝ}�F��^�@"�H�t�a��h=-��f���fP�i4|�Z���Mp�7�j��M�!Ѿ