��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P��v�"<ߞ��&'��k%P碶�R�ӣ�sĞ������FY&�q����H6�:���M���$��5
�J�C-����no��AjQdd����:�`w�@���Ey�r}�d�����݀t��&N��z�l���Im~��!��)�ݢP�̥<���@���#���R'��^l�YQ���=L@����':�K�+< �����
�I���EǣEg�x�&�w�2������Yj�+%?E�AT��{�h�t�z�vA�^�����SZ޻i����HZ34^�Is7Vr�ѹiLث�.4�3��H�{	Ih����o�5�*��y߿]��LA�M=E�Q3Z8�R�ja�h� a��~F�F�ѡNph>��\�烏�5�-�e����ϥ�0�s�
+���L�ӦZa��VT�!$.I8%�������8I�����ĝL��q,�I�	 ���vq��A��U��&t�&TAZZ���j��!Ψ���?Gܥ�C�Q{�U��
�q�W��`K�&b���"��2�-̋�ay����3�7T�tq������ѩ�	~��p4<-\8"V�ԙ��r��hU�� 5����
fE�W�l}:�
g��gT>s��*$*B������M-^�*d'.	ړD�)/��q�D��uh���k;Y�Ed���'d��u�8�9�-�/юNo��r7B(%��[X��k@�f�-zq^t�~��u����)��23W@;��M��	�:8/��Wթ��dFR?�yf����bo��WV|lP��D�d�}�X3ׂ�ݠ�$ I����
��ٟX�<��.��GK�ˣ����/�3j�G���*o�mxk[��"5��6p�[V�� ŏ��e��w!@`[�tfAÕIW��km��jN�R2����w�o����'9�hMO P�Dtl�Ær�F�0�Y�*[��z	��Ɔ�[�8Y����^��:>`��ޡ�L8&�LH�[4�Jt	)��d󽻫M��0�-�%�����^:�eK��;O��b�e�Ϣ�ЖQ���K�>&O�C�)��:�'6�Gx���c7�׹Γ�A8�#��~�r�楘5g�*�a�*a���޻x�&��}1>R�]4����lȔ�=��_|qL���x)"�6���m����)^LoDu[�����f?�`�j;!P�S_��C�x�0�#O�Q�y�4UJ��_�2<�Mn�q�]d v���%Z���j�}�#2�ck����n��3���}^��+W���;�	`�*$-��m1�w��-@�	.����zA��O��5��U��"�ZJES��%�8�n�{���M93IE��ڎ��pؚW��H����3�j�"�x��c����a�s���'��P��d5V��bL?�g�uI�
���*z�

�n!.��Ȅ{���z��Edb)S7�����6
m�aK#��7��tQ�� LB��PB
�$��a��e�e��2<h���k��A�	�A44O=��8%z��3Uzw�q������J��2-���`0b!�,y*�0��w<���i5)jEƂFu�}$Ǚ�C8���7������������"����g[�4�����
xeQ�ѝ�B���E��a�/�����{ �4~]n珯W�v[�T��_���|�ht��Ș�t=�ᮓ�hp+o1��6��2K���hC�0�*k��%��xyp�B��1�⾷s��. �|�Š^ڒ��3*���P�[�1]��7��.�U`��O����2kǕ����O�q<�[h&G1��Я5���Eh�S[�8RԦ��:���.�
C�9��g��PbT&1��^)~9��n������Xgv��Ņ���q�
&�+�7R
z�Xa<�"K:�$�w�U�ݝ��2�5ݒ���K��-����J$��)�DP���5���	t�^��t�w������Aև��Aڪ)���᭟ �@���=1���������@%�t`a+��y�x��r�FL��g�Ah�r�������#g�][��r�`����+=IZ��vX{a��{�Q~}���Xc��!�Hҡ������J������b����6u�K=�G���VO�L_
=��U}�[W��F��$�� �=����۲�ޠP������S2�2�i��z��8�������H�oQ5�!b�s�t�d��f�(������`5�5��D���,���*$8Dߎ�Xs1b.�`� �0�J!x�RA1Hש1��ѥ�g�	jE�x{B�����n^��G��%*�ݱT�\.@�(�K�9*����Jbͅ�Ϸ����q]��U��ª���B1�ڔ�oX���[]�������U�<�����ڭ�V���E�ڸ�����7�{3��B�<�6(�m9;ݘ`��^��{��&d �����rR8���F�bY�C\�?�j�t:(RY�7D\����������f�\ԇ�1�aw=q�_�6�3�mx�fYڄ� �#ޣ�]e�U���1U�_���D�F��<�f��B)MX�L�x��/�9w���	��F�P�$x��u����ak��Ǉ�ÝNn�UN�m��Ij�۪�"�G�˟��u@�`l5`dW���,GON0��ΪX^��7�Q���K�����d��]�V��b�!�s8� ��V��m�d�Q��IYY�_�W��'g����[���:���������%tN��A�$Ʒꫧj��p�%���܊�7r��;w��2H��l�el���J��E9vP�u�L����r:�0��R��VzT���V6�,�(�T�=;<}N��3�/�v��s.��Ζ�:Ĵ&l��Q��q�N���L���Á�P���H���RU�_FQ5�R���� Z���<"�YK7�O�a�V����jM�ŵB#�����?�±�����Ct"{'�7,|���� �?����*��_�x�k��d�4S�؉�\���n�]᳘f�.O��"����5�:����i�.��q��:��N� �#�w�a�g	����>���ْ�g4Z� .O�G���2�k���qu�7@��������(����O��J�4"G�1�~tr��7�����\����� �A���r��T1m���M�w�u'����
����d�W�:G����S�5=r0��l����56`S��8�.l^��ę�.'0���8��5A,�Хk#jn=��Z�,��ð,��H�J?Z���C{<�Z��������i������7�V,VZ���~�|1��1�+pѓ��w�M��jD���@O�Z�V}�A��({���8"""��q!
�&a����Cz�7���xI��ù�9��k5.�V���WO�t�-��TYc8EG���+�[��l�'�zO�ܬU��;�( �ž��?��E9!���e4��UT��+`�kHr��n�bN��͖v�[C�����˹���GĘ�����Pf=�3+{.��M�m������:/k�/��w(��X�|�Cc-� s"_D^F3Ι��u�!����w�c���^�תG���G��� 0����đ<�X��e��[� :X�1��tw>�:�oc�:(8I
�dB��>)ULP,��s�e��{>D.��)_�xW2ĭ�4K3Cu���#h#2d��]�ʃ�ʦ���L��1 ��3Qq������D�C��.�^ ���&u���?�t,�U7�~�D���Y�����K�OQ�8�X��3~YV�r΁y�GƄ�U�,q��Z����-��	d�;�-�H��\�Dol^��ڐ��"��/w�}��~d�".A˸��N�~:��7���oԍv"~[d�Õ<i����H{�qv�[�k<����3|�#O�{���:�Q���[��z�c���;�~��$>*�Z>m�F�4n'��a���9�+a����"��:g�g]&��-w��h�|H����=SO��mm]-�Д�� WK�ᒺ�:�:�:�Py;x|c��b3�Gd��;Gp����Vc�G �B��L�r�*,8c/pIO}�;����[�d�FD���M`�?|���i��� `�2�Cq2B���t�HL]����HXU�?�b���d"i��8�١Ә���֙��=�!r����
[;B�:j� �kmy��1��*5�z�?G�E�f�8ϖ���A�Ӈ��Z˕�k�,����^���`���}@@�_�L)��ڇ8#���OkT����=*)rz��b:Yۘ'
tH�]&;=�[D���< ��4X��VHW9K�E,b�ٝ�o]g��vEw�� Y�Y1i���-��
�Q��<���<0,2�ܼs�IN=�$��q�xR�Q��!�Ѓ�:?���/���mu�	�eɁ"���к:�'�mC$�H�j^�ܧ�p��㟿��[�\��2{�k�nέ&�1�j�"J�-��I��*��NEI��pÐ�B-/�y�5��g�H-7��n��X(ty�j��gY�U4	����]��L����@X�����F���9<n����;�F���;	}[���Rqf�\�w&��W�ҷ�1�:�ׂ� w��6����ԗ5��,@Si�����j�hi���;R��,�u���X���QZ㆞�fn�#'��Qz"�I�4T���X�z�l{>��o]a0�M��6j>�T�eq�1���_5���W�猧��b��tq������
�D�y39�^� [ZB���A4�A�0��	�R�iY�7���Gz����,��}�� ^�Y��,T;��@�&ID�����,P�F��w0 |��z?���s?����Q����4�Ќ�9�⊺uf��/����wi�>�����S���f�����]�zA�h��qj-��h�?v�����>Y!��3~f��Z��5�0g�#O�c��c�����N����B�vLi�����@��g�tB��ZC�1:4M61d��KPk_875Y_�l(�Թ�vm�a�J��x��:�O�G�M~z�(X���3�\]4��iǙ�Q��%/s�P��;5I�{����u&��eN������E�6��eV#�U_�N��h� ��h�R;R����U8�~/�Ac�#���!�˺�;'��O��~�0鮷�Ҙ擱�ͫA�