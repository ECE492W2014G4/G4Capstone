��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>,M�Kߤ�V�P����W^�o��K
͵h�����h�
�;� X����x�Ep�*���'�p˂#gD�4H��fZ��"4��V��6��cq�`�7խ�:����%�	��H��\	516�K�W��K��ֱ��q3/I��	�0�j����X]Pa$3��	���l�W���Й�̸`R�d5�^�m��	��7���_�7��c��GT����T�6v'��d
g�Y=׎�IO�p����[m����.>4*�:kCR����	s\/ux��<���rP�!��c�;E0�*\�����瓻�_I&$`�vG���\] �T:�����Kj����7�e�HY�;�EL�+޷m��;c��i�Y��#S@�h�˕������6�Y��u��1��a����Z]�T�`b�ǽihA���r�(0<N*���w��Ϯ�s� �i��� �<�X�V�F� �CCK���2�:��ςO�޽��{�['N�@����*sV���s>G|q���
q�2����G�%��MY��ԇ�8�s&�m(�U�(}D)����n���Y��-z)p��6�=��x{1i1zw�4l]�A&���gE�������Fl>a}�	�}Ix�h�M�J ���!�/k�B��v���ՠ����e���=@�E�HM�����k��3*/�N{d'L���Y"�dnT��SؘIHl�O�h�b�I���.D�Ԛ�s�~��M��r�������w;����̆�`[�Nw\�R��ګN��f��%�h�ۄ�q�~�p�]���w�H��r;~�=b�
ǡ��Jv{Ԫ6%�'��*�</O�u+E����'�����8��"��h�����8B��[f�W�e0��4��f�)5�+iP���:֚EjN��6�-�놹́����9���I�(�5΅���8����U<���t��r�h涧���!,�`��U���|*�V�V\+5n����9��!�rƌ]�Ee��M�Inھp�(\�r]����v�yQ�=N��h���>a�@~��DVd{�}'#
g6�>�*�AY/I|��9��;ƅIt~��2g��� ���s�D�uq2�z�p�UG���Z����9WN��Z���?)�6��\���Z>�^ݺ<o>��-N�Km�csɷ�&�"�NJj1��g[ecn�|��H�j��C{�SQM��7�Tɏ��5_%#�^ P	Z*�z=7ڻ,�;����%�	v#9�u�=��"ӝ5����5Q��KNaS�(�0�2F	`��;�uNV����y��U�q��ـZ�(yi�-����>����78�s:�5W�<���EE��$�Z���YY/IP�� �B������@'K��
t�-�,������d�`׫����nM�W���Ͱs�����3���~��'��{q l{������OX�菽�qj��Ϣ���xA aLD'��0�V*�8�r1�Occ�گ�Ig--���d'�m��^��}t�>fK]����D���sOwaz�i�9�B.�>P��*���\vB�=(
]s-���j}�ob.�e/]DԽ���L����,��ثL:��M1e��l���ʋ��C	�Z��D��Z@���z�*9�Lz4K2l�H���L~EC^7;���%E��H�R��z�:��*1D�j
��L)-u�K�{�E赅�:���Fv�|�X5/�2	E4��	�/�羹��m��4��	2�����/;�)��^��ѿ>��/=�iPW�1Cj(�|e�(�߉���K'�̎eSKw��
ܹ�k�g�v���Ϸ�8�9��f�5#}�V�:Z��zb�wb��!�x��'|�fL�������yA��h�����E�pD�����@���9�0��u�"���li<��P�1F)�� Y�Z�oA���NWnF������o�ZI��\���@?v��8u�WڧC�b��Cl���
�'�J"O���=�G�r�ĥ��;F�։J�Ye�v�����3X)��3i"C��3Lm0VbY���B����"g����Ő��o�ff%�E{�xД0(��c��i>�]���2�Ɇ���"<;���E=��*uh�������!��`�b&����T�I�3Teϛ�b?i�{g���� ����՟)�9"�Ւ��sM�'�L��^��z����:>k~0�b
V�i��ǛM
�i54`��E\�ã�<	�^������#u	B�B��=m�MS����C��ڞ�n���Lq�ܝ���]�����D�6g�ESC���"�����%�5��2������ʕa7 �����~�)��5���$����R;��ֽL�3	B�ʱ#O/�WF:��������?3��v ̡����tf��ݩ�?�S��n��}���Bt�%��͌�[���F�M�
'��-쾅��;�O@z)��� �S��~P����=&Y��$.k�a®ph���g9��pYE�DN���|�]�X6��4���۽�ߧ�=��H�r�N��\��h= 街*��/]CU��c�}�U����Ðd����R�۰Նs�`8Ҩk
ZJ�B��*W�L�����Ԑ�WH{ 3�@�w3�wr�ݪ�	�96ҕ��w�=����Xy�_�
�/|02�{?&�߃��Xz?��)u.���2�q���I6��u��F���!��k>&�d@�����Vh�Gno��f'�Z��v?��-�b�l���ɛ(Z�)�I����i��b|.R㠸M��ȱ��b	���Q�k�\Ғl��o��CLto=q]EHֵD��M9�m�H ��ր��6�	�ia&"�*.�l�d��eq��@jE��i�b���T_t����R�?r)g���@9Z���E�QV�U=�lЦ���&��+��"UpuJ��(�^V8W��M2Ic; 9/Q͇��.�խJ^�˒(uh��KtӘ�����
�%>��+N	��
�>K�	k�y�$O�"W��� T��)��"�k��C�W� ��Z7@ُx~��q��Ԙ�4#���G�|��ӕɐ��%��A���/�'s4\���%D�-�[�v���I��3������#��b΄u.�B�UjC$^D���jxnT�,����S���FVd%<S���v&%�^��h冘�ޞ�_o�/x;`�D� �8&׋��T�u��c�fbi������<��Fy��a�=r++�5Ar	������)����wu��d�6�g�;-���FZj���[�$�*AX��b���&lU꿝�짖-��wMv�#f�mD(��G|�^Y�ց�&n4ba u6��1�������"�d�ng.J����6�1���T���jq��9�?�eiN!1���� t��d�6?��$�ц~F���c�N��5o��h�vvFdA�(=��k�CpNP9x�:,�l�Ll�d��h��<���#1�v���B=eי93} �
�R�Mo4��c�,��7B6��^�|��J�DS�'�%oo TY����E���˕L��J��Z�Hy��YD?��H���XIp��&%�3;R-s�� J-��aTA��%�W1+�2y�����c81�ݭ��	�@��qY�D�`���f�������r�jg�S)a��jfY$s�T)�"E+5ϸ�!q'q�k�h�QwFd�M܂�/o4���sP�i6����u�|Q&�b��يM9��|����@3{6Xx��Vt/u|���VZ�"(�AĘ,hZ��[MI�i��̈q�q����]0�`�h���&*\>Vr%b�����.���Z+���p���9���.* j���R�"Z�p\NCc˲��d����د{#S��݀�$w���,��NWE�ʘ3�K�F<:5f�9}���t�
��z�mT�� ���)|4=�=icT���Ȣ��X`ݍי�h>#Q�}"�J��fk������U����&�W�<��blNT����"U��U��a)�a�"��O,@�.l�:�������i��k�yo�A�R�&�Zw�ysF�RP��c����%` ��H�N�?+il���n�0?��$�` ��5\(a���}x�y���[�ݭ�K�?+Pȱ���E���n>b�:2�lᠬ��!�����T~�!���1�&�dX)�,b���_�.tq7�@���S7���6�K���6�f~���25@�u�_/�C/�g��սzŤ�L=�dV�͗�R��zo:��'<3?u�D6�1��ʽx��`'p%������h.a>�-���{o8��F�kӫyG&��|[w]��K��Q����sl�d����Kb*���69�L5�zY��nF�h����se
=Qh ��I.���e{͕:@v�F���G"�P�0�?cKG~`ǺHI�x�9�*%yf�T��Hg-�A�Ś�'Ǿ(������<?�<%|���>�6ވP���Of�b}a=�	،���VNW����LR����O�@EVE�������_���~��z��MȠ�]
ye�>:V�:	�>�bVẕg��11㝐p {����w"�f�37��by�v����2�HɃ _��;A���`��s��&~E�Y��	$s��(�O��E���V���6���q��:��J�l����3�ZY���!*j���U�tu����a4_"�W�?�M����o�6�_��J�.@Y������5)}S�e�Oj�ڒ ����h̨���h~���%qjS��bi�1Ywo��e��s���Y��X������O���ђ	l��TW���4�?Pu�zlǹ5���CB`�&�8x?�D�!�Sр�;2��|�2nѯq��@�T��ճZ����E��QM�O�	+�ɟYSb��Z��y4�� XUP=O�{��|����PSp�����xXH؊�Ǡ�=�D�(d�	�{���?˞^Rͱ�*�l��'�����;��1yP�A	�ñ����]��6(�C� �7V|�WͲu\�\Q�k��r���cO�����/�I!ֽ�6Ɓ�t� �t�Q��8IZyT�t^9x�F�rk�[��TOY��,�"����v'���a��%�D� X�:�?�O~a�O�bqV�5��c�pܭ�*��õ��7�}e��*B���
�VaY�g�%>BT�t����ǈh�����#-i0��hpe=��E@��	%��1�=Ъ�f��z�8|i�$,��l��y"�u���qJ�W��-I����y��9_3>������`O���8�/����=Yv��O���Pk�$�i�^'�	
c���n#�vo�=�W?��� >�8���v����T�iӒ:g�������-�oD_����pV{����ݜ�)%��(�]P�R=�v��REj��%ټ���Ax.�ic��V�fi��3���$U��[��l�)#\U5�y�
���t*��l�0��*`V���Au�8�ڮ��P�����p�]X$W��ʗ,��٫�|���x�L�j��l��1w���#��ž$���\��_[�c���W�Ғ�]��_��j�&���aƿ�hĈǰ�;:jy����n�'���BXV�I��J�s�(�k�|ô�ո���c��`�ݶ�	5$�SQ���m�|��@nޔ��P���Y�$Qm;�=)[2U����'�����44�[Q�^� ���I�#�D_��=�Y��	'���	[�V}�?ƆL�B�D�|w���������1((v�`'E��Ec	��P�ZҋE!T6�f\��l�V�n&&�f��&�}	:�$h7:��KH�i�t�S�]8�x����?��p�{u�w~��x{/~����;��Ĵ�˼�	jSu���#�Y��$���T(?��y�𣯦Ö�/�Ob-�WFP�C��I��7?K�y<*ve�\��罥�*/�E�<���TW��z��ũ!�����S9ih�{�h[��A�P#��x�g�r>��
��f`R0w�"r�cm�-	b�q}���.B��r"X]��hz��,��NE!x�\%�t��
�����9��E�(�l��;�V=6j�� �^~�]�'r~�u^�ǟ�s&i�<�[��T��5��[�������Hz�����=I���,_<F������pww������9~(��������ԍ!ꚕ�B�������1V�ʦ�3�!3�:;�U�[��J�gIo�eKí4�����a6�יo�$k[R���O��r���)QyQ|��= ,�4��jE�܊�^����`�	5�\���H���Og� �~��fh�g�7�'Fl�U�Hwi�1u���m�����bpf_�)�6��$���[�_)��Ό¹��+��^+*���[����^�A�Vy��'O���e�X��ߞ��g����u�y�S���bg���wТ �3R��d=�P`��` �Rq-
�./}Rj���ѿ`�k�� }�� R^�6��&�k������+<5��6���
g���m�Y��Y�u~=/ݓ����Y�|o"\���G@�?��J?��=���y걀��+]��4C�4CX�g
j������AF� �!
��Q��w�C��g��]BW�࿡a����P�LU"U�D��M��F!�XT��H9X�m���Gj��,?fsTRD��
x�XO�7Y�Q��ei=��V����c|�˹<�!q��-Ӡz��uڽ+̅t����".׎)���I�c�d+���O���-��x3�ɫ�b�����y�H���S)���鈰�]�O��9���o��4� TR�`����6�XŔ�rr�t�ٿ22m�^А�w��c���l���*�7���U]�^�����yhl��0��>�E��J̞2��U�����< mg��U� /�!�eԜ�ĝW��4��:��l{���gY{�����g�7�%�G'�R�F.���%����|��ɧV��?Ġ0+}��x�G���t��ͭ�
/����Z���<� 6P�Ö5Ji�]�Z�u�Rı�bB�z�JH<^A5w|�r�:��F4|�ک�4���uf{�8����rl�kW)/�*�K��͐��ʁ�x|�¾��Eü���3B�a�x��� ��q�`1�s�O��y�,[Ax�m[78s�֤�ю�yM+��B��N5:m�W0�'��c���UEm�-��Z�����x��sJ���c-W/Y���.�r�a���p�r����J����$a}��O*���aI�.��� \	ϳ�Sݹ�x���SJ���*��v���e�;
�z��PU��	�Q�j��i�9�ap:ɷ��}��
�Y�k��)w�{?=�m5�z�GH�d�Ly���b���V�Pi���I�Y'��	�Og5�r����v�����3�t`Y괯�B1�I�#iG�_����ߚBO������2��92������]u�kh=�W��ߓ�_?������ӗ�Y֋a��O�(�7���	\b�S�D�r;��>�,�������0xaud��+-_���0��4�J�F��7,�G!�c�ل�����"�Z��u�~�c� )�e�n3]���;=%q�ӄ����� *�T�W�/>�.�����C�ܘ{���g�1���
��S/��@�U�u{�w���<��w�ڳB^��T�(�u���ZJ�����ж�?H����pti�}9��g�B"���MfF�@,	n���C6�)��0_H��Iv�byk��x���v���&����{!Z���COU�m4����3繌����s�+ꌿ?�\�@r��d=�	����ڊ5��,k���R"��x�b)��3~�J|O���#'�9!��j�	��Z|S�Ul��/e�^z���׸b���-���$�h~�k]MF˱_���o���mUP�� ���p>�.s�e����S�.Hº7�|d�f?������<��8�4��{Ċc��Ǚ�����8���ǄC��&Dɮ�����B@<��1����<6�<7b=�`\WB�c�,��Zj��I|��n�p̾b6�cV	�x߬�ʮƷq.?���HU+��m���"�&@	l��Gf'" �ae����xrBΝ���Y�A5��q��nt؍Xa��Y�������|H��cp`��O�ۖ��,00,�AN�M�4�s.\�p�{��7	�iZ������ʞ̕Eအ��4�;�}�<����C��Hc}�:L����KK�x/(lTX>��i$����"'ė�������=grg���Z���j�tkܦ~|lR�(�D�~�������t_�%e��8��*��?{8'U��BX)^��>�1b04�D�b<�[KY)	���v�	���e�'_X"���/OF�g4&Zc,f��?�����8��|������R$!P���Q�G7����*��uZ
U��	�\�	w�Ƒ�M��k�S�����|�T����#��u����L���DR\8R�ǈR81��q����0U_+�m�0��� `ŅC���G+��C����?4��\���"�m|̩`ґ ���ó�h��#x�{RoY�n�c��g���+�W.�s�Z������k�k�%��E�l�S�����s��]v�������N5xC-3Ԣ���eT������ʏ�S�ʯ@�5�t���o��64˦�C���_�1��%��M��)$.n΄?�g<A���xІ���Rϛo�o��lxܔ��ֵR�Y8�a�����Y31��}j�)�(�|y���q�ۣ��N�:E�a`�V�̭��휔?+��<%_m.�ajM��	�Q��"�o�Y;��tۤݏ6UT���[J�AOA�����m
۲����������S?(��t�������/�d{nŁt��V��~��Q�r!�'���%�d.�b��0o�VT���h1�Ǥ�msgF�&�A^I@s�vT��~����-A&3T��W̑���@���&VlOsw�����?cG���|ۀ��<'�m�fzk��YY�sV4�Xu^�D�)]uv3��p~��pL�RB��t G]/��F]L�.�d<�w�L�d7�e�G�pצ�]S$�^6�[��v�+n~�|%����t2��.��߼��-�:p�T^�mk��v63ut:r����ľ]U�3HɳS_3�yy}�j���p-���x�˟����f8%\*�@݇ۇ����ӟ �I5���Kc|o����ô˥I�X�TΤWYP��j��t�![�<�,��*tm��2-,�� eF�y�"�b��"�PI�(,0H	�+��i������%)�*A�|�x�7Vmҋ	v�@�xÓx٥k�n�/�g׍��x�%b;��~�Ek����K�X��eŽL�,�j9A����!��X��=��%)�b8��<~�â���������;�F��8[�djUP�&bZ}���c�����7%} ��<K����d/�B�;b�+�gŞ���� �M�v��6��g-�o66>k5_��5�R��P��no�x5Seo�t��(F�J�b"Bݽ\����� 9�?������l\��.l�����f@\�ÕP�B����in�K��_�m�]څ�r�Sn�ǽ৩���c�{�y�ٖa����e8J���{���CqT���_)�����B�y����v�L��e&mI�)�-����?5(����Q�������*rDy�,I��-��R*0�WjC�P�
��?���)��i�9C�^`�Nx�}�p��P�ߴr��{�Ϛ�:Y=
i;�z��,�Iq�����~�7�S�\��@R�	�̑FKJh��!�W/P�{�-x<b��\ѻ���c�bߥ���V��ϼ�V&���;�I-o)��}���0oV�w�>2��~���wHrC�v��(�/��D�n�k�e"֔�}3m����E�8c���$��#���9���+�3��$s�Q�y�ǝ��q_�a`�r�!?���pAEd�G\w4�E��M��.�T��Z=$�6w�����qb�m"��;'/�����u2\ȋ�&	``w�O��B�~)a�)���o�n�o3vO�R�߮��>��b��a��V�<r��.�W�s �`��wރ߃��'���jaA��V�ZL�Q+C:̪H���*�����o�`�'����`gv��<>���L
F�2@��G�!��Z�ɫp{�!Ԯ�D.E�M��_����� �Z��X�`��Dƙ���q3@��*H� ?�4�\���.��%��.&gV�/6�ZpC��o�q��>YI��H//7�l5!��"۞G��h���$e���5 6OP�i&(��p�ٖl[;�?N�I�z)�:�g6o�~�03���@��*$�� ա�Q.d ����8���v*nBE�̋��w"��>n��g~f֣<��On�В�+��0�4��t/��y���h��4w��24���x��_��x���%*r�y�ҁ����L�u5�Ap5�`)v�n� ��媆��E��C�h+��$��i��G�c���L�my>(ݲ��"�T|�5"cw�y��sdh92o�J˾e��2Z ֥p�IH �D��箕��) i��xܦá�^�w���z���2GS��]6 ��E�Ƀ*��T�l���".4�ޥu��Ft���{�PPB|�螡��T���wZ؝K(,N	��&�,��7A[Tݮ��n�(^q��Jt&-��%����#����\��kH��ފ�)/V�=�j��(5�m�?�#�fP�N>?�.k���9;���o�t\��l�@d�<jZ�0�wHKͣ�|�� ���g���q��9у\R����P�R��đ���\
b^:/��j��e��FF��lL�R� ��69�-u��-����S�wk�:d iQ��K��~���U{��2���V^�ʩwB�-ӣ`f�|�Bǰ��xId�3�M�g�Rl*�[P3���ްm����.�ET�O�\�k��[��s�0�&�����Mp��X�[�+'��й��T(�8��GyNV�.�`��N�FN$��/\ɔ ��wc*M�?d��p�^�Ir�|���4�4D��}'���\r��7S��¿i��03<5PÖs����73W_�N�>�쐯�@%��KS���(�W:�