��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_����m�e"kxu�Uٲ"#oB2�-g�j��h�p� M T�(�P�+M��&�[���+�=�n9" �2)g�ݕ����r��J)�a��m$�ke�xT+�ol֘B���zUz��}�+F�v�yC�V�`�W�#ƚ����?��J%!�i+���5�����5!���o0ٳiBk�욃�ٕt=V�騗Q���@����L�?=�w���]H`HO�����%���=�UzRG�m�ק�-�J�'^2�%������ޘ+��ؙ�7��q�̾�M�<Ul��z.�?p�
	tnM�F�xH_�K�W�+	������,R�$#[����ν=�i3p��YP'�h8��@#5-�U��r!&_���D�,2r;b�'{/wǠT��� ���ܑ�h��1����=������T<C೬ܐ+|0Y��њt�a+�.�Ya����$f`�E�>m��*�����vO��]`UJay/�C�>-;�$^�7~�r˛�9l~P��R���l���;x��/��u��s�&�u����4vG\!�=���PX����X�����^���������G�]����j�Pb����,u�,=��8�;�4"��D8��G�^�O�F L�5�.b��~<�L,� �7MM�>��LW O�F�G*4�Dm&ܷ���pyU�s��E��ڢ5��d�l�C�*T,A����-�Ը���qD�� Sq�\�Y���R|���6<�Q��>߽��z]��wB��়�ȣ�$�;*��+U$N���6TnRP����x�d��_ݥ�塯�����ef%E�O�j���C39���GO���r�V��gH4�vv��G���`�9 �@��v���'�~�2`��#��TnKx]��qr6
���b
�0S%���+��<cn�U"�+�iJs�kB3~��/b�7c�0/���_���H;�Q�5޸?� �O��Z�g�Q8����{(��@�=��g�y��ĉ�pTi4u�ew�EbI`��%�d��S���?Κ;�2�Y$�ٺ�e|��]l����[�7ᄲv
����1��"�]]?�C���z�Œ��w��	|~C��7)��Vf�.+~��]�>Z�����m�C��wХ�[�jXΫ�G�%S�]/��e���l9O�X�rJW|?��������4^p���cZ�l�R��& �0s�����"znCSt0�M E�c�b{I!�+�/!��5ׁ�֊������"?h�7��	�m|��O�)�����"�	Q	�+B��)��p�;�l��ݓ�M|�j����g�9���{��VG�g:rg�1�r፹�^Y�/{�Ǉ�%
��0�0Yפ�LaW�$kw͓�����j@۱��=�	I���DK��ey��,�1B|�ڄi6�N�84w��*D����a��XVA�9E��Mm;�־�M[�9��Ty���v�qb	y�KYQ��h��!�Nz!!lK5=Ϭ1�ݖ���F+�s�~�
�!��	ѝb�6���JX�
�Η����[`xQ;�9��C|�pm�'Rb�w����z�[�"^��F�A�Bx~����H�=�lζ�:;�ʚ|N�R1]s���?��%���߉��q��\��u�ںt9�K�Bj�(PbӍ�ѝ��J���"�p=�8�4�Xmaݤߴ����~뭞��ǛJ�7���
λ�N�����KPA�rz�R���X>r�N��XQ3I����1��J�G�qm���8�Y�2���O�h���o'4ض��e��sV�c��z=u�p�%Yf6�pOV���`$gRVá*�,S�]��7뷶�(r�� ��F%�X���	��a'��į��,CO�S��y�"]Ʋ
k����kq�)�m6��v���x#l���}U�fd�X*�R=^��2�*R&�����q�%W��i%�k�^��4�Ft4���1�7-̹WO���#�놲5��N�=ð՘�47�b���HqX��שLG��Mj3��#G�<��|gBރ��7�$.; ��G������S)�)�6���VAo�2aɌ�$ʤ��1U9}'MP�x���>S7��t���!&f�	Eyb~�VCx>~�'hD$�pq�����Ŏ6Ƴ�b/(s>\�D�g�]P�:�+"Z��Ñ�qU�XE�9?~��0�&{n��e��YK��0~��W�{���xb���з���<�9{�(̀��⋄����J��
���y�CE�ׄ�������r���o���y8Tg/ �D^��+��耏�͍� �Ͷz-�����O�
��=Ւż0�S�j��̳g1��e鍊b=n�P	P�!�fŘ����t"[�'�C��h������h�t#����d��`A@]�&E��8}e��6�|��
Cz�y{tn�٧}��+~�wJ$l�i�*��aE��c���/ރ�|TU\�Q���n�����oq��l����2CE�4��6Jl�N��`�_9�����K��4#��g��E��K�T;!T�a�3/W�6�f�t�ΡP���t�PU�/%s�e��<�-'��V3Q��Di��I�e�yʸ54��4,Iq-�/̩{����m�z�6�r"��<����7�V&���y;G��o^�GL�|�W=]�+jý"h��Qf�Gࠚj���0�ɥ'�ߣb�`@*n٧z��G;�NA�'Ŗ�g���=\˴)�N�?�o\M�e_w����1��J,�x2��9Vz���TNQ���gһ���.T��Csg���Pܮu/_j�X���\�� �A^�8��h �qh*_���m�O�iPIP�{����,U@d�����2�-FO�Ks!F��`���p������r�Ľ