��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�"��F9s�`&���a�oq���F�g�O�]�<ݲ����eCL��D���{�5��8̝DFI��Zp\m|Q��
�}�6C���UnF:<�jΈ�2�����<����sf�k��,jڙ�����2��X��Ss�HL��	�������+g?���N�Ż�����|�v7�{M��VNB
��Rs�゙�Ld\��X�'��R :�J���^�����kMkx�Q���3!P}�e���Z�Y?.�U{�RP	�)��lI{tI(S
7ZF7��R:]��Ѥ�>aE�-�$^D�źXr��}�C�]��c�1�\��,Aj7����C�	�O�s45���.�,���s�y��Er"*�X�C	w�l�SX��+��.���v�Na�ᴚ�b��ul��TY�l0~���M��(8�T" R$��T�7z���i�1 �X��֨��5�x9���9�"�O�5���7��*[T��Aw�2&���1K�w�+�w�WD�S6�0RߜJ��T��*ڟ���=(t���4J�$�H�Y]���լ0{��9J���q�K�i/޳s�Ƥ�O�qc$Ei��fP�~��2u���>��;~%��x�� Ӎ�x��IVa�+g�����E�)�mS�ZN},�&A_�p�>0}����!6��%̋��N�c��R�.����T��8�>n��'%�Δ@v��nϥ��~�"��>��s�@o�Z��W ��Udqi����^Dr�l6?���ֻ|�a�]g��Q������q��Y�d��V��j��`�2����:�Hv�H��Je`+犳c�P�r(Nd��u�#�:�g��W-N�<BW��X@S�uNY�����B���@����n�FU����B��H��\����T�rn~s��*�PJi\eq�ţ��嗘�6gC���6U�/�D�F�vK@�����F���%�2�B1@C�g�|�ܑ��$~�u҄��D����s�O��'�y,�=q��q}��!����I�װ��Y|��dJ�|bmw7��-&��-��W��-��||��,��3����.l�+S�3o9��N������c3 ����Xƒ�Åi�(Tf#ڎ�m_�ðMJw(�2Ȑ�`
�Oh@�"g����	��S�S@��y<��J*��������vu�(�s���7`��9_s}a ���HGl�������P�˕�/�c���a|�D��$��J[�q�,w��qQa@�M�hH �D#<93�R8��=�r����I%zY������h>*i_*d��h�E� ���dɅP��z]�"�E��>�������� ��Ǆ�4�9&���_)�w����i�GX����}����\����Rx�XE�_9��Tt�D��l7���!�^�fn��2���f*��sÌ�*�\��2�����3'G6��?뜋PV=,��ߘ�F,	�:��VR�ܕ�X4/n���y��S��Vf����	�����^.���d����$ēj`S#+m���RM�?��u9X��wQ���=�K2�8��E^��ݷ����k��z��J�h�D��Bfv��ze�*xs��@����w#�����D�ڼ_��5/�c�L�/���&W����mش�RW������p	)Jb���ɜ�Y�i�b�����T`�fCI6Fܼ$��B�����z�K?���,�P��|Z�F��hW�}�jR��e-C�\��<Aي��d��D�Y���L`95�[JS�}_PAK�cٸp:M�O	!P�_:�a�@�������5��߀X��9�0坧���&X���ŕ��!����N�{d���t�k�ip��ftz�?�t�F�w^Ē��h�r��-d��ᱱ�Z�{P	���W�֟���f��������彶���ڭf�M��͐�<���6��,0N��W�-cﬕj	�K�C�!,5M7�T�2-B�#0Ҕm���$�ܕ�r�㖃ǧ�d��G��#�q�[�,�h�il�˼'�n�\�\v#l/�6|�u�y��8n�`DS����k r�3@]�&3��'�!~��rq:�9�Cy�+d�ѡU]�>�QK�,p��ԟ�5��Fe7+��t�ő�YsZ\ϲ�3BO��%:O����^ܞ�:3�y?�`"������-�̖c�~����,���~���+<�r�]{�N�@�9j�.]��N'U�&p�ţ�k݀��t�0L>�75�������9}���$
+�Yy�������Xی�Sޑ�y,�ƠEk�\�sP�f��	T��Yn��v�5�H�c��-���<���o6C=PS#��ÿ=�$� 򁠽{�OL&A�ҏF���Ҍ��Q�S�G�7��ޝ�U�1��t��cgp��
t��ǚ¦B�tWD��0�r�:���,U:��DdJV�� �;���%"���:w@o��o��
	��b]׏],�`F���Zs�w��&�K��T�'�b��td��t���F�+6��<R��Tr�\F�����*k�����cO)k�c䋲<��W	1dw�����S�LJa Ħ=�T��n�T��?�������"�,���#[�8j�8ꍛ)<�N滑���0Wā�L%w\P�i�2.��q]C�ՠg���� nS���
w3C�C8ײ��Ua�'p�a#���vċ��=NKԏ�R�N�ҕ��Շ�nNy�YmllTb6R����DsS%�~/��/�#�ۓ�B�,��d1��w���{zx{�n������.�v7T�7�׍�ݴ����'�I�鼛a��@WaZ�j����6�x��.eFgR���Ɲ�����.�UC��w��-��`���i#��x\�U�Uˎ�:`6�G����,c��y���z㼳#h�.B���ª	�x�}H�խ�ًA�]�%,�V��r��Z��䥽���v,lF�y!4�]U�?E�yם���/�?�/(���歽�L���S�a���_���*�1�w�)��$'@D3,'i�z�#�Q�(���*N�2:�S����ºs�K��Rp9\��`�`�oܦt�uZ���r��6j[�`��;tSWh�Wc�%��[7��X��2�qd{��J{�Kk�\�/���|���p�?;�FR�Λr+�>Q� 6�4��v�y6T���Rh����[&��#��ҏ�Q�-W�v��*�2Vj �	[˂�B��\��^�Ҡ�R(˶{�$�Dk�k�(�!��í�z��u"(
��(�ڼx�ݹ�74�!Y���ެ9�E�,��vU���O.F�G��YP�"1 2�cܼ?E��ۗ��w-�`������`T�k��=z6Y�"���:.X`��&�@x�3ᰢ�]��sچ�@cY�Z�r~�ٕ�զ�BR��ia�r�5t1A��ި�y\ !lG�?�CȰ|��E�KAAFӖp�Y1��Ei�Ԍ{/��B)'�dE<V�+�K��G�g�6�o�.�K�~�{	.	-���R��لә�uBO�y>�DJ��K�0*�9�����ݨ �C 3��5�+�{�!I.=�?Xi��S6f�^:�1)��� ��ؓ�VbA��KlaJ�׍��Jt1�FQ��ߣ�\��C��$C�^���mi�ܢΚ�2���T!g�q������h�(˨�P��G�����Ug�#Ϲ>�r�̗����BC��wW����y����6,�����B;e"(7`����<o���ic�j-�R���Gr��,�-�zL�����>�Is��+t��2˳0S^��o����Y�O����5Xc&�I�/�܍(&�X��f%�*��k#)`:ߙg��KF��Dc�|-��@ݡ���+1��+=e�Yo�wr���x:�D�A*w��+z_P����{衭��7>��}����w��W��Ε�Ο������~=�����R���~���7nLlr�ѱ��}-;��j���`Q~�����χ�0�Gar`�� �4��FR��q�X�ove&A*+m�?g}�o�=�抻�g�	��S�]I�p���fd�>��B�L$��o�*�hpL����*(����{LG���8�����@:c�[w,F3��LH�]�A{C@�u	���AXֿKN�ML����&;FoZz���o��kj���
/�:�%���� �ᔈ! R�0+H!�t#���y�-�`]���9�����'A���أ����,�=r�����0�GyCL�éN1�g�3ۮNQv������I2@�x�罈E3����g�����]��O����
5�
�����yu3��t�\0�<�Ѯ���A�#�=n::J!Y^l������<YELw������F�vq��&�(7
A,+�D�W���� �{G_��;1'�ۣ
�NsK-%0�ai�gE+I�e�Ŗק�i��3�6zƒG��`1~t���X��,���f8	������s�Ўk���iF4S��G���ؑ�i�R��Q��@�H�Tg-����g����!�����|~�ߏ���hh���5���>����M7��*_&{B�Q�A��c�����GU�9�b�X�����S�]�l��{853�Ō��-Y<�@�8I�E���ɕ7�)��f����x�P�4��t�~ܞ�S�6�� q�Q�Jw���Ek��.b�@��c�%�ښ��5va�5��We�ŗ�b���P��`�� sa��*w�v��5�.��u,�
G�}|�Re}8��j��d�|)�YU0���g=?��k�+���w��\�W \⋒X�V��#��k~�b��.��\���w��m����Ӗ�@|4Rn6���Q�n�p��&�e�C�Id��e�л�����q��� [��6��]o��!U8�ħ%_�ʱ6k���"� *�T��V�Z��I�q��,Y�0�=:�HC�V�C��-�_.?��z�V��?e6���-`H���"����deBT��Q��R+�QpsW/�L1	p�� ������(�r�:��shx=��aH#���r�0s�c?d�a���I[Ћ�5��թM����:`(�Rү�-��O�C_9���klv(�� ����#"����D��}����`���-�x�h��f��.��p�<���:�	��J�8צZ�� ��F�R�j��;�+0���GL4�ߴ�����lp�{�	S$�� ���2	���z<������Ĵ���D�����59wM@�sG苝BYH���&����/Mc����Ա�0��e����>Z�,�{gr"��>��N��3��_]�8�ućT�I�Iդ���d���P�~�8��}���
�;�i�YT|Dro��,>P�ث*��ۡ˧�^͎�`Q�.¤, O�?O��b��5��yHc��ї�a����c�-�PIA[����+f�W�vE��ش�vhO�����|��k ���Q�K=�qD~T�d&�$�6��4��ex�:{�6F*��sܪ��{~������������V�d����"�O[Ũn�v;2N3꾑��
��嬡=O��({�a���{��VLت���d�ޖ�W0�`q�4	�4� >�k�s_�m�"�&.8%`?pV]�v=ߵ!��n�-�n�L�@��4w�F�b�����m��R���ˎ��y'���2z즹o���دZ���g4v�:��̃睳F̝�_NƎd_Y�!sp��4}e��@T��46��u��X<�V<���E�a�����0cO[��ψ��}>VAH3��//�>���D����SdF�'����²#��۸<\#�b#b�J6y��O+f,�u[�~g>j�@U��J�PD����q�]�>LW�vrS�m�x�	钂�^�5Dza�j���1������i�#J�>i��r}&�I�$��y���`94�G���w���FH��ўN����(��2������`{��Rة-��3�NNk���:�������u#�Uz��2c�9�IJ;��������UG�L���o+Y��#�eT�N�X�x��o���3�=O������,&�e�3�� ��s���@.o��jlz�����uI�a�\ƝĘ�q�W�b��H-f4�Q�g��jH�ޖh���0c�W��\3��^	�=S^z��i�GW[�$Z���|�i{�v�qĢ�]9������N��I}�3��vо�����Ko��eO/���U��:�c�v苁B�xS�*K�Fs����R�l�Q�:E�o@:/�����3|�{'�}].*c�ÛK����V�7�vˊ)wSv| #�7��]��Ա)-b$���DN~A��L�H�wÒ���Þdq��=�� �oY^?& �Z`�ؔX5V^�}mB)f�O*���/ d�6N[������钠w��6�?Y��QH��eP)��:QqJ��&;>3�S!���j���/ ۩U����T��O
hy�7hҞ����{��j�2��4 �����Ar-f�(�Q�::ֿ<��3]u��!oY���_���73nS��
�t�]8=���!���~�.$�W�
��>O���o���[���J�ˑ��(E[��k�3�)4v��uI+5�i�cX���ު����r!���$	�ʅ��G��B�8��R_	q�5�\�_$�%�81Π�w�����2(Sq���H8����b>vmp��L�����Az�Bb�����M�{�0������W�ĳ�"�1�2�qV���-Q�p[v�B��/�@�DRKW��=2�oB�Ϭw����_�|���w3EP�����CW��{�Y�E�M=C���g�%���"cW<ʆ3U�	>�%j*���-�ã9�zet]m�Ʃ�=kC����Zm?PHL�U|\��o�S��13DS��]�OꝞg:?e"Vd<�=�H �Uೠ�wNC^q�4���a�I8����f��zД	�GK��O��2���J�zl��J�90���.%�B���^���.^�����w?f�E����4�zB���I`]n*�0�D�C����>J-?�S�^"�v��
d�G�摐�K�I�=�Y$�Az�m»V�
��y�]Q7`x�%�7	�7xv/u�nż)ЗR�1�@�SbU���M|c�}�N�����7Td�s����$ܚ���c��k�7�&{�����g�Cf7a6(��i��0�hSHt�õ�;e����&ldds��3��'	��e�`,�琞Ou�jdU�a���9�w߄�*m�]H��c���rZ�@p��O����g�&�8�͠O��S��Bsښ7�_(��a^��g��ar�N����N��ub��L�ސ:�h(����QxJ�s�*u7�*o4�����1�0<W`���G?t�0�&6��<T�3���Ub��Ƒ5-�{��ߖ����pv3˦��%��9]����8)�8���#��'����%5��e#-�a�U�׋�p$��m�ܰ ��ex;[v�yc��+���w^}���go��^;*t��'�ơS/�����7�s6	ɻ���"J�[,��g��Hҝ�P����ތ��#�k�����#C���� c���#����Yj�H��M|���Z��!���	��H�w����i|��j-���&�͋�������{u-,t�aBqW�:(���#����륑�L;�������`+��9�����ż���� Df����͗d��A��^T	��#�<�1�Y ʛ80��0y�ٗ��: �hr�_Hp�Ns�H�֐v=ފ��&�l�[���7�Z��=����c��4nw������>a�i��j0S��x���0ރ�Le�L��+��}�);��7�V��{�`��V�M��5R� �6��u�&��(H��П��'�����?FԉF�l
\��Ƚ
ݨ����}2��&0�����OMIw���y}59�rSp�z��h�D��C�o�S߰�+�љ\��=��M�n9X����K�=_	p��%
�,�U'e4Tu�I�}��2p�������2yZ�����ɕ�{QL	�kNU�x9�
s �	���t|�8�7��]�0a����B��`qŇ-��A%t#��;���NFgjĝ^%E�ե��� JO#\�[U�S~@�И"ż��!�Z��c'D�X#�^���)�aB	��p�#}�o�R��#yD�a�,Z�pؐ>UW���T^ш�pr��%ؕ����� �F��W��Tm?T4��F3pP��	@�V��"�:;�s"����ћ�K	t�!2�8�iI�(�|5�1�h@�P�༕#(�O���L����)]��VZ�4oQ[�'z0�d��L�3�t$��Cr�p֣
_>-`{�`�Y��P�hY��Q�F��j��*xQ&(��9f��%�՗�<V���Q���G(��C���ꀎ��V����PߵK��b�:��=��������*�P%C�K	��A��-��@�΂��G�$������\���c��W7���C�X�K��Y������ �[1���X<�3O�<S�y�Ş+s+ZU�]C]B��M���ֳ3m������K�.fp�X���T���l�
ϑ����d�If����(َ��F5>��Dg�v�gUE"��"�Km� T;��M&��3�~O6��Lπ4��g\��y	8����(�!�$q�79���0�������p�|���X�ȭN�'W��v��i��u�xOG��@� �)���V"&�i� p�N�l��j�/>C��p�3� �D���=���欜�����yWY���k� �N�GY �� o�0PB�δw� ��X�8��ZCk��ط<j�G��+��?����v�_u�������.qW/��±D�%�>�y���g6�0�w�N��&�o�� J�1�4Yb�s"2�������q���H��!��