��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|�L��58b�Y��u���ۭ�E �i�s�D�9#3]w	�B��(�Fͤ`a'z����1��n��n��oD�DHU?K�N�<�].�K�3��d}�a`F ����.5aE�?jR�(��_�;�4�`P�VG$溒���UK��1;�+)��w'I�Ҩm�X/�:$Dv4�XiZ���D�̠���όr������\Wb �U[�=H��a�b��g�~j����a����¤�+�A�ilCN�鬨�P>d�ؾv��꪿.����p���Yl��S|��Dp������$�0�YXIB4��y~nQK���כ;ǿӾl�<��8\���5�<*�rBY �h�-��M!|�{�uE��Q���Ww���aA�p�������1;k�#<mP�X/�p�U��|����!_��{�#���m��C��5m3�fK> ��G�%P�t�:��l�����.ِ����/{-�� ��"p�¶@^�oC��ҷUͲ��.7H�
��w�NZ���:u����h
����\�F����X�) >����J�����X�C@���Jw<�y��PXS ��W��������O(��U�I>�vd��bXȵr=��*E��I�(�6�����ͥz<�"����#0&�>Ћ�<�S����Aڡ���0���d��dT"�//jR��xI_K��z����㍗8S.v��̵��&��D���KҴfO��'�І��*���Q+�>��^G���kn��-�ҧ��E�>�A$�ۊ��ˠ��,���̢�N���
1�;�g���T� Jy:�JGl���MZ����?�$����F+���ŗ� fX�4X��<g�W*M,���� �:�SSu�C����v������������wTUmY�Q�a^�n��n�7C�w�5�A���e�35^ʩ7接8ƸG�T�wl�R쫕���Fw��1�"�a�ﮦg"�l�
H��m`V5�"��,���"�p���H*&1'�x=e�`�>�}��x���d�6x'w��R���� �(��������N���u�.P�֒?�7b�mk�2��C^N���\j��Aiy?��V����M%k(�ѩ��=U�y�K�V/(��1��n;'F�No��YzG��1kK�j�GQ��,4MI�b�e���(�m��Bx�l� 8�zR/Q�$+�'��$V�=@`y�����5 a�����Zq	":�������W�Pm�ˠk��e�X�A�ի�$�A�����}��U&v���ea��5��zy+����I����>�N9v���e��EDO�&��e.n�g�?���C1	�����"��h	��1��Y�ć}����[��Ǆ_ѹ?w`$T�fe�J0{�@�_�Wy��%�#��@-ޗ�r��/�z|�R��7�8
��-�Ya)ܯ�e��l_��bR�g>=�ڔ#��x��Mw����S�l�|�D<j�k���m�{\�/]%.�©K锟����ɧS�c�T��q���)�Q����ڐ�P!c�������Wp=��A�䗞 �cu��J��W����4�� �{#8�G�x�oטO����7ݸ-���g���s�d[pK{:U�_ ���P׳�t�%+��V�`a�J/�/�������'?�EV���W<�#�c;���1Wr�+��:���GJ2-q ����0�b�=�_���L>N�-#�?�|pN����� xN����q�*XXi����;r����jJd�s���W�Q��3��f��C_]��Рt����F���|9?�vA�����ʹv~�v�޻sd#⽾��"�1ج��[�提���4������ݪ��]�O��f�-� R+{�0�_�S�`�>'W�X�.�prr#�����G���!N��}[Ѥ�&�w�9���I�kn�A�s�>�ɷg ���?���IF��zai�Q�X��ӻqE�lވ�H�?0`��H�"�Y %Z��A"��Zљ��j=v.^�	��i��q� Ո�Ь;�c�:�s�C&�g�E�=��\���WU0i��݅m?��o�NX=��6���Cs�.��t�q�Q\R;ibS?R_Gr71\M�S��P�\z�Y����_펑	(����s*b{��"�2�D�&T%�'��B��U"[0=�(�w��#Y�\�^:J�}���h�>��k>\$��`�b�������?���K�#0��]��Ib>�l?װ�y�א�CF�g1���cw�;e��I��L��A���w��A�K�@�X��\��(�h�tO��;)+���Н'H�s��i��r�RSt��Aږ�0�.�S"��I��F���{��u�0l;�_���)%��y�������Y#�� �E���G�������?�L��>,����k���V���[Y�N�'����6����734�^��ۯp�T�؝�����UD!~:�V���y`6F�tc������-y�v�� �+���]x_��OM�N/�wpBۿ@�z�l�\�$�<����xhb�ƖMoH���w|$7!�#TB��	n�H;c��<�/���b
@KJ~��O���1�uŁw�p!ĺ~�m�ڲp�UajG(�;U%Do���26e��� Qތ�NS����~��Ě2���fT��H�g�����+P(�T*�qJNk[:������f���5&�ҟ�w�=�-8,RR`@qș
�����F��~��!�l��$� ���D�P{Tb�3r�/����_��(�kK=MV�b��o*�0!����cɊ}��{0M"2u����1fx�GԾ���d'&�l�e�ޡq��q���;WD���T'XV�S�
lq%f�m����� �J�kxd�ݶ@=IhB�p:��Y���j���ӛ���8Ӌ�ot����^��h(�nR�����2l��T�MǪ��WgE�31�O�[n�=��
 ��o��"��p�exUXn�������f�f���,��.
O":���Obź���KH�ʲ�)0����X�?�C�p!F�a�����{�b�ril�R�\c�PЯ�vdSNM��q>��n+b��.�1kڭM۽���^WE�X�#윮�B"f�m�6�He�ی,�X�OFI�j�_W���bL��3#���o�3���p=�h�� ݸ�M���s�~YKM�-�й��vE$ ��v�6V[t�N6��$$�� 4 �쩛E>��L�
��I� ų�Q��զ?2��BW�1�7�	6�Oc����:��F5�p�ħ����&��jEy����&�u�|�zX<�X��2�&us �*����出��+�U�ťP��6+��0������:��r�,_���}Q�������Δe�2ه��Ҧ;^>\