��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P��v�"<ߞ��&'��k%P碶�R�ӣ�sĞ������FY&Uu1ڮ�*P �V����7�����F��8G���l��UsK?lM ��ɱI�:�8�ʭ�N�Q�)����mPe��Sk���ޱ�2[<b�b�&�p쀂��7��ذk=4��F�>h�r���sG��<�[�Vv%{��f���r��[ ��~���Q����Ż��Pd9Ƹ]���'�e3+�{�Q#�^\�2�Zv3-���˱����U�@�H/l�l��d�"���F������'G�@���g+	Q�"n�&[y��4ۡ�.a�2"T���jy���k��Q�3�s�{Qv�}>�^EŁ@Z`����p� @%�#D17s�F��"�DMW�{H��I��J��U'�PM���9-���{h�7.+	< ��G�o�?J;<���h�h�(!�_��);��EsH�i,#�z$����5cZB/Җ�����T}y���|#�[�Oϳg`-�i�2�d{'�@$�}�}��N���-����P�o�=/`��6����5&��84�](�i'�GQ���x ����$��J�����Tn䄟	�_7���i�Ao�gKLj�����
 ��y�'c�7 
�1�P�RB}���t6��C;��є�+R.{�	?,��R-�Ӫ��?7��|�'��2|�'n-@��k��D��IH'h<�iHd��s�=c�Dy���&ٔ�3+{w{�|3� >��rѸ[.`>��$�Կ�)��O�9Hv>#�	�o	�� ���ܨ�eu�L�4V�O1�|�4.�5���U� ���;�F�A�	oQ*�Gȅ��,@��?�4e��~��C+�ʶ���Ո�>��0MG�
Y�6A&ي4��P�}2��N�ZA^+�J@��R"�3���r?K�;��t��5��Na8�!g�;�ߵ�Lg�']�|���Q���6hT�!oqTHO�f�D�j�鋗Ĳ\�Si�`V���J�{�b�`H9`�i0Q4P�-�����"�w����3<����]{ΘW�^��)G�Mb�h��"B_�OվJA�'�@�v�a"�s!���jX�2�������G�`�A�a����EŨ�����ڗ덂���u��f'�F�<X��r�`���&hu��c:Ǻ�`rɚ��Et�V� ����6����1.�����yr��s����*q2J ����K��h��d <v���> *t{���i�6@���Qk%�ǪPG���Ev9��('��4tQW���m��v��Y��E����2���h#n��,�O�e��NT*��~DeK*U��?�c�?��freO.y��I �ﾺ6h��_a2�ߏ�$C��sg���<��;��\�k�~���i�K�:�&7&�1�����~8�mP�ϋ���A��.˝��X�<�0N�,0J_6:�g�P[Y�a8���h^pv�F?r��=���2���DVb�D��;�k��͊���)iqY
cU*�|';��L�&�%�j:j���F��3*����s�eH�tּ�����:PO���b�U{�]�R%S!�CV�3���ӴŪ�["���~��?�S�8f��bLʜ4o��5�{�,C�S�e��t���j����n�MD�$�����������w\���֙�CԷ��n)�}�[(��f}82 ������[d��K�_�g�[�"&���.�S�wD��y�7	+A��F��T���e)|��ۥ-ٯXC��Y"?h��F�[J����WS���}E�P���~�4���}��\�cG�4���P���d��#�L�,|XeX�Q�\`Z(s:�g�_-�A���M%�����9@v'#��ﭮ}v1w��=�x��$?\Չ[���p`���L���~��Ӯ��'&2�}b����R�ů_M�i���G�;(;Jz��**�ܜ���%n?�t�%8ĶQ�d�j�|K�����A�Y��y�'zk7�5�CU�,C��<'x~���(��ƽ|-��F[Lw�����N8G� ��n7u^�}V��jT;t���:���u)/��� A9�S��Bq`��u(�V�X�z�ɔ��6�d���Ƿ�,kI��Ș	�h$�L��!Ai4	}�?�����:Ç|�q�P��T;��ƍ�u!_A��}1(����ӧ"QM��H�z	� )���ޯ�z̊���Ld&����B��[p�%�*d�b]p2��I��S��( ����o�?^Oҍ3�h����_��c8a%�����'fSn(ex�Q5�im7�j���kgeH?�II�����;`�a��(rĉ���ǢD� 	B|�AOݠ@��jWDΠ�z�)�cj6(X���B����ܨFދ��O|374(���md�5?_P��Sc��0��)�6���v����]�� ��V�7.ŧ�E[��<�p$օ�?\kn���V��10�j�K{��Q�6!<c�e�	��w.J#4M�c�I�F��}hk4@���W�lyt|��3���l�$�л�u�t�i�~(���B�������hY�s%�6����i�����YgHp�((����)�e��b�<+�ם<Ҹe-L�_(8�\�݅�����t�	�"(�������h�S�mN��Z+��Z�ΉF�� �lm��!�� ��5g��!�a)��xӯ62�sc�bTI����K�Y��C��t�W&O��[=�����{K��w�{&�#��q�h�	�"�'�_e��dkG�w�3;���u$�� f3�NZ���v�!�м�����J�!��wGN�`+:���rV�*��zU�C�}���f}@���I��(�A:�ׅ��y��1&�7�p1�ӵ�PגZrzǼ@�I��i$���L����"�y�����C�\��ՙ���g���3��8Hi33\~�`rw_n������J��;Ep���sZ>+�R����R�z��`���x�-��*�?�y�@����9V;d��.�}a�H��]�KDB?�q�F��Rl�=�;�SW^�Ȝŝ&b�����8��Elabp��'���3�G!;��^�.�4M�F��;SZ�0�JA�a����9l�D<~'��ޛ�|o�	;%q�/�N8�����%�8p�nKxw_�#q^�:�'e��;�d@�*3����8Թ�p~6�оS�yv�唠��Od#�9���͠;��z�;��=O�]Γ��t�vgQ�5	����N�K���ދ7����Cx�<%?����!tK��Wٴ�@۹?��X�	��q�+����Zh�ʾ4x�1=�>�-'�����J�A��WJ��)ܜ��9�P�>8?b5�!-����t��+��tv?�.a���h�G�?���p���V�*�[k_�22EX��0�����I��������	%�53G���~]��}�-=9)��Ytm��̋ό"2���-Jx����8z��J��j�+���+��x��!J�v���.�`&��9�px!='�D{ћ%��x����[\��F%[$� ���w(V\��;L����Vjas�G�%�ݱ9���T�O���ei
��#
� ͬ�fNwO�3%
��g�aQ�����D� �"mAe�-B���C²3�D�!�L��T���/k��:����k[����M�������{y����kg�/rS�A6�'X��X�z�� �V�]�k�Hox&ľ7�*��x����,�6��ʹ^�.:hr�d*�]Y?�ڎM�+P�3m�+��cz j��a��u�i�d�����
��k@�(.b#1�sU֟[K/�� ��sֶk�C3ܘP0Z���K+io`����w�I|��]����0Ͻ��B�TGf)���x��߬�+���:�	c�P�M�2�Fb|�i\쿆N9ύ�=ʦ�4��G0���GޟqǺ�ԎRz-I��+�'�s�RP�P�pq��1!.SRaP�O-[T�pO��07G��~�3=�۸��	���B`=�m��I�)~�<7_V�G�A�ܚ�W �f��QԢ�@��VM�����3�7O�!��fw�@Q��}ݞ���O��/���.t񈸤�y�3
�����<�fJ[�o������u�m����*�,I1��:5��I�襖����̖�˗�=F�t0��̷�/#-O�F�� �5��O�7�t,�|S%/���'�y����e!G��(8�x=�|~ټ���2�.��-��6A�9�<4����AH�r�ʥ�U8���4<��kn.��+���M5Ajz��`�ۇ���f
�+�뮶IV�Ot��π􎇖�Ě>Om�M��"�#˽�.T}fzuY������E,VXf����'������H��Y[=�����K��oFD��`��w�S���{s?�Bc�)�k�w�YR6�}{m�`r�3˸�	��v%������(�w�6y���U$���-�\����r@����l|�iփ�{���۶�f���1�D�`�ٵ�gu�|�u�]�'��!����=#������y�Y�oԖ?�q��*��V��tk'7L��W},��g�q��ۜ\tX���|��uJ=!�2��6��~�$_G��
��}�#�J�?A7��fȥ�o��.�T�����V����5I����ϢZ^���2�m���G�VT�% ���	�N�njP�!�%�=t�7ġp=�� �B�`#Q�w��Y2��߄E̢0�C\�6�q��p���G�̀�=Ƨc���5���uO-c}�Ǚ��闒�5���J���3��u��nࡴx��I���/��ug���5� M��L5�S�����2u�5��ۼ9L�xl���ei)��~���I픝�<[h�٪^sCE���o�/��[s�Ef� v��q:��5��])5���qI��/����3i`B���M\�/t��bX|#����a�-��V������Up���oP��f�{m��q����_�ڌY�8���Jz�z~�Y�c�+��Q��Es�@�1��`���;\����3���v�>��p@�vs�x�9TI^���
�w�c��j�WW�[nV�:$�S]��*Oi�m
��[�pU�#t�{�SZڷc!?��<<��Xc����/��|�� ��O턺3�0�E���"��o0���H)�JW���r�o�m�b�K؛~�0D��n��vx�<��;�j*;�L���W)K��o�����^�~Z�Bҋ�ѹ8@� T���������a�֫����Y+4�^Ki��Lr��ĭĹ��b5���4��gZɥ3�#E�&+�j��h���?<�q'�Q��n���̈́=1Y��K
_�kĆ �iKX,wrbGN݈�Qҭ��r��k��NR�����-|u�+4�А>'1���yog��!A��ְ���kI��M�8v�ˈc��Yz�I���9�[�*�kAq"���sQ{���	�u�O��7	#D��;�7C��ҩSЌ%ƼA/K�6� @<\��^Q��ڟ{1�;p�>�8�dU%�;�3.:����n�>³>-�����O Zl��b ��I�3��l_����:6�x��q#j�݃D��ј}eI���x3�c}���M�(��0�J��!���7���C����ݏ�\�܇S���iZ�1��.W|n�d��` |�Q�[�"��t,b3B�kү���OɹA4Aq#a�\Q-d:E��.ǵC��)�:3�PCh������t>>�]�����#\���ݹ��������v��v��l�m�wt��K��B�q&_k`M̃�upH0��*u�1'ol�"�N���]8G?u�w�*?�2���ƹ��h�Y���_(�Z�ٮ�h�����&D��� :E��v��i�����e;��o��1�76�Cb�i°���9E�C��$q	����"�Ri���I�<��>1m���p;j�վ�����ź��@eHL�j![5�ŝ#-�E���ۅi�OCz�=��j�=$=B�si;8�ºR<�Pԉ$5>l����@�
��t~������;X�|���9!��5�Σb�^O�~�{O�Q��ݖ��ps�:Y�gG�iu�~:]~ =�ӏ@T��&B�՘`7G!C܈ca���.�ѹ9"�}�Ϫ ���m��6���j�t�4�H�.�Me-�\��"Z�|"��ȷ`ET��
�9zT�U�����@�/=ș��� �8oﶠ\�8��!0� RgC/��JY[�x֐��5�=)�ǚ��k��kC�aV?��!���R��<g
���K=Gz��~p�x۫4�A�ɮ*�6��i��o��jҦ�d�#�>/�9:e����υ��k��U����D ���c�����I��)L���YP�`e�F.N�xWF���dUx,��Q\��4��o6M���������ԋ~\���� X�
�#��as��,���$��NƤO+����|�~9ɰ\��e����N�V�&�iy��EF+{�C`o�$w�@����}V�l�9���`;Y��Z�-l���޳Z��/�!�WƇ����~�R�˅����(ө(c�� N�Ze�ɻ"�Q����H�8���!UG���y�y_x�	�"\&�h3��ajO0ٲ[\��	�|�H�����[g'o��k�"�l�ޏ�3"̬���9�K>��������ф�A��{Ox�~��"��B�l�����'E���{y5xp|'��LQܺ��X�W�BS0��˘����~\��%w�9!�	W���+�'@�v��k�+�gl��,u���B�S,��t�3|0�Cg�u���7���p�A����F��hX��d�����45�J4�ۢzVY8˝�:�(���h��`��[��CC����SKƀH��:If�q"SȨ�k���X�ЫN$
�{{�w�����%:��4qz�$�i���f���vE]�?����+ݟ��I�uP��s�w���!�훊*�a�I���>��E�c���_�*����JC��3=|\@��hk���`/�	�^{���;���o���r{��W�@�"�ڛ��-/�#�x���5#�G�tS���uit�kF[�//\T���\��X�� �h����kPw����q0��Q��ꋡ3�p�[��TQt����NA�ع�Vr�>�H7���L�0L�(��a��>X���J*�w�]Z���%����\0l��vA��� [����;g�mĭ�dX80��K�L���H�PG*��#�������t�`�Le6�깥8��`A]n1����8y�ֿ`
ބ�9s��5��32����n����GcT��S{�R2,��rX�ӮO�4�t6*�m/��)�w2�K%.� _�*X����(�\�s�W5�o՚c!��!��ߴƚ��yF-� ���ml�9��.f�lHZ=���h�9��i_!(ki���&�Vj*ٙ<���p��HD�T����7�~z�m1[<,>�Z���H�SC���͙�/�Et�<���$ɰ�)^�#�FR�(y�*Ag�VX�Bz��6l�r$�M�j�󠬯�X�]w3�2����S�EDk<�(���"C��8o�z~�]O��0�A�L�T-I���%����� S����7�9[@��HY�s�czpo�_�φb�u��X5�T����Գh����'�o�KV��}7>i��U�Lj���7�	�� +1|ޔҭ�q��A�S�B�I���y1!j��m��vf1c���5N�7��H�*�����L5�I?`)���= ߏ�q��w}�I�nO�!cKh�d\�F�~>���[�Pí����hrPq�4��l|��L��W�$�$=�Q�d	��i����u�`���J�e�U\��ɲ��p�R�ʺ$O����˰O~[P/$�>;>T<]�(���J�Y�ێ��� �����{GU�'��%�^.�|�rߵ�foYw