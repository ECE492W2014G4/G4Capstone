��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P��v�"<ߞ��&'��k%P碶�R�ӣ�sĞ������FY&��9*��L�y2J�ǰP[�
�@��ȵ�i�W�`�
+��T=O��h���e��ԛ�ѣ�s��|K��p+!Mb�\9���	m���>u\ ��	���b��*��@�צ㥖Ƌ
��x��m��~92 ������Ȏ5@����~:|b���ߥ�I�_]+�������u[Kڋ�K�,0H�UՆ��}9"��ԍ0!�n�z`�	d�,2:�d遛��F�,Z6m��;H���F���� �U��$]���:K,�1.�M&�R�&Z�Ə4gu���*�	�UV�y�|�p7E0�yܪ�jkT>�yV��OӘ������Rd��(��Z�;��Gx�{NG��Tj�����HAz㢖}/�6���ҔT���Z�~?&�v�8&9�Ь�F�����ӣMvޙ��6��=@M�5�0��rf,bos��B�Z|8z�R/A.h����&RZ���Dr@��u^{d��g&ǀ�\�o[NQ�f��&�	b&��*���|`��;�t'S�Z�Zꮫ�/7��o\�x�n�s��h@{b���E�_,�\T�����a�-)�T�o�f�\����xl2+�"�P�Z-4w�/@Ԙ	A����㴐~˖YB
Ss~��-ִ���M�/#A�
����Zk+��9���ZE�����-E|:W{�2UE� N5d�<�;ͣ��J��g�5�Q���e�ދ�Ec�DNt�о���bl?�7��ܘ�2����fRt��\�m.�"�(�Yx��|�����X(&f ~X\7*fL=k��$K���~z>;������r=���v�S��N+��d�:I����^sA>���?�4�<N�BX�(e����:H�aָ�����'�{j���L6~�R2G��6��HK�j��t����A"��}� �Ȧb�%?u���7ma� ����Y��Po�dF�3 |L@[�ѱ���3�O��d������\-O���p���F3M����膞��ܟ�JW+yY�49���Ftg	nX\;��eD^�80�[���3K��7Z!هS�i��Uv�H[�l���K����͙_ֶ%�L�V�
,e0�����=+V嬲<v��=�.���/���D!���@I��|
�A߳�Px/
E-��p��5�m!Vȕ�4�Kli���G�J�|���3B¨l/�!9Z���MĬ��jp�f{�n�2(YF!n�č���@�ύ	���&=�h���<��8;@�߃u��`�Q<ePgeGI�����+��ֳ�������;f^��� ]tM[�4��M=��sd�ەU���O��n1ڙ�s�R�u�����R!��ˍ�C��Ӿ!n�ZR�S�l�W�s��~��U��w�?gp{�A�e�7
�ă�j6�P��1��ѺJn����
�ʦ���4��o$jހ&|����-N�`�#�ƕ/��[헧�gzZ:��]Waw/r*��?��4�X�u�FP.����RYf�3�!���.�'��Z2q'gD��{v��J�׹*�p�lB�eU���d��H�}z��E��8�Ɋ��6��Tͯ.�j�a[�~��y�d�$���D�C��6<&�[ymp��T�}f�-��M�q@rcid�g&�HWX�<�Y!�γ3q}��#:Y��irg[%��ĈO?��8��O�5�l`�>�"ȡ�YUL�Q8��6(Y]�"o)�-,��Q৾�I��1*�8���}�-��%�i�r�^7��I���� �8���8Z�/�o��Vga����y�VQ"��D/�=��HA�bKs�jğ�b�E8�*o��������P̧TI*���ު�e7c�>����"9E>#���wZ��ς�ެ�*�6W�դ��Nc���vj[t��I
�3":��!B��7��ו6ndB,Z���Ԧ�]`@�OKz�gd�$��"Ҙ�Q��b��;H��u��eT���&A�`Nriٮˋ
�sIExv�L�Ϛ�u�����j%_����ؙǋ�l�/�������kt�vNc����/�oݕ����o�r�5MDs%N��� D���}#�����LR=�~ㆳ1Oא���c�B���H���X?$(�`�?@����^ϡ�B��2�������3���h��@��߮6q��|Ne���B�����t��À{J�l/��û��������R(�=!�l�9���j�����u=��f���`j):4�?�?Ol��{��S��z����@����J�Sl߳k f�n|SH���{��h� !��Ꞗ�7~�2�lMTK��>����R���H��2��P�s�a�=�el�
ސ��%Fź܇�D��rw��{f��p0�Iр��O L�����Y�'4�������ڬgn��ިIWOay�����!��=h��܍�`�Z�Q*}0m������UO�.l����\{�-$�Fީ$�z+���bw4�B6�L�
���T����S����,_��6��J���N}o�FY0(���l/6?CIf���@��c�&.N���D�ԙ^��`1X����%t�!���̀�F���pm�I�~��Nv���F�3�kfr% ӸB���3g*���7�_}�׆���Xx8�e���߰��s�1��)3\�I#�I���61��uhW��Y�%̪
��ꍵ� ����\C��vȊ{ޜB�!yfs�Jsø��Z1��Y�	��3�z�ȼ��g��V����cZ���#�#P���x�X�t;a]7���m��5o���%�܀k� ]�8y�Ɛo.�b�xc��w�;_�n���t���(��#e��E�t��Ј��P���ė��t���P�p7Ls犉�<1Y~�J#4���R�A�J>���D{1e��e��9�J��A�=����SP1G��1�X&�7خ����d��0��Fbp8��|i����Nx�Ii/�3�jZ_�:8ZO�.���]W�ք�Ɩm|n�yl��Y'�vKt%%����i�{v�T�{��a�gn�
��2�,�4c�	�F�(&u�4�ZMگY�A�ab������	��3��D��������m0�A8�P�_����8d^�-.�i%9Z�S�<Kk��3�����������V�Z��*�= @i��hP�����+�����۴�k�zH���1�Jt��o+	q����GY~�T� �2� 4M��S ��vnf|u>��Za��%�~���8"{�^ܕ��-z���4�qy��vl��kI�=�n�w�$yo�-B���f͂c�(���3̡�������T�Q��������{�	�ɬ�ft��A��h�F�#�Ġ�\��dW:<�^�+�s?��v�z�
�a���d�o���w�j���ݚWKJ
>�5=��D�K�x�Ϸ1�孌���7�%a	�T�Ȧ=6��\Ag'�۱��J�W��~��6̮	�*�	�)�gK �7������A$�,�6�|��B1q���6�o{U��9�sT��(r�k�E4˅��"�p��#@#t^��}�=)��r0�u7pǯQq��"���$�jS��^A:��D$���6E�ь�`��h�p���U���H�ۑ�<���Jv����Q���I�#M�����(�j=U�� n*�z���3��m��4!��ѿ�T�T�[sN3y`�w�,�߽!��ޖ*�HN�s"���}=БTL�����5�(	6]�bt,��'���p�;�����-:���[Ȑq5�����R�y�����Վ֎s�����8�]fPp��YF�z}`���Zq0� 'v��[~�WO3�����C�Ԭ��$M��n��t\�FA�9���%�4g�)i�aSh_r�������_��⟥R*��m��Z ���;P�ܱ�2|!���^~Ki�h��@Jǻ� �~a���3U�+�gAm�^�E>GL���¨��+�	'2d�X�O��E�g�׌�Tkqښ�%2}� ;E�C�c��Y�����s�Ä�̘��M�ޥês�
u���"�F,F��� >����J z�G�s��nB�,��*x��"U=�����,��F���r��A]����@e�譈6F�&`.L9�Cb͊Ju�p�N���F�b�i6��k��7"j�{��R��=Ct
���5k�>B�tl��>�^�x���n���k.���tO1H��_G �LR��"h��oN�V-P5����` ���xH�����{c���mw䳒�%�+��W�8���� @�C_�o^n��ݡ=����ӿ���k�����n��f�R�d����H������P���~_;�z��?[��ěiI5Cw��B��[�����[��:{�9݉g1��wٍ�2����#�A��?�S�BNü��&��iDOFhz�*�N����B�����{���@���Kz�d�B����5AP��{�$�v�������P�2'�����y�6·�{|t�ք�A$���M��
wbc��8��&�ȭ�>E�F"S��C�u<��{�9'�{��P��(��ߛl�L�5�ء
�]|u��}���RR�QUt�%�@,�a��t-k]���1~�068�,��1�yS�W�5�2�x�������ܑ�O���x.�����6C�!.ؚ
Bv�kS�0�_@3���}�y�����3Ԃ̤B6�= �O:)c���"��n���B�4����7������R�rv.�X�ѨדΰĂå���V������r� `�K\��$�;%�V��A�m�o���~-YN�E�( %�oFl�=\��C]m��aؽ�.�!۸���sÉ)�p���ʤ��flU�'H!������Z4vT��F�Z��I/d��o8�l��h����"��%Ȫ�0��XB����Z)!#p����
?⛅��Яҭ7������$�W��L	T5��P���E������f�*:4�OfZL����C5��{}�6�tL��捋��gU��(Q��(h%��n'% x�S_�.����]_�o
D��i��KrI�D�&4����<�g�5D֥aɽ�Պ=��Q\����T����04���3N��!���!MGJ|�3���8�Q �Vw�����J����1�ՙ�<*?J�ݹ��j=��{�mn[���A�Z�$eu�7�d���qc�\�q
2D<	�5�_�A}��ϗj�ٝ�iZ�t��Y�Pe�u����e[��ͩ�[��O�j�a����nX��'��U��0�A��g��	)n�.�?o��/@5_������$CJ���l43��Tb��^�����aEy�4Ţ�/��]�?D_g��'�߱C�ax�]!��݂�>ʌ�����Hj�A���qN�ۆ�>�I̍V�pzF�3��<����}'�I|*"^����6j�?�/� ����̅����OߐheO�,Q �E��_���EB|�S�ct5�H�\�����abǨ�;��C�N2�|��R��2�@��g�6q��߼��Fu:�F��t�rA7ȁ<r
�ЭO�~�~h顺o�I��ɨu�$,A���Gs��r��8,��yhj�W����+�O�*�r�
�M)vm�������I�<������9���4�(lPل�u�Ȱ�Y�i~(��$v��%\V\��cs{�t#���j�ƻu2Y�u�^����e����r bq� &��J���[�Eg�J'b����!*��������.=��n��}�|�
���٩b݆d��nё /�0u�˕/�Us���i�Y�X &/`Q$�2N^��|�+�xi3��-Ve�<�,������e7|�y�]�C���H@<�H_�#���;K#I*$��N�G��4QP&�)1͏	?Wf���ڷr�� ��x�/j�>K=���59��5�HS�ʒ�I�'.*�3�˓��H=�K������ʞ�#퇰M�it=ZE�Y֎��m���$���+��튤�ְ�R�X���u��۶�*I��&�rFא	����C&P8f�u�@�������l��"�i�^[�'gn��"v��M�u�)�w���{�ѿ��wbS��ZX���tz�E�t��\�BV?�x�|�-c�>��cIͷAr���IO��[eGr��h���;L�-�Ƹ?�^�N��)��Q�l�Sի�vZ�H�.؃��ό�4D�cAu��˱	ǯ��Me���=muD�Z�����3p����,�Çl���H"��YB����y;��b���g�/�)Q�A��.�0�	�M��\&;i`�=֟�����"ի7�_�7�{�_Oě2'�����H��$|	=�8�	���$[<�Nܪ���V}!�8K_&ʎ��v&�G���͓�tv��5�oN�`4qƏ �7��@l[?�^l��M��ۺe�7+DbeE0�Z�xK}��o}�;:+�%�k���H��]�3��%r����L�=S�}*(�o����/x%*��]%���މƗ|^�Y�O&9���\Z�����.B	��r.{\j��A��2:��/�X�! ��� 8Յ�f��H'��რ��֭8�m$ޢ2�[@�q]��̮�u����$6U%��>�n*�@0��)�Bd�:w,��.=�z/�co�����¤�dZT׌W���`�{'���퉷Ka(���5�ۅm��'gޕй.^�iЕq��x�ω�u>K�C�ѭ�'�B��74��XC�"�̰݇,��,��D�G�t�"{hR��)��euT�Fd�(9�8�=�|�~��0pQ%����*���Z,j/l�:��,��)���8r��o��1c6kHP�i���6V��֓,��:�C-��5���C�����$�3艥9���g�l��Vu��� d9#h�������GJBl���`�c�u�a�,�(�\��9�`�-#�����|;	��uھ���