��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>��`HX����5a8Sjfm~���*��
��3c��N����-��REK�!���tո�Up`��H�րS�E��јj��f�G�8�u�h�����8�WD{���CAJc��k^�Zi�@�MR�q�+��.ɏ�D'{��7�s��ͼ�T�Cҩ+���<K rM#42���fHK7���
�l)R_�͘:����@�ԣNZ
9�'@^nJqx��ӨK���`R��?�O�m|	/��ͥ����I���Q��� h�L�+��T�B�7^s�����x���=,���^�{�����;W��Ʋ�)�����9poj�����_�l��]�x\��~�����^E-	���o�f�"z��W�􁲊�G,�4���mC((��v��+/"`A��������0��	����������轴��D��� ��t3°��յ�r
�0ۂ��?��kı	�\Rw�{2'�\�T�$l��f�[&���\H��6��o1>�e0:6�!fH%X�bo��7�} ��c�O]�C���PL���iR[�m��ޤ_�!f5��ϓ&�H�����<..�4cC�s��C��4�k���z����'�Ъے�jȽ�%O�iA���y��s�Nn��7�a�]���v�w.Ҳ5~�����B�v8	�u̬��y���>��nխ��N,#U�OnYN��$�m�c9(�FY�O�2�<�� Ԫ�o�� �����Q/�f���h	_c���ѽ+��S�������j?�9Kt.�q*� ����x�����KC�����{��o���A��Ū���4�/gsC��em�?!�ҠU�f���$U+1am����CWC�M����M�������y�K���OjG��e+�ɯSU~g�����[U�(C^�}$!�{��i ��ϸx���5��J"'g����'�~�
T�y�7F��j0r��*ӂ��oW5W��&�P�-'�	� h[-�9�E )6k��Ÿ��m��p
 ��+ �Am�4�P��ӧ_�{��ʛ�g����C�]��~ϩtɏj��V��1D߱9T�6�>���ǯ��B#j0�2o$|kו �̒n�RNPY����"r�d:��w��=��q a�M���%<��M��-ga>Kq�п4<�`ު
�¶�Y��O�
�^2�8���r %����ҥ��2���5��d���-�!4�����?el���&'�K�g����\��s#mau��J�{;�����\����������7���k�
pӀ�����߼K<1��^�c8�PN���EO�m	έ��#��q�l���؊��
���(�8*���"3��T���J��u\��%J!�,E�{��1F�١S���G'� ��ْ�}���n�w�O�65X�T���������B��ae��J|��{\�V,�7��4�i��dN�����WI0��?o$3�x����;O�t��NS1�i�5
�u�](���U�u.��c��ʰť!
3R�a7\���O:�
��;��
Q�@v`��ͯ�U��^~*@W�"�^q��~��ڪE��C�#3�������1GgYGk>�}��WgߑY%י�2Rˮ2
�[r&
��[ƭy�����]�ͪM�.�����1����w�CC�*�IJ��ye������C0��Y_�4L�r��I{�m�r�o)��n�x�dQy[�\}yLzދt��xm;�Л�;�o����
�����`y��p-�paC�������CSB�����u�9�Z�?A�MXB6�Ǚ@�A�[W��]cq����!p�M(��lᙡ)I���yoi4gB��c��ŸuK��&�~��g�Plϡ�����vV�tmA��2?ۦ�y�ԲY&k�'�*�KK��\�	|��"є����EZ�R�<7�����{�������=�tWK�+)l�o�u���wR!���f�}�ʚ��<�Ո}�[��-�BCCT>�8v3�w�k�Z-Aq7�8 %o���o������P{N�Id��l�����nJz��Yz<%��`º\<�.#��\&o�;���F�"�w���<��1��%w�iз��a�T�*���'�~7�w�0��fN-���r��@��[n���Fpt�r�*��	��vA�ކ�/oŎ�Y��L)��sFۆg�4E1��Wճ���23{�i�_��o���V�.6+��Ȟ�:ٶ����.u�7�|�)�=��n"�t�����N�'��p	��ӕOB��֛���s6�e`�5�L�]2���t�
4�U�FP��=�q)���0��8u�VF��Es�;[yg����PT�ώ3^l8��2�]:'�"�R�@E{�e�f�b��q�O�f3���J�Z�x��	����9z�C��ȟ�%�		�&޹@���^�$�8τg�0�U���`D�;9V���f�}.�qxzxan?՘�w�|��C(�
]�$. �Eb�ZuW�̀�ި���@gپ{�tU�CMk 'B�<y�I֣�������'��e�� �ӧ2ėw��C�*C$7�=ܓ�4���R0� �i���G'���;�f�Qwl���U��0n�z���������TB"�OQ�{� �r��u�QQ8����M��7�_�-�������}��k����V��f{Ⱥ�n���D�s�>�L�]��H��:�~���@'R4�'�H�Ȩѥ�6-�qKlO��lz��f��2��iLy��&A�4IA�ْ5��WJ㴱p=O��R�	�N5ؘ#Bm����կnP1����)�Kɐ�<�s7]GC��Ș�{�9�����<�s��[��t��������ţU<խS�i�|Rt�$��(���ucԬ�H�����XK¥��!�q���G���?l��ܩ���Z�sR��lH�DR�Hw�Jk���:��ltzO�"n`G�U9��0KW Et�I�\�g�/�� '����*����΢�&q�<�o��i�wyU��o&�N��xh܋�gF*�RiW�'V�f�d�W��a��4�"�J:;���emO�U�_+����L/B���.��u�K���202��|��8(�����%��րTX�x�J�Ym��zH�w�*����n+n���},�U��l�#O07&$�0�h�.O��njbT�2���������w��B`)���pz�����1H��p~uex�fό��];(���S����=/7ߵ#��4�H�C��|�L�[pQ���J@���1�3�{���ӥ`�ٻ�nm��_���0�c����������k�%x�`a&yjl<#R�	��e������r�8�-Cl=�e>t��
9��������cR�-_ͼ��x��P�>��-!����(C&M�Y=�t�sg���7E�~DJ�4�(���Q�%����N\�da,��j���F���<�ߦڊ���oDt�7�3����a'�}3z���ς9y������V����n���{>�E�c�9�;N�������}
w�@�r;����L�=��!�B�MթE����{��hs0�����%�{�3I��ZK� !�Q�b�dz7k�2Bd� 7�Az/:�U�����M�T�����G����_n�Lz}�,/z7��~fE"�\`l�/sn�����^C�u);_����&��*�)o�w�e��,|��ܔ��^�[�magxf�a��h��z�x�l��u�<�d橱p-��)8��ȭ����(2x�;���}�D����	j����k2��ye��@˾�g�|q�=�6���޲-D�[�D��%�DaS@-�B,O���ƽ@1 *r�LQ0}��l��Q�r����	9�f��Dp����G���sM\�bm�U�m��	i�O�1�(��zV�KE3��^҅?Sec��i�jݐ߯��B.�"i(��E��&��Ym̮�^f%*��<�WuP:d�!�-!�3��RPN�~*A�u/ĉ6�s:<�)u��>��2`���7�.S�Q{c�����ډn��v��\l��.���װ�.�J3�寨�X��]���~�?���U6���@�2��{�Ż�@{��#V̒wս�8���"zmh����ƁY�� ���@_�K�-�S�q�!���*+Z�q��V"�δ�����|mdA�j \b=��Q�Кb�'��ϼ�7Fv=����6�%ڸ5o�'�T��"Ga�� Q�.�.����n�f(����~�R$�eַ'�lT�z�8O�Emmp��f�
��{��2W�����jdSP�#�`�L��C��f	G��Lb>O�)�oL�D���R����q�Apx���S�R2؉�8����`���(V�2ٕ�(�;n"�Vj���ݙ������5/E|�l��b�1����p=OG���4Giube�pt���yO�@�3�Lʦ��̰�A�'Y��r��y N;�����v��G��y�b�U�^���(8�e!E��a��'m�G8#�S�Sue���!WG�AxZ���(h0�S|-uI�`[�J�a� �**]���{�^cU(x��>�l��$�G�N4]��ɟ��+AB9���J����w�o���W�P��"o/sB/�`:p�"K[��I�;�3>���	�Ig�+*�[�7/���;��>���k���*����˯���M�	.�ş�XV�g"��J�����3���+C7�)Ӻbl]����f�D��R�Y�������pl�t��V�9IA.��x7'Ј�r�dK�݌�\+KO�S�k��0�zC���P��$�
��b2�[�w�v:-~�0�˗
���M�����/K����T���c}:�)���?J���K��|�̀�`a
1�l/W�7iA� ���J2����8��zM=$�e��'���bn1��`[����!�Q���5�]a����ѳ�>�o�q�K���C�-s���@S�	d�#���<��� ƗuN墚��	�_b���6�AԢ��^������ב�Pvc�1́���=x�*�)Æ�'jU�w8?^���R�إ@��U�|�h닞�03�-�C����V�'Ѯ��+�J�g��T�%8#�~��������l�]����ġ����d�ZmB�����_n���l2�*�.G5R���\���+�G_��UCX.�0@q�V���|S5Y(�ė�K��{%=�ثN�b���;�oz��4i+d m���j-�jΔq:ހn�=��
H�L����$�5u�Dgj�
��#��񪐞�;��D�|��y5�EJ�Άڧ�����]����T_#d��w�'�,{��V��sBa�|��%���AK��Ac\� �E�"�P_@��f ҭ!c�AK(�XBwbl�A�����s����ƾ'�� �<CR��n¬1���/��|ﰲ\�D�?���� D�UiG�v3���!ĥ�b�'ksqx���!��#R���#A�;įi��5���-�iU)c&��U�������_}M�H��5&{��b�ar�8s[�14�}�k�c�!SӰ&
�������g�*()�G{~�O����'��Z��M�ix�}e��\9<E���u�yc�Z��{VV�r��/���䎁��%x�ܠ�|9���2`�4g�4,1{#u,�V."��>��;=[*��rs-/]
��-G�_�/�)�S<�>��܆�"�ՕS����������1h+�h��J���j�w�(Ao�����V�I���?5�8S�����\N�:RΖ�ak������ҹPxF24ۋ�/�����Pһx�k|L�>����9g�(�]�G_z�ָ�ڔ�ԕa��(�T�7���M�h�8�����y��@�'¶�z�����5���k�OU�
#}&p}5qqD7�+��?c���N=_�O��G�\���aq�R�M�w&H;p���f�b4�mSg$���%��j�H��i�?�Y>��j��2��u�6�b�T�w,�s,k��;�O�ui�
EOXr������T�k��9����4�DĆFjƲ�Г{�1j���z0��usM�m�W����������Vr�}{����R�D
-(��!��lM�dJW��jⷞm��
��G�B���?i�;�,�G�~k�����]ud&M�h�@�/7�O_�R_�b~v�>-	qz��OQ|��`�c5����goK/�7qu��/Ը�˙�6��F^���cme��K��?�ޝ�F/�po)�'�O�گWţAs�O ��"� ��h�M�
n���/,`��xe�F2�񎊓����Z��Qi�e�-��6\�+0��J
2 ��H��C������*Дl�f���2�9B�|聇[Pyq��B,(G��t3	��~�������i�6�7#�r�2E,�K���<������H�3�ǿ�3���(y7���ˋ��T�O<��N���觋WR:��ݸl#<����F�a*X��:˟�m����r�a�57g���L�ˏ'�g�r	$��N�����z��bC�Cy 4�6�4�lm)ZJ��<+�d�}�+6��������^��w��*�S��l@�t��=�Jw4���*�*����9�Y�Pa��G���*��l�o�B!&v��6U�Xf a�=-��j�b�"M��ChEZ:�j�#6P|/��.�L�&X(&�1?]`�'�|�?�k�W �f�wʄc&|A���%�"��9qS?	�Y��l�{
�]SJ�g��D�/�=�A�WG��{#Jt'�����`٘�������(!E��{�I���oF팯��`���bL��y�vFʃ�ߩ<�>������.j
�"/���=i ��P�]�.�k��am7e�a��)Mt.����na�SX��5���!IEG��m������I<K���ێ���C�Y*��GD��>�QP?��Of2�T�����M�A�����C)��ck����}Nq(l��E4��$�\���AH���_���^O�{��l�����.u�4�I�y�U�&�#:��4�bUI����G�>�%��f9���:���~f��|*x�R-σ�Jҽ8{���:��y.��Zd�UJ{���"�� �����������`�f��;�,G���YP��]���Uw#`4�E���짨�o��0X�|�z���^�w��,4��]�MV�v1�ml��V�.]3��{#���S��Њ��98����Qӝ�'��捬촪�=�6j�L�	�>�/qe+�H}Cެ���!����c��2g�4��z���x��'-w�I�����> ����i��r��WEe-��k��-P9`�s���(�Y���W�t��k���uml:WĦ��6!�CіmX�5o#/�����g$�m�Ґ�잋{m�ȗ����s�5�,m7>$8����=�vģ�<r���h'gB�����y'���ߣ���^�����8V/�r��@~Wrڞw��ZcI�FMV�S��!;����a"�O�gy�"^|r�����Z����֮P�&��q��u��-�����V�շ[��>.;e����H5�4K�'H1��d%�#ኺψ1��M��1)�6dAF�Fr��������(��bd|:aT���j�>�R,K��5��Me�|��������!���#D%R]r���8�!Nq������2�ycS_BkB��i�=���=���Qu�Yq���Y*f�u59t�?�v{�D�7�Iw�^�u����Qz�z�@~�@2���4J����-�p�8q�t�hݰ3ג�ϷDe����zv�ʼ����6�=1G/��~@Q��ә�>�`���K�]�,�&!��T�m�:4FX��-/k筫j"
/:Wq������5y�$F,�x�YTQ�G�������=�XJ�r{�E����W�G@�'�N{WUK`�"!י]@��aȵPb�z�T)�w�Y�])�R�3�A���$�VJ�������8��=hm��SZ����<�Q�߫?�%�Ax��y*��twcft>^����X�S����݆��ƪ3=�!�Β���U��KSF[*cL5������O�ȝ1����3�n�A��A&�� �v�K])���	�]W�o]�[�lRP�M�{����y�Җ�Y?�_����jҋ6?�۷�j��Ѹ�j��ّ��:x/�?�}nƬ������r/�9�CwN]�����@�� �S�� (�V	�fg�k2�#݂J'l:<]�d{��l.Ӥ��]i�/r/7P~dTʊݮ�nZ2a6�v��*Ίe0����IX!,��+��h�s�NO�S��[��/��u�I�$�+o����&��Aqʒ�tvK�̎�sJe<o�������p35��v��i!�>��V�$�x�rʀukuy�� mﬦ��Y�X�������d�B�hbü/Sze��%#�䙕#-vZ�ƞ��[�X�����\�����L\d����/�,����L���eKƿՆ�1�w\��v��ai���bD��L��R�)D���������5� "�P�|�l��)^u8�6_�+�GP 2�>Y��!�G�;'�e��4�U�;&r�u/�C�q��4F��҉�x�n�xIy}Ю�S��	��+�=`���2�.�.���CTP�e�}�����?�u[K���a����ֶ��)�Z�-���O]��Sw����U��B\6�ƺB/7�N����)����mdrafS���D���!Λ��bw9��@wM{���wt�b[���k&긚��C�0⌧����*"�
��b�l�d�T��!g�����1Q�1ln� �z�H]l(2��8�J��|Z��i9lv,��H�p������H���v!�w~ �Z�S:\x���-���G�>�M_�q�Ã's�/�݀�MoH�#�G�b���C��;��8��êJ�=�`�A�:�q�V\
����{@�RA@��Ҙ,�1���MN+�Ln��ThB��Q��ж2L9R0��[�h�k���v9����9�;U;8����Ujߪ@P=�F���z)�"�BW�Y1Q3�fw����pZ��V �4d��
�n� 3A��H�ܙ��Se
���H������xo��7�`�����Q�?���_�G��R�r�h�u�m�ܝ;P�|��y��tQg��h&Ę�/L1o�������Ņn��l�6�z�7r�IQ6��n�J�5���'x���efX�b���nF��Z?���E�&��G?�w{:�nwQl3r�q���X�ZE�#������>C�Ք�h�NB����X9^X�`��LXfk��� g�S��h�+K�S����]{�#�&�وb�L���.ɇ�T`�e<�<�k6�H�~��H��p6<ݖ�^���|,�ϑFDr�������	d����A������O�)#@71k����Z-�n�Y��}��oz.!�	i����b'6���@8nHh�!�ح"���YWM�����ԣR���~�ѣ�ݾ�o�]�K��%���]�̓��q7�����5l���oz�B8�[�9ߍ�e.�^�}��3��9����lq"�?"'��d�\���IB����8��-XUs��3�P	������V\�vgN!20/8�Ƹ���l��\�4Z<�kft�!��K9vJ5��2�0/ i�>��1�%a��5;�Զ����]Q��s�����$��.������ī77.T��$2UMo���ǧ���Nϝ	=��f�d�G�.&�5$�� ][1�#���&��Dbϸ\Q��GC�P�Ǫ��$�n!�VjAn�]}�]���t�'7"�.P���d][u7�1' ���A�v��b���l&T�h�0d�Z�[��;pv#8RG�����2b��jcn=�I���a*�g����!�S�֏��L][�u7j=����VJ��T�`�٥U=&�>]�Z�c;D��h�ү����e ��Jt����9�Ftc��m��)��Ec�?��p��u4~]��WNc=r������"�I1�����ko��d�b�ʪ���cUN�4t"��\� rg�s 2,i��#��8 gҙ�_D`nq�	AY��]��aW�<hj�چqU]ZJC��ՒDZ��"UZ�s>tF�4�g�� u6b��n�g�q�K����ر������ 4/ߟRdg ͱ),��������!�H?�Y��dmQ���n��'�v�r/�[/�����~w�~#���`�rJ�\8:���	\\=�d_5�_�x���4��)���:�������$W��.�k�tY�R����M%�z��m���"�Ef�8��DOF&!��c��w�h��|���	����`����2�S��_5���q �ċ}���ϊ�0��28�$;� �=���/O)�$�zږF����ëV�������rh�a��}v2e�}@�4�kB���L
��5��-[�$K��!RB����G �Ca�� G)���]�l��4�Яp)��.
T�.���q�3t���{<�E#[-�Т@�f�6�ӗ��?���ɣ�� ό[׳T���-�G��s��t��[Z�)���`z܆h�9=Ӡ�h���IY�*G3��R��Gb��ȎƓ�!����Hg��+����u�$��j���í�~"G�� �K{���QgRH.[?ay�y*�)�uIv����V��Z��c8�6z��df���<z���Зl{���a�]#&�_z<�5!�#V� Kw��G?��e��~�lS&ě~��#ۢ�&`�� -/wC�̀X�^�U P@z�N���B�9	�{����y��^�6��4�?��<�,��8<��K�{&RZjad\�*N97}E����P�pҞR��T��bƴ��G ȅ�*���#�x(,:5R��9����mG�0����EI��؏�k��Wɪ^W��y�Z����QX����a���<�(1)��G+������JB�w1����6�m��9�R*�a�}�K��;��e��KU�Ƚ�ٺ�H*8��
�+ȿ��>�&��l-�vb	`2�����Ş�||��:R1�J�PQsB�J���]�d���Zʷ< ["��T��*d1��\F�K���C�
�f�!?�O��&���-�dh$`{�=:�h+�-��·��������k۬OfDm�j�mj۩�p���]2�2"��k�לV?%��E���r�
íl�a�ۊ��eq��È���H(LWVvi�W��+9ީEHo�	hY(�e�ǰ%�502w�m�<᎗�#n/$���>Ώ����/��a�4r���Z�n�Ҧ�QG�|cv_��yRʒ����AW�`R�ݍ�
Q�Xibl�Źf7o��r`�c�y���'�Pk'�O�W�<Ѕ[[���M��OGt�3떰b�ɾp�_����~%�Ž7�K��g�و!(/�$������8����)ɼ��@��.�؁�b\��7H��qu*E����~ޡ������6b0wœNԤ}��Q5"�#�K*�l���o{��cee�Kx�ꥠe���b�)8��<]E�(l����7�?���G[?�td��G\z����o�Z�JB���c9S	,��ቝ��6��~��J5Q��$�Z�>��y;8[sg�-(_ܲDo��M����A����ꭵLM);�tz�o5����-�<׹%��tS�������1f�(`���o����48`
�Cr'>$�eVk��$n;�mk���i�N�9�|6A��:�t4jn�+����ߏ�.p3O�򬿖�_���m��T�MpX.9S��Ŋ0cQ�@���w@jE�0i��31ߥ>;QeR�zU�k��<�_
�݌E:�c
"����}}��$��Y돑<�Ry�n��[�vU����
�(�G	wU;5.�D��	��@C�&=O38���X�VĦ]" l�S/|�k�x4£��9�5D�q�"�����֝t�D����)�-���r��ǳ��.�=���@� 7I�.?>"R�jM ?U&ܰ�́�/'v�ii��E	r��n|�*�ndu�U�ڱ���������
&�4��5�q���`�D��*=�pЧ8�e�rocGEyф�4H�|��9'I(ʨE��9P��'2����|;LN�X�!��&�:����E�w�'ʅN�|b�1V`�IE̙���ӳ~��l��%���T�usx�,�>9c4$��Sp��6�[?'h���O4����atM�;r�i�4��l=��:0�{#��c���ϟ>���*���.�? ���Kצmࠛ�k�R�vÚ$V[��>zJ�E<�BY9�B�����X�3�+��W�\5��C�D�#��K⹕2(fˠ�g��d�����
�.XN����G�r���{��h��X%h�|�k+k���L}��9)'YW���+B���)=^-(kz*�U�����g����T��DDN�&�����y�-�R�u��(���{Mŉ�:��`{��lD�#m���2=�o�a:�u)���d(n�H�����kZy��Y��͜`�e�o5dX�/�Tn^2�g�Z����z#$�����8�k��b$/��+��.3���W��[	����Y<��ҥ�4��0Wr^b�}H�xۋ$Ô
]�
��r�:L���Z���b|�&
䴟'���l���b�&W0$�I,殣k���d�w����c����+$��FI�i���TT�Q� ش,u��Cs�f��.]=H��"�յ|�9�h��i���O�t�z�%� ��éD9FD/���s�e�V1Y���(��L>�,����O�Mr�q�V���'��3�c��u�1��ꏟZV�� ���&�������W����e��ݗB�����YE+�B0�֢^`��r��k�{��<� jV�O4wʸ���em��榻|�C��2W��m��?��
(�s���'0#�3�q6Ke��D@����U3�NP-���3�:����f".�H�'L�9I�#B�>4�J��c2�w�^}����ƣ�ǻ�*ʓB���Y����5���S����<sb�~�^j�sih����,�]�V;�1�,`�\$叒�0ؗ2�sTKˤx�xojgRd<���EӘ��c��)ڲ�<�}� S���U])!�~M�W�Q(D������w�U)R-�k��6B��S�$�g�y*��d��Q���;�㦌qaR��A
K���?(ߪך��#f���=�	;�{\���D���ƈ�B(� t�4p8�����D����K�1�`����l�~�s2m,�.��K=!�l���!ҁR�ӝ��}�9���l��2��y�K����j�HCFl������E��=���[׾�!%C]�*jhIŜJmY��ۧE� �[vg7�@j`�]*}"����z�̈́��T��i&UT	�҆s���h�V^Ȱ�(C���`����c�t�Pò_�Ǩ�/��b��E��^�,��zg�ͭ�Pd�hzȅƌ�W��]���e�0_3�j�]�z��3bL�0v�xM(�p%<���D{g�AM�o'�acG~�sF�U�Tк��bi2�yM,G�^�(·!�1������}�������H(T���ד0��F����r囡,��.���σG�*C��m�v*�e�~'�W0����'�d8����]i����q��*٩v�	��R�]��{����p�fzs�moA�=�de)���,�c�AE�o�gLjef���s��nS����Zpf�|e��VL�'�������t�<=�w�6��(��C{�!�`��&bC��W)��٦S�������<?+#ʩ���5 ξ[`�l����<*�p�
ᬃ6
1�5�a@�
z�"@�o�,�Hٍ��d;�!��I�f�Y�6vu-ZE��}�ϲڋOo=��4�ӎ �)�v:5D��o]]�������{�����L^#o���r���������TqF*A��h�u���C�N[\q�?��G*�+�Y-��{���5��DRȟ�"0Q5��O� ��R"����D{$Y�����P^�s�� IX���zg�U?t,�ҽ�"�Џ���-p̷Lj���Pk��t��?�c��$L'����"�� �g}Ei
"BE-D照�z"ĕ�=�s��QHY�ZJx��D�EB3�*3�p��N	��S�c�b�K�G�'�^�96��e�|��p|<��ytO�̢�ۅ�Z�,��P_�p�)g�ч�v��pكu�Pf� �����<���Rhl�0�\<߬`�o=G�4�0����E�յ�������kk����k���u5������g�+@�<U�����r�[ӣ̿LE�ڢ5�	��7���C�_�P	���b2mj�O,uNW��߫��8恭� S�AƗ���Xmi��]`����F�Q6�gG���5�����=�� ��u`�3'�����fv��������,y�MiIO�:n�V���'/A�M����+��'����]$ h�'mc\�/�	��1��1��x�j��:�X!�y�_�n��%2��kҫRu�afq1�g������O�/�J�N�x���e
�֕�'��i�]3�M�R|�ٌ�!���q����0�]/M���2���]��ݷA���K�D����E�:��շ�`�P0	�ȹ���5%;.�s}��`jxN�{�x�"����g(L�8��f�K�cV�G�;w�I�<�a�D�)�0��C�lw�S�ul���mCci��wB`a��y�ٵy�!�g˥3�t����"WF�c����Q�	{�w� i�R�gV�\ܖ����ˑ��?	n�SZ�M�)��;�1���7d�w���댠T�8�#��S��-��`��Pz�����Bͤ�����Q�`����9���wc�H*t����u��N�׀oU��w��ʥ��pHECB��&q�d�.$,�P8����m�"9�j�YIP��@g�[[��td�(��g�52��cṆo�/��$�+������r�ه�DV�3���&eȠ�%W.�ud	x��^f�m�"
h�|�P�@=��g7C [3�!�éKxWP�I�HrR�6�" �[�*�j�=�̑d�Jy���cc��%�C��jJڤ�X�^��=*��_N��z��D�HQ_��=��ak>�G6�
6I�bZ�3A�y��9����q��E9���H��?�.mrǃ�2��.�dˆ��蟍1��>���Y*^�d[2�7�� 8��׃�Y�\��NS`,�;�@u?�����*�g�t�g�ё�.-�E�������)��8h�h�H�n�)o���#�}("�a��y���n��1���B���?�E�F���W�fJ:RW<"��D_P�>��ۛ����Г��97�_���]嫲t��$���6�����̉�N� EK�ŵ�i�<hXl	VK�a�����h�Qց�¸�]xoS���]A�����?H�8���~'Pf�{�-�;~>�;�   �?$��x�������e�H��g;ei��~������4��U�wf���W�[�߹��x�oA���e�G���
�~1�r�I�������J�4w�0$��@9�9�W�c#�1��`5eO��Nt��3@�i�5
�u���,$�rB��ؗԍ'������as �mF�׺�l�/�e��).́�}AkX�N�å��҈�0�����-i��3�.7L�dF ��s53��s���V�E�&��i�&����*k3�~@Z@+=��gw9��bjpِ)���;��n��C��� !�p�-h����Db�+�����6\!�Gr���Hbc/^4D��m����Pp[)��@��
�V�i�bP����7weq���a:w}�K�n��"}q�q�G�&�86Ϟ�ߥp�H,�ې�0O��^ �A�)!��`����˗��ixU��<�c�{�d=�H�oF�e*�\'���9�D9>;|�ws����LD��3а+w���.�x��,U����"$���2Lc.�c�:�$%Fu4�2k���Ǣ���oH(��u�E������A���qI�jY��`�.��i�k ��6�MtlD��y��U�,�`'�x?�wXo�9�N��>X@I'�$Յnda�Lt��/l�@����X�Z�S��~�"��po� <K��_��H���=NJ��!�Ukn�9�'� ZC��}�M�̏��3밎��3Z�a^}�ObT DrI�����zw�����̆H�3�f4�ZoiS\�PU|1��>�y7q�w�}���1x堰�A��Yzo�0һd�p�c(��f��^@�7���9�<�F�?1垮|7��<]�dD��9�#~(��M�/�P�h&�5���/z����i9�C��UOC]/��㔞]A�@��BP����8ۉ&�Y�q\�Ѧ�h9F�q�lg�ڴ��'�W��4����x�Qv}0�sY�F[Dk}�z��� �V��d�A�ם��ے�C>u�ب���n�I��0F|�}u�m�9���u)��=�L��n�����r�-u�����׍n��g��D���m��^���>����t����D��m"|��i���L�K�.�jO� ���@6���Kҧ*��r������oz�7�v�{������#��vqΝ�T%c�@*��w�bEײ�`G~�:�1M+�ې�1�]��p�,���/{��~��pKM`š�,L\I��X�����:	L��䥳R�? Qx��ѵ�)^4��[�>u�����!�v���1� ⁌a�f22W���0������!;6�k�yLA�r������RcSW�9�4f>�hhl�DW���
-<�<1\�:�D2�&�o���T
�f�:�<�[7~�z����&��lU�d��E��J9�7�s�SY!��`�{�N�j�.��j*c��H�m�w:d�
-i�{�#�
m�ץ�St0m�t3j���İ�Ҍ96�Č�!�Dr���H7�)�����L�����.�ð�=��'��a�=ײ<'�����J�\��=в�*K.$mb�J1�,x˺Oɸ�1���of�A
��P���6��Yc�AGQ�6$#%������m&�Ȕc�cL>�q	����4"3qTF�P:Q��U�l�f��Pby9���H��+��?�UK|o�3�&���(P�
��/k9����|����N���f3h��l Ţ���X�AnՎp��#�;>��ۨ[�t�Zl�����m�1��g'�K���b�l��D%�gU#��ɯ.����;����.�*O@�=GW2�f�U�R��#F�bu�&䠰�o��F{��В��m�FH�BH�N3���R1��aᅪ��%6�R�:�o��l���.ܑ!s�9z Й����@Ua2#�#u���5<�(�ĥ�I�Կ*��t���Ә�ɺ=,����{��R$�EY$5�K6�w��`B����g�KyQ3�&�[.�ۃ}����A�9s�޲��|9{i5i3�>h͏�n��aY�	f�� ��������)�	9���*���:P����e�/��n���{�p{�4xY�@�I��ֈ�<�YȽ���CW����v&H�c�9�!(�W�Q �V� �la�:�X�A�j�rfpP��R���9�"~�[jR�n���{��@��!>t�""AJIJ�{uQn�%��Y-%�7��Ðļ߰84�%�<��3U���p]|k����`�XE��}����>�6������9|c�`-��0�0���WQ30nK�"����b!�ϻ��;�L���EJ߽���$?O��o��ԼU�C�b���oU�P×�/�Mӹ�jg[����@���*?u������� ��<eA!u9��:�*���;�u��̽�H&�Յ/�U,�4zE��DFqb)2�.�E��ڵE�sʾ�}r6��6�X@Z��%����2��"�W�sRr��؅�'Mv�QM��TH�ǔAÁ"lG�Ҿ�p�2����Y2sTE�Pۋ�L���	
�r�]O��������x�V5����~�>��!��)5��r��L;�^FY�w��9�ޟ�h?z��q ���$�T2�%i>�q�`mw��������@��Fe�Ҵ�|]#�<�\웻T���!�%U��_��f��슃[�`�u�E�	�$da�����d��t����3�L�L_�����;��N� Wq5�?���>�c�;���� �
Yݎy��ӊ���2�h1CU�埪�aT���-�\H"�����`vtkE��ŀ�;"7�D�R�%�Ŝ"�R�%�,����D�"!�Js�Q:���O;���]u�s�J|tUs���W�e��P0����Ӆ�M;��J����o�=O���B�)r ��d�b�
#�]�4)����y6>�[3�ۻ���Z<ڣV�u�����sկ��EaG"��VX���v�~�P�5e�Mök�oE'�7W|������Z����+]�E�� d�:z���d�8�N���1{2o&K���u��҈�����-� �y�hO/i%wء���:�+�[�%*ǐ2�]�7[�T�/��q�V�I~��y{	�5��G�NjL¢�9�D%�g��2����:�#$���~y۵�\���ܘ��+״]PJ��Q0�������$7��?�����R�_Էn-�!��6�&q�Ė��C�뒏Yq
��"|j�(Ն��F|A��ge�x�Zb;Z�o��{��K_�F2��m�w�R�#� X
��~d�G�����Ly��p��W=��!�ڑ�K&�������n�[��j�zO$�	s�N��~���]�z^�O��*��"<���a�4�cD�@�kO�a�ĆZ ���{ b6_qi� 6z4�9 �D��rU�}M���3c�d��M������7Xf{�iţ��1@���w�9|�N��Z��F���2��� 2��)�� ƛ1*���0uI�+0��o�>$>�~޴�P�R���2�^�a4�!T08����e��>ǠRè�F�f&����RY4)H�?0�k�RD����T�NUH�!��Fǉ��g n�ީE|Qt����˱0+�����X����'�F+��!6pt
�L]�dL��_. p��&~����A�I��N;�Ey3����yb�2�j��_i�����L�\�
�U��JE�����]R=;�م���V�����-3 +%c72DX�����򨀫s�5~�2���/i�h�o�f�ad_��Ek�e�ț@UaUT�R�D�RYu���.3:I#"���a�P��_Y���ڶ,y0�\���r*B�܏2>���a��$�ޟ���(��,�����2�lnxÆ]�ь.�)f{(/��7ٱ88f�����K��"]Ӻ�mm����v�I|ǁ�M!��ŰrK�#�h�~��kԿ��̨(�����q_.A`MA,��5�;6K
��>�j���2�.�~���N�Bڼ�u�'<�C��#km�4�����a�#. �2�̧�ι�< �>����{��p�A����e>��)t �(\x�0�扉�<�	�3K�Rq�{��vB���r����C����]+�\�b�]t7m��s���U���>J^C�[�YO�H��L��5;�-'����'�����������]�~k�I_�:�f�+b��_����"����|eH�m;z�&�U^�(x���NzC�?�(u���u�ob���B�_�'H>XQd(�<���㢚����(�ڢ#��[�{#���Χ�h�q�wam�J<CA��.��X|���B�ƳPx�k�
�np3��ϠD<����/(��9,�����Y&�Cp���)�6c��;vbf^��xW�uGd��C�����t@A�hY��.�KT��y�̤����
����5?mە��YeTgr��`�)&q8�h�u��C�O�ޗ&���/$[&_b𦽐��40�2D* ��uG�[;�t1�~�tOc�a���y/'������F�ň�~�ޥ�'۲875����1�§��qW6w6�����$A�Ñ5x6ktMI��
��f�9z]�il���O���|	&A�j�S��(^��br�����_2�D�BL���e��~�'_�Ej64:���HNt'ب��,�ټ��������5^3G��~!<����o�{��q�	VR�a�g=ٯA�TF�e:�~�+��:��Y����7��>���U���*���9n�	�����д;��LPْ��Ո�v�x������w4����B�pR�ONn{WA�%�M�*�4\R*�S��!��Au�}����q~v�;��x`Rj}ىc��҄�@���q������x3`XBw
e��G+3?���*_�[謣�畃'\˻O�)�v���[���L���/K��\���2i�����K<P�%q\����-��C	1���j_���O���&��MW�O��z=���?E��X��U����M���>Z/��;ղg>,�yUr�亹!$��D8.qI�l��2}�$��!�K�c(��d�aUʎ��r�`�����,���itV����O:E���2tP�K��e�GB�����S�i��֝a	ڀ=N�����{
3��D�r�n\-�����-���Ι�S���3�MH��2D�I�#lO�XlQ�a�e�_����Ym��I��Ł�{\ae������q9h��%��Y�Oq�⚋��h��Mw2����8�V��m�Iq������y<X��qÛ#d�-���2f�+�C%�XX;�ک~���b�zd�9���ʝ�^ �b�<8+�_���D!C..��۝O�`7	P�WD�1�I�W9M�� İ�%��go�:�dB�M�$��*f��v=dW��Z�飝���F-Kw�,�t�A-~��1���}�-���Ɤ���IT���$��1Sk�{���9�.��e�eG@A,�6�Bn͖o��W:e�T�,+�m�ש�G}��c�4-q��Q0w�s������FZ2��K�Y�V��і}�27j��r���I�����gՠw��ן����ߖn/��"��O�m��L9&����Գf�=A�Ѡ���~ILKa`�ahK>]::��rGV/e�:c?�ȃ�>�{�}v�΍A��ASqa�q�#�^�OTSB]W�oM%0��Ҕ�=�ٵ#Y�h���<|F�_`5Ɉ�p8�A���"p=;�z:���B��|�V &SG`"� Ǡ�X�ߏ���:�Z1�B-�H��Տ���W
"�hs�$r��j��34g�L�b�YY���Ne�Z:����S&Ikc�JmH��U�aΐ8�
��"M��ʨ]I~Q�{�tA	��ښ\�t�f�FA@�G���%�f�F64�
��7�L��dl8�X����i�	Ĩ�6�b@�z;��Y��� �
z�͹�[؀j�w8��qZ��#����X�խ�=���
ek,Y@�<=7�����W^�nV���pG���F�g�۶�s��<�>��YI�Z��Dn���ٝiy�B0qn��w������A4YN�/�N�������Ǫ���q&ĩ\f#�=�P.�a x��oG�#m*�^oQo �*Et�W�J�`���g��o�0���H���**�G_�t�(�X���p�Lq9d嗕"�Gd��p�����d�/G�;�n����l
��*e�WQS�����x���ԥkLw<��.ٟ
�A�)��9ZR�M�Y��}�A����Tݮ/��tm(g�;��y�Bs���߄��h�5���R>S��M{��˳U�K�I*T�OD��m�u��)t�,ι*-�Y��#;��2��d�&�*t�{IT�7��,�ǯ�&�&�bb}�0�S���H�O��TKY�y�~Z�#r��u/�px3���SID���-�����n�)�J��m69)��l�֐�@ܾ+�Cs,���{� �vT� @e�B��k�NNʖ]HY� �6J!���'@Q�A�#���7�j�椂ޭ���ʀ
F�7�����BX]V8��"P�b���:�/Ӳ�4?l�0��B6��]
ٗ>c]0��#�"�4YB��q.����d ����V���$�,%̈�\i��[3Rݪ{�.�\?�½��0>��������(����7Z'_�w���ˊ�-dˏֻG'� Px%�}��Mk�^�_*8N�><��{�`v�U�M�fkq����w�,�̂}&�/�*Eˠo�-A�0��o:���B��Ӟ��C��IE�c�>���T��O-5��D!�K"�bVii$-Ƚ�`J��T{"h���u�������X��de��W������Ն��*t���^�=Ǉ�G�dg���-�~jg|J0vɩ'j�D˾��ض�� �yj}O&��`��Y�?�fj�Uf^�!2�YQ��u�:m��T��5y���:����!�7+���Qg�r��c�G�(JYۜ������&ʝTx�>����3|P��w?���q!�$�T��N�O�B�J�?��sƽ���A���`���3�3��t�
/�coJ�ǯ�|e��w,;c<H����<{�ͦ&�J-�dT�$?�J�Y�_ϲ�So�v����Cs�b�xJ�1*O��^�1��3�{��6̜@�ݯ�/�EP�t� r� I�̋;R�DT^ULt�pZU�g4X <k�k]ׂ���C�a�> K�����.���@��,"WD��4�P���d�] |�oi�)|)ύ=Ӗ�ea����%�s|� � �9)W+�w���ђ��+&�/l�{�Z?I�s�o:w'�M2k׻�F9p�� ��$�T���e���sޯ����bw@�� ��j���*B|�@�5|}��9�<��~������51��(C����!C2B�cIIZ���7�B�p��*$)���0�e���s�Ó4Q63�bz�Y�f�����2ְշ���k�{���&9�JSp���A�\���6�pJ:�$�i�O��U:����RKc^�s��Ic��L�?�C�7i�����{T��
��{N�ZӼɗd���A�\�v�	����@+gƹ�A�.�VPr�D���hvۘ,Ws����ߦ=79�#�[z^���{�9�(�S�0[��2n1��`��8_U�Dqko��wD^�y�C�F�aȂ/2rL*�Y�B�1~����7�I�]ܑ[��"[}<'�M|F��֮��>�I��_pW/���q��������Ђ]�#�����ANtu�Nf7�����ʳ:) 	�p"�i'�$+̒v�:H�H�!��R���ޒ��p�i��!Iֺ�9�jT_x ���BZ ��~�A�fr+�G���Q��q�Pt�<H�E���:���(��S��^ueۅ����詃�M-��;qA��������K�)�ˬ��x�9։L�߽�Cږ������剳�I�$J�T����9(��CE��y�<�r������s�g��{p�LOD��³���to�:�!k�����j�
¢	� ����a�T���
���Eb�##9��ד��-���'�_tJ��䜢"�ew;h�B�(סDf5E�(���`���Z�P�X_�#��9ưd�;�L|�go�{/�����_�k`]D�
 b&��V���;�~QaҞ����5h>(L�A��\����-�TG,�a1�i�^7��,��ێE ��議�FǆNƂ�N�W�?�X�#[��\.���㫞h��Lz��C�$�n�Yɷ�N�A1��}�ó��8�HR+�[��c��e�3k����P�{9>�|6��Z��nM��c �Wñ�c6�x�톉	u=�r��xP�b<�y9S �3��$邥閱,� ���!�=�� V�u����I���]��``�%���Z�)�������|m��m�qS����n��z����đ��	����r��Up��oS�6"zJ.����C,<tX�@{5i�]�Ш1�-���s��d�]Al��m-)�����;&}��x��0E;ɕGn4ph���;{�_��~=���p��5JHg�0mk7x���h�o��`$ԲS{�~����v�;T�N�K�ܠ���|刓x�<Q`2�ߖ��9/�2�:V�~Xr��*�8��򋚗�̆.��~�B>�X�{�o�g�S�>�k�0���M`�\R�g`��D�g�W���sT�ڏ����;p_a ����K���u�{�1�jO�CϨ���mjB�6���+;�L����ma����KrZ��{ �+�ǀ���@��K̶p������\��8��:�|�>Iig� Su�֢
�u{��p����<3N4�,��R6�EJyV�ٔ������	��d@�U�"��"��6G����N=�i]�B�J�m+��V�����a���-@5K�:w텣��A	K��Tr������\��7�P/�1��!�&���/���̎�N�*�C5a�F�Ƅ�"ɏ�i�n}� ���`�8���Y���]���h��*41aKT=y���ocI��^�<�$��|�ꛠVgMw���l8n�ƞp��ϙ߫� �'�ΛdC�������FJ1�8Eׂ^�5е�%q��Cߛ�d�T��|��K�w�o���Q����QA���3��|xo�e�D��K]�Z�ٿ���@\���z�r�
� �ˤo}9��6wA�ɷq�x��F7d�*��P옶R������PG:wxB�,@	(M��wQE)�[�)������Y46r��R�^��`d���C�Z�Il���]�t@Q��������%qW�2����,���T�C]}�K��^����=lfl��
��b�(�gX&86V�31��/)�*b�||�X�x�|�;ࢿ \Y�ˑ<�}��R���2"���(b� o=bf����q���p��}�
ʣprR�f�\ ,C�v���8��9��_��N�*�\���o^NK�n���V܍�K3l���L�կ==�A~lyi���OS�	���0{_S�/w��i1wb[9N�q/��ު[{(,Y���*�3���)f�_����m?>[*s#�9:��/���e{q}��P'>��A��DY���3T�9���t͢C��k:��B�� ����s�yR(���wm�<~�����|CʫCXQ����	��5w�1a�"o�4��:&�7<�%���o�tH���J'��}�舥I��Nw%��vh��*p���D���$�cq�\�e?M;Wwb�ʹ��'�@
��7���)j/Bf����w�U^�X���A� 5n?����6�p���Ȇ�����b=}�.��c��B�ݘ�#����j+v�<7���P��|ULJ���� P�`c����o���C�����+EB_�]�5|=�3r��*�x�W���l��{�r�Z�}��0ИA$��x�_�?�� G������#��5's��7&g\�yx��|���|D?.�Bώ(�p!��1��'�-i�o}Y�����?
HBa0o���ߦ�I:�ם���z3
�l<��ps��I��X ��E{�IM�r]���ΪT�NX$���O��I�ed+՝BS�O�z��}�c{4�s���4l��A��S�Z���9u<�X"7*�!J��+{�������F�FAυ�]6��h�n��Y���4
^��m�k�3:�G��N�0|��
')�@�.}ձ4`�9r�H���H�Y����H_*B�bpHf0�/��x?�����!	C��Tߡ�J��AsaW�_�Z&qq	�u��p��UAҊ*�֋Tc�t��I�E۽r���e�uyf�1/a���W�|��.��3xWԖ� ���@CK��%���ٷ�K%bhZ>�>��Y��>��\�<i�j<v����a���b�
p���? T���$n���=���f��lD*�,y�Z��KE��A^ ��"����x�w�d#M� Z��U ��&��n*+�>`�+g�p�+($��F������su��(U��f[q8����e��O�M�t�D�s�7�dlA�j�1��XZ��9�נ�#?���>������,G ��U��.�����sA�PD�A���N}���3�;�qڽ4BY�i�w+��,��yn���R���P���>W�5_�?��8 lʅ�A�w��,U��e�p�yRxK�GQ#؂�����2��oeZ�2{x������;���t�6F����wr���s�F1D�s�~��]"v1[�=�M��q�5���a�	���IJs~y$LK��w/X�9eK�n�(L�a??g�ČK���!en�\	��h�&}a�����)�n�
+�=]=Y�x�bl��y њC�lX�z{`x	�����:��yz,��A&�y�W{�������wݶ�?ɯ&i�SNf�A@�j�x���Q���!0�9_]E��[v�+X����TWW� ���q`� ӦO�3�I����f�$CH���FT\�+���hI��`�4,ɋ�s���S���LfNA��	�gLG8[���/���g�����B�S����+;`Y4 MIiuz��^�b.��RuFsr�Z��֚Е�.�QU��;5ŕʢ�C�tL��C�!M�����3��>z>@�6 T������~��eb(�����3�PH�瑠Ņ�I�h���qQܰ�T1l����j^�>!�B�:��F��A,�މ��G-Ӱ痫�D��������5s�J��noy	؊��Cf�����d�7�y��qș����*�>3W�sň.�!<�D� ���G��{t�Ԕ��p$>�+>xMe��PK!)1W�����Nۀ�M�6� �h��5�<���\��Wx�@^+I;��e{��C3��@���B�[V T�����S�1��}���R��ɓY���(^`�A��T_5E(�� kr�Y?��ߖ��0��d�?xX�o�D^m�g�8!�\����'+a�h;Z���#T���e[�|��Ғ�+"K�j�LC�bP�4�\x��6�lF���$(r�7{�̐�P����$_��Y��E��g2�z @FP>�s+�=���PJ��V��$���du�*Y9��Cs@��1~*����gN��O9��`N
��Q8�q"�E��/zJ���j�B���nj��H�pq'��pt��/��3n��'q� ��a _D����D�ݜ$�	�5�~���i�t�pk�a�a�*r��w)G���`rr]��a�'B��hC ���eިR.�#�����ƻU����Z]Q��<���:nn+�Y�n�d��8dH��f�5y� ����*DG�),�h�&%e ���c�b_���/��=���]Ƙ���6�@��;g��T;@�V�x�O�XA���~�5p̗��3�8�}pyp�#�Y��&�s���Nʱչ��:� 2��i��Bg��t3[�����Ӌ=i?W�$�&z�B�dF��%��M_���iޠ���� ��-���: ��o-