��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P��v�"<ߞ��&'��k%P碶�R�ӣ�sĞ������FY&�~l&	'��O7�A�c��|�.��d��Uڬl���ʚ�������5B�x�,���5-�ܷ,������� g�r���œ\:s6�u�-��?s�Z�� �[T�������aC����Y�L������f�P��ǦY�PX���K�B����dى�GK�c퇬��9��U�\$�g��q���!�f��08<���9���hh=fY�3jx%Z`#����|�V�L��6��u�Gp��pV��pqB��3��Q�����<j�2���#ܭD�����ׂ��M6��-�Ʊ�}�#�x&�*>SK��B��������V��N3�l�29�|?#�<���;�ᔡ�В��Pث�9��ej���M�����֤k�\UU����i+~m� MF~�7B�"��tT��d%/S�.M��iy��8�;��~@���K����̊�e0iȸ˵���?7�o�Mj3ۊ��B�yH��*C�yȍ�^��s�	�3]��T�BxީV� ��҅N[@�̑���%��& B�;�k}I�P��Nt�{��\'�N0��XH�O�BU��[o�C�I�w�}�p���P0���ϛq�k!��o�Z�#KNӤn*:�{��IZy!���ݼ�G�k'G� jͩ`�r�x��7�MG!aʈ�^=o#'������^��]OH����[�Ś;��m���8%,���ۇNe�I'�����f�b�pށ����kT��Sm��|��ږe�惩ҴU�2�
{M�k��?��u� 3�A>�~�Y\5ꍭ ����������&�4*>�	�wG�1:}�Q��U��u!X_�>TK�;"�f�yM����J��@��$yM~bҮ�fz4���C��x�-�}� �r�Jo���/��,�ƨ*�U�h(�*h���.���R��H�����K.k�
ۡkg�L��^h,պwY��|�I��S��L�F��gb�y������.��V�s�_��
%6�o�xd6i!�n�~��{��.]7%6_��6�Ǳu�$*b�����å:(y۷�M՚�3/���,a��~�yv~���5��H�Hհ)�*�jS�ʿ7_�x�~��j䊉E�+�'�n7��h_��+@=K����+��cү<iA����ѫ�4�ؚ]��l�a���=��g�M~@���:	n{���_�3�w��P����zP)\���6�-qW ��)��DI+yѶ���R�/��l��o��F�4IxA����舲[}�SD�},��xGva��3B�V$:q�3�D�Ըb�e}A
����H��+P�����d]�&��cQ1ϐ�b��y��U2`M^�sҫ���Y7�*x���͈�!��'�ufAv!�C��J�cL�V���Y�q�0��)�
N.�L��w���N�����<�ȹ0��.���(��X�jB�v{��K�)�Q|�n���.����c�Է�'y�H��w��\�\�W�5���tB�G�<1
Xm��P��� cVXb'ћ>t��>�f��'�5�Ӡ��>�H.6�P�5��ǵ�ٺ��C9İ臆a����!�ܨ���^\���}c��rwf�wǽv�[F�G<'�e��ir}�f�����6U���?��Ɉꄕ�����P�����z�+������s����kQ1T�]��P�*��uK�.P�
�f���im#��0��(�L�~���)=.���P����ɵ�u'G`|&�*c�"m�1���co�	uf_�9�y�L�d�}<d#1"g=�CXD��2.�+lQK`y�\�l�L�,�cF�hd�d��u�I�K�fV����!"m�kr�T?��_������:-="��O��5�d��-�m���+�U��y��p����2�@��ֳ�3m�s�:{�p�N5�h*6TQ���2 ����\��2HگO�aa �� J?3D˗���Oz�N%���-�R�Y&�$��aD�og҃Z�h��Q[4��P�T�~�T&%סO����$5SJ�u�:�S�)�x�hp8�P96I"��y{f�Bv(��"Eِ�N� � fI�nG��]�G��O�K��R��z�O�QV��n��F�jz 8~l_�}�:���k����C��&--�C�M������N�Tfx���u��`k��D��'p8�ш����&b����t|1������d�lIS�FVӍqA%��l��<*˦蒵ؼ�!,�����&-�D�̍�����Mq����x3�Kl���m�h#9��b���� `��V^�4��	6�%�p���#.�)��[?��Y��2غȐ=x�D.�U��x��%�a��8�#֏����Ei�%�ӑM�J�~u$�8̚t���x�,����#��Q�Qʫ�@}F�<Ao%T�
w-3��.�ܛ*��2�QD�����ը�2���:���&MJ�mL&�0��#rT��¾u��JRXs� ��E��s�Q�Gq��v�L=����9�����Q�?��D#�c������4���V��������J8�ݶ;��6������ İy��PtP�� �.�ZɎŖ�"#�G���]�q��S�jβ~�����A(�w39}�փ4ǴΞ��n4�VL��=R����db�Ż�ZV��?]L;��/l�P����M�2v��c=�� �)�Y�x|`�� �,J
�'8r�K�T����Xyz	��W�¥��C�Ϥ������
#��4��/譐��ð
���?[�G(P��:��_�/�	^ }�� `�}�D{���?�����2kV˞����Y���z�K(�D^CpW�}��0�S?f#�Pfn�l�����V5��ڎR�7����f��R�xX;h@�4��c��A'(��zqs�/)5ÉƷ��j��4'�v�5j�bs�㕰�z�N ��-�d��8E;~^;��<G���[������Ok�� ��(��N5>�
6����@���I_>2��ɿ0N�XϞ��_/��Z�.�)�GV�_>�q�.�g3$BA��:���������_��ɏ�f����r@4$� ��ӎS"��֑�O���ku�B����g�s��=�qg���%��]LΞd�?��h~�w\��+��ѹ������hqB5ޥڷ�n�B��8��}����e=p�	�%�;��x��y0����;K6��Û�-��?!o�,��q��R}�R�w$T6��h����ȉ]���`�ޒ������{�����ǿ"ז�l y�⹵����޴հo3[�%������!6�9r�&�U�9�}P�8����g ��z��W���܏��/!��hF�j.�IE�~%6��l��7��rN�}��D�.k��{,�z�,!���3#�E0��WF���� 8��Ԧ�|���j��n�1PܔTog�<�Ýw�����E%�)����	@&C���霑eF��mk$�ہ���̝$m����I%m�u�{���� ���,WU�oB#]��':@�\	��혪]���%乿�i�y�����mu�t�L'o�Vh���H�r�#�����r�5�"�Q"��</��	,�-�ׇ<�q�6�Åv�4�UI���IlV�7(hA�Ž	�������FP���M�Գ�Z���JC�L�܋�v��zT�Ђfc&�MSNT��'��|H�ɝ�i �E?����0x��CMˌ�L�}���z����?��$&3��C��;4,T�%��Q����l)
�@�-�Z�օ,�e*�]��\�+9xb��J9�i6-��9$-Y2���^�w�j���e���#����+:��9M���E�{�wh�fR��,�N Q���֌tG8% ��K�J��sF��YId;���+�-���.�`��K�m�j��KRY��^H�A�E�ba`(�Y�t���^�2����2WF�;qF%d��Y}���@��rI�F�	���(���-+����ȝ���"�o�Y�G��@�$�+���Jc;��lO�jk��hl�Jc�F�bM�=`(~���f,��4eD���V&�� ��-�&�'W�76�)|��zױ&BC��k �]����K�-���&ɴ;�D���t��(8~�\�XQW2��}� u*�O��M3M�W�V�֭�H3�GT�����q��46��en�{�ep�T��#ZW����!� (} ���!�Ob�4b�XrDkG��d-5�c� �#b'EԂF�VH��;���Yk����U���f"����6������b"-Ѭ�R�3�
	[�@�>1�2lV��$�V��/+��<@&�VW���Kv��Y��,����WԘ���#�xr��$��T�Q@��b�VF���^�ߌ��|�N�p!8h��O����pꛊ㇓3�Q�]pC�ѻ����T�Gk�(�av�+�L/��i��oP�׉o���Sͨ%�ޡg�iWڻ�uM�J~9?T�[잊�>��Y�&)Zہٵ����}�+����p�5ۿ�Il�<�%����|�vɛ�d��6��/ad��Z���?rL�+�/�b+HI+*��nE{��R�N ,u�LDu�Ha=�I�PtN����P)�TO�Bv���pl��
�9M�|&@O���$f��Ձyl�C�T��pjH��خW
l㍄�./Ƽo6�K�o:"�9��Ėy�z;�|��f8�PI?q��� �x�$�Q�S���{	JH^�%���B��<�Ɲ�Yh�hݷ��/�`�$�7`t��Z�\2��ة��3�
��z�9[@)��������CH��F�y��p��[eǠQ ���ܵP��i��>�MN i�^�!q/H�T�[C ������>��d{��Q��ŗ$�4"��;5|��d�0X^�����۱�����(�ڠ�Q�.���ne�\��A&'����F ���;�4/-mUܩ���Kk���r{n��r;
�t=�����\��Gd��m ݬ�����-~co�La���Ɔ��g�O��IPM]��vk�@a�? ����j\ �0�y�|Rۂ���cJ����{^[vk
�Z���LO-��|n�(�re�>� ĕ��>>�<�F��\M�_@ �"��龜�<�7vy�'����x�?�����@}��]}�� {�ՌҶpr�䮩����w��!��\�r�=�%w6���V���zĽ)k��ӎ;�.2$����`
[�D���-d|������`;�Y���E�<9��=����^�|$6��?0�T?�ppS�ϛ=�l�ի�]��O�(����u	��AU��-p����&��tK��*.<W���DngNY�$��-[r�ů����)d��ܷ8���e1t��H�U6�⤵��3к =� �[Xڍ��%�rZg�\��v���Vd^UW[M-��XK���@���~<��ٞQt
x����n=��\�����mj�E��Zs��U�*_�7�f�Mq��B�|n�#���}S�.�$��ZƩۮP8�~��>H�{B�\kc�-���r_��`ܨ32_G��x�Ǎ\m)τ����5Iehx�hkA;Y�����v�,Q�:��D흀�U
͡�FF�4)���z�U$;h��s	wr���+����ׂm9��;_�����������%@.�tg�7b�6�J�9`G]�!���Z�*�Zm�{G�D��G@�w��z��[w8��Q��@�sl3��Y!��Z�+r�:	���H,q5`M��	ɸ���jZ7� m�59��k�jː�#p�w�KUJ�]�3%.X�K
��Lz����=ջHl�)Tճ���@1�q�N�Q0����SR�>bu,�ʋx6��	�����n5�4�y��m�$�8��c �Xp.VK���թ��%*�+��z�T�k�L�-��G�:����L9�u�C�����ZUG��L�Px}BK�E}<d
�B�*\��L����K^���K�_�,���]��1�|Y�~{�}-^,�O�ެS��.Sx��>X�Nr�Z�N��3p�_��������P��t��u���CLL(`O�m��]oV7Z�M��:؍�^ظ�R(p�&�[*E���2��G�lC�Y@��y.חMlۜ�䲻KyC׼��"OR��5C"��1�����ȪߖC�0� #�$�.g��Ǚ4}ڋ�ݻOt��p��}��%|R��Z�e������H,{j���
��ҿ����F[��O��3*�_F��C6o�ͺؐ����k�7C�����{�4��ڥ�p5؆�\�%Q�+w�g�\�D�/��`��橨o�DF'�E<1�O�W� ���*Y+�rbٖhs!��C��1k�W �;cm>�c#�� N�:�μ��8E ��lW1KQ,�=���6b�Gi+��[_(��|�0`���D������=$΂�ƲPx���4L�}���ȏό�?b$�*y��k�$���fb2���^����׾54S��~"<���x6�����ws��N��ik��3��9*b��շ���8G�9��ìd�Q�g4lRv�H�` ��J�
�"���1���.��4������
O�����Ix���9�j��6 d��>&ף��rb�C�'@U�Y�Ǜz���c��E�����F���2����m�D  ��̃��b҄,;�sl'(�I�w��e�-�@@���Pjy
%���ADk<i3����C�{�YZ��+b�߉����Imt$��AgZ,P��?Ev�9Ƨ�ήa�f�`2D/L���7HN���?/�KC0&ݓv����
y�:��G�D��7w?�I[�nDn�����͊�H�͂>�e�l�\�q����ɲW
�����>��Z�� Ԅ��9��}��0[��V�j?��Ʃ���ɐ��*�/O^�DZΉ8b�^T�$��/���Ui�}V[vg'�hi��[EȎ�
j\e#��B)�i�q������l�����WA���?eo�G��
Qå�=�'���㝕��u�on�*Tz��R0ա�E��F��v��mKxO(�\,��a�@�-Y���-�8�b
_[&��-62�!\�����TBA��c�q]XTVd�D���U�#LI�4�R+#xY	mb`_�2ᆂ� v���"Y������_��E��wA��E���(��ʀ��m	�eVW(�˪�xroi���6���� ��/]�.���Q��Gc�2��.��TD�σ($�s���z�T�׸�R�6�S�)&8޽0XR��h{1�b�vДkF��6���0瞍2���./s'���"��`���~,6�2�<�+�MF����H�i������k!�� �EQ�Dv{�Ӥ`\*�	-A?��B=�6���Ѡ
A�26�U�6ݪ�)~����V��F`�L2�X��ز���b
�%y5u���dZ(u��u�Q1}sV�a �����c��KY�+�3�Y��sw��*�NȻ��++�� �K/j��9��|���Qr��f�����l��.~�>F�SgT���/�!0�{"��
YV#ϙ�p�#_�F��$�_��e�%����ӻ�ڃG���"���6Ő��֑�&�Ks������PP�ؿv;^�e�ǏW��ɞ��Xbl'u���H ��i�"��.}
�Ÿ�l�^��c�Mj�<�P������\.N��ф�z\�N���a�2�&�F�����# �(x�.L�66��?��=���R�5��aU����o%_y��\5���V����9��h��;�Lw����:Q�#s��@�C	�fg[зn؎�s�r�/��1NM��}ɸ)~&�@Oe2��Ej$��LF��W���_�sp?�cy��u<�]SR�;�S����5߫	W�DR�P�l%�u�r:�+V�@���s7Өm���nt�v�}��("�qf��q;��j�5,D%Ҍ���-G�%Y�(��?{X�Ŵ����Q	P5N���2H *=Q���*T��,h���(ڤ�?#��M�;;o0D��5u!	�E�ӹ_76�hnz�����/�/�m�#2�틠����{�ȩ�!e�6�b�ө��>�Sx{���x>��l�Ff��T��,;��p7�9�f?�����b����qE����t6��7J���ވ����7�"[o���3�u�y��m�3n��%�b��Ń�;Ίxt����$'�v��ᰴ���ak��eӠ��o߂��/�&�4|�ڳ�������������i��Z*�(��^��Hı]FK�-��/��b���rI�
�Q[����
��8�N���g�j��c>���8[���Vd�(�J<�*K�r�g7��o�A	[m�����,&T7=�W2�M�a�H��j�0Y����0B"��.2Y¶h[��]*�/�5���^��^p���}@�Z��U��_�-k���7rO�ʜjԡm��	�{I<�Z}��L�,=A��nN�M�Z,*�!�>|��dr8s���:'sR8m0���Q,�{�)W��'�,��UTYm"$��;I�d~ŗ9��}�G��6���Ѣ_zwh�lfL�n���A
�� �ݞD�_R���O����ۊ��ز��Rͻ>��l��7[�S�B!�����6��r~'i���g�j��%f� ���e�8ڢ*�e���^ �Pv���mB�ɢl�w��}Q}�g�y��(�e��\C�YS8�F�~4*��#Hm���#eÝA_>�w,�}O�/�G?q���緋���r�����୯�쑈	��,��k�����B:x���D�\��&���]�˖����}g)=&_/D��e�6lp��9��9H���l-,h��Hu�}y($H�-Ә#�tǲ>viu�0�63���aP٧��=l�Hr�&]�S�˔T8���D� ��[w��ch�	ې�������G�<;�