��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�۫k�۸�m�i(b[�{�㇌�]�i�5'�`;Etg
<������"0F��}�h'��8��<���9���-�j����,W�_/�H: 2���x���CH�^�g��$�Z�d�5��K�S:�Y���~��n	��]H�C1��C�#V�S��7Q����u��p�Yp�ľJ8�so��s��v���l�OK�i�ż��Q�LLa��&GȹH��i��B��K،Mʸ�qzZ�a��W�[�17�#>i,�,s�l�>�����4�Z��1�d�^��{֐�S��6Ux��҈��դi�{� zXh����\�%(�ܭ@�0�qyi��S�UvY��V�5��_\C>c�1��/�`�	�n���L�0u�c� ���Tx/]�ʇa$�Km��8#�S1�ܴ��Z��j2q����/�����C��b�*�#FDLr��"�7?������FF���a}Ŝ���_�B����7����d'��A�@#^������ݐ�S�p��Du�ұ�~�5{�N���K�m�m�
(�����������t��rqA��G�.�n�^������&y���e)%���<j��F�1�o���¸E��q�*`���d9���%�i/Ͱ>����1�I�S:�BI�A�+����_���X%*5.&q�$��-L��u ��
+��.b�Q�C[���o���������>�T����`��i����2Ș�q��5��JS���Y��-s���M����R�l����|��/��l>V�Α��Y�����ς��Z��6��P���;$ߨ��x*��~�X� ����E�zPi�*=]:sH��m���Hi����V�N��z�������v��Y:ē��ZN�3 �X�G˿����&��j�`�1�7! ���@U����-m}~G�����+*��B�HT�ԯAsk o	��/�*wۻZ�W���� ������<TnF)��8g��>�{��M���R�<��,+#���5i���Ad|x��'/�;�����e�YJ���L���/8��H����ݽz���3!.���!(�V<���0c� S�&wVm˿D ��L6&#4%����d��M��O��p���#��a�
��B�QȠ�
9��TK4����#�$����̕X��p��t���
���\sC����q�U�$ڗֽg����������@oǕ���C&(x�U�gP�h��}�fy$�+�{渿��4I�P��'jA����N�TX���=}U�4Dz{���3�������e���US 'C��ӵ!��&��A��mT5Q�]�<§��){l~ )��,m�CX���vȅrVP���<+��N�1Ǚ1&МԨV�5���nҲ�~�:(�x5y+�?�F@�L$�kX m�%�4�������q�^�'
�o���M� ��Ǆ�ْ}JR�����2���z�W��X۴��� iSQM����s#�]��9&�њ��1Յ����$���T?7����#�Hu�hS�K��ӊ�̂p�4�d�o�EeE"C���G�n8�6on�U�&`Z����7�ds�B2S/_��&%��f]��a�̃S5�a�jb����Y_�̀e�A8X[+�h4V���l�Y�Uj랹q��d�O�C�ؙ�����`J^��,%͊��xV��UoNzs	zk;���T�"8��6G�HAA�hL�e�t�g6,Qn����rR+�χ�Pv3���[:�J�z�K�A�C� ^"fũ�\�t���נ���mߨ���1��ϑ\!��$<�R)��i?Ȍo�#c�p��XN#e�簱e����
��m�A��wx��O��G��~%,]h{�d �-������f[fb���F�&��3�3�P�\4��ŉ�Q����f�wg��ɘ)}h�%<K�Db�P~����ǖ�	ЩT�a�Y�xh��4	X�.xŔzӳ��?�ML
�Y�/���FMQ/&!��L�4�{�L�����Z�9.��F�L^;�2
 e�s�@U�%��H�葡;*��OAC腂<�7R��G\���1VǨbL��I|�>r���	���i/W�{���;`/���+�޾��d����&�M�H�_��Sz�j������/Qm���E��f��l��<z���w;*�I��!��@c�W������=к�Ph\EMV54�LG��'�h�z�9�P�D�CGp�|��X�P	�^L��U��+�&TA�j�4�*9j$�-�3�r�B��\q9�G-�W��(�[�����W떬�'����ɳ�����f�>�I�Z�q�Aq�0ړ`R4~8?zJ1�b)�^��0ݚ����B�~�s!đ�ZC��ΝS�+�2��
�̛��,����2U���גA���p��%��M��M�xL��ޔ�߈��Ϥ_���g;;
����Y� � %�� Ym���������I���JI��^<��=J�[�Oqw>�g��Ld��S���w�`vކ�w2#�#�{�3CJs0��aZN�p�+�/hql�u�'�i�S�\5���\;�~f��џ;�� �b�VPT�m�?r�T�v�]-�F;�Y ��qKN�T�9��h3Z%P�C��	�(�O�7���qq�E�snBC�]�0p�{P��G?��Z��_>�o�6�?�ދK��lN��x4R�aQ���Z{Ow<)�.W����K�(s���aF�����ms�Sr��-�����daf_��t�)���-�e��}1<��^�>�T�k�2x7�d٦��I�lR���iE��l�T��%.�e1�F���?�s��uu�>���4�넊�G��'
��9{!��t6b���u���̚�2|� W���Ĝ�	8� Ls7�E��������#�T5]�P�;�7l�{����7������m!�"��D���r@�����Ƞ��[/��U��}0���-�/"ƫ(ym�����w�]'���u��
2ޮ�(��P�p[�ӄ�"��<}�?���$�"�n^�
�ڧx���|~���2W����M�ϯ.�e��hKOQ�78���� �mǶ@�I�plaW.�\ ��c(AK���U�}�%��I�9�"qPZ�,\��$����2�7�� җMV>�x7���l�sv�}2hHԉ�W���%���\��B���G�JT͚f]��S!D]�6W�����gRX���� kf���d�CPr�ɏ��7���&-.E�z�h��^�����߫�[X�Ǻ�`�71.@��n�+��z|b�6KS��v8��N���)*7�J��R����Y�{r��T�[T�7!Ht+B�%chꦈt�<f��A�͓��s�Mu�<��蛣f��zޛ$0<&sQ��d\��{���*��ɇ����|5��"��\ct�+rr����Z�($�t2�N��8m��.�(AJ9�J����Drq�I���@Hx�| �٫�B�N�7/՛;�[td�Rd4O@�Æ[cŅ}��^��nO� �'�B��A_��NkI 	F3�]�XZ�U H_q�]3?	�K|~�G��.�7����,��@g!�=��Tu۾}o�e�J�h	a�XyŐ�KP}d���p�U�c+�e��������޻@=)��T�
;4f�y]��gs��;���{�<)��_�E��(��}Uk?��~15�<�N�O� �����>���nw;�����
BŞ䯉@�R���pN�p�a�)DM�������6� El�ު�(�Gl���~����~�b�q3�-u�wfN�RO�v!�5����L_N�h�����c\��_�]�b�ް�l�.�w0��y�rf%&[%����^ケ#� ���$8y�F��>X�v���^���gA�j����߶��runq���+9�`�����֤��%��$vM���r�3tr�g���t�Z��Y0�c���B(~����$g�&*��m��� ����/�����h�&TeNm0�S��<1��,%�c���ADU���މ�a0���P��a�"D~x"ܫ�h����ޣ�K�徑k�r�s�HF] ��v�տ��z^�����U%b��R��MO#g�w� �T`~mҪ�L��i�X���v�ǣ��4�ϸ����=�l��^E�2���"��2����'`|�Нn~�$�lΌ6�oq&�	Xj�����[2̤�o�kx��JZ埑�|�w$������\�5�wxƭ_Lf�յ�����#*���P��=��ݥUe�\z��By����vd���6�rt7Y%/��ĸ�i���j,L!�ށ{���G���"�1�Co�m���
�K�Q�j<#�)��g� �7BQ
n����J=^�d>؍��T<�J���f��;F�
*+��=>�t�Z����(eG$D ��!�¥�t�"�����d���o�p�ʲ�ЭP����>n1,&�"�%ER���%q�Y�R>��amb^;�*X7=Mm��j��,iy����fIJt���Ir�� �8Nm��q+�~W���=���2�6�i�H>~V��G	����f���#Ue���7翝�S~s-�O�q���4�g���9;F�KB%ͩ�Ok��zq�n����j�C�ժ��h���l��ȵC�˞*���߹KS�+8q�_�W�4/Ħ��#�Z��b�3^Ck��H����͎Է�����}��)�����5|��j�n��GW(�#���4m�@LL=�1�I����{���;��>`G a�D� �)���C��݀��}���#\H?f��P䯞g�Lت~Y�aݪ��O���JfK��,���K�p�{eJuqb�6���'���lc���q�V�YU0�0�E��廐���������s20�R-��� l��-����������K�&��n�q�!�Lֶ�~@<SV�l�݌H�":	���4��ME�\���!�)��X̽^ø���Ӄy��6'+9f���D��^�o��ʀ�ɿ7ܟ�~Ľ�zV�����B������|=���\/�A�ا��kCP�v��N6��ZS��Kd;�����k�`��PJ܄�=��2/'(�9 �݀�^Z��`Kݦ~w1J�����B5�'���i�f�ͩN���~Fr�K�����c�E��|y~�o[�������2��XM�,f���܊d�Q��G�����]��)���+��ps��{""���0G�@2[<�t�E�����M����7N�X�\����i�Y�Ќ�y�jj���\S��({3��M��X:�Sf5�);0�5�(��dO�|���XF�9�d)Z3��"q��)��g��}�Qն�,؆]������ NwO�%:��ӐB��/��=C����mɕ��11d?�7�Z=�64�|���e�u}]����������o���#����m[VBUxԚ�,�ݶ\����Aq3��.��*\���_�h]+?��!d*lt�ls*V��%��_�;������:K�<��D-$LUrѠ�9)�t/�7K%�Ԝ.p��)	��hy���]GP�V�A?��1T���$����$Q�n�|;⌖O%d���0~��U��,�4Mݨ��Q8�]��ӥ���K��(�&`Qh/�6�y�P��dZ몽���B����0�������վ �� �����I�nG$��pF�bxT����@)��'�Q��Nm� sU�0���7�Q �Ey@ %�J�0
����`	Y�!R�mk^�|��!���4����:]G�Wȶ �d��#:1�o�`��������!�nZ��Y~�����v*�g�|aQ"*��9�J{<��z;��u����P��_[:����h�aeZl�'�( ���l-�ψ{\#T_%zM�/��Pd�����n9>�r$�Q�GE��+�3�rc8�Î�����c��6�&�x�{�N���,�L�ғ|h��ӎ��܋�oj]YG?QZ\�\��}�\ҋ��6��3�̃��v�C�nF"-pe��=Od���ht@�?)e�������ȏ�?k�8ga<�!�/u�£��[��KtV���x��<��r�0���=��'͵w�����jY3Ċ-Tu�c�kFg#��1�K5�1��}^r���d�n���������(�=���T0�0_+�ZYb���
�����C�mR�~���c���J߇�2�7��ò�tT
����*Sޑ��"��g���zr���*EӢ��PuM���W>��[&����]�ȿ���S��*��O�#��Fg]�^6���p�is޶���b�Ŧ��
�5w#�m��*�����Hb|	���h�T��~���[A�ĝ1�	Y��]ϊj���{UpI_%��$�_JU���x�;�O"$�jc,i�_�ĸ�uع��T�N8��ܴ=�-K[��Z���_%�Y���i�ɬ>+��7t[*�F��@Ҋ�������+�D�6��`��f�P�_��)�FUW��Wnمr�-�ƾh�i��WkH<�]):j/N�
��K�����A�G,����)m?&S�q]�E��"�S��̋P��)`3�~��F~̵BL�6[���퍖�m��U��V�
��#΀ʭ���:؝�d.�7T�_��*���!.P�w�z��\����X��t��1�+Y�^;��?�0���.�g�0�yR����V�p�t>�){��� ,b؃'�� ,9C���lڿy�I���e� mN��xyn��(��[[����h��b�(�R��6F�Ի��Ըf���B�岊 �f*3Cs�c�,�P4t�;�Ot����F;�Z������A�Zk�+&��hX�9�G��';�+�!�/~���a�:1	�:mk(O��=�[�z)0����}X8I4E4���������A<3��]1�m7��<g6\��v#?��Q�偀��7���?^fh�j���Gw�ذSM���*�v��u�U;D��/�[h���ğo�\��S�p����t�	Q��"nP�E�g�?�����o��9T�i�^r$���%h2=���D��H�\�&WWR)����UP�a��	����N��+e�?�|�"���C!�A�N�N�N!�i�E���h���G�㪘�	{������/�=�T�mR�����0���� ��-��}����"�Yd9i&}��)�+̔Z�J����Be'@O���=��1pb�<��X����h���X����e���î����O�F����)~�PTj7l�I���b��."��y[etD!����:E+�#��>�0��#X�M��ġP��.W���0��K����������Rp���,d�$}�|'�.�<_�6-��b���b@\ʦj<�3���9��tx��}/*� ��ǑI���:�U<���|�mQ�L�6�W6����-T�+|��{M��M�?�i<�q����S�1X�QDn��a���T��4�fs��1���ڜؐB+|���6��ILX�T�V���,�0�Cx��vqP���|�0z��?�L����u����a�09����t�4�jubWAU��M�P�����ՙG�/v4�9h5���gm5����>�~y&����^��*N��P�T;>L���WwuϪRE���OY�p�Ʊ�k�w����Si�8(��LՊ���D��&}�t��5��:IFb��ŽC�4��=<�ߗ
����Ú����F�Dɷ0��.R-6���U=�]4��G�����kvw�\;H��\7���l�qGr;dH c��OQ:/�֭��Ȉ�9���ك�ݼ��������':�4h"B,"�#�J[�����nL�c�8����`/�È�r��z!�L���rU!5lv�k�L�0�OIUt����b�Z��p�+�!�\��3رF� ��(�����R��WO¹�Á�?[���8��wtt��-zl���1s(�����f�e�U*f;���-Й�)S�m1�#1�vL0-��q�7s�����l���yŰ������Z/����&⩎r�@1�v��yL�N1�&�����1+B5&,d% �D5\Ec�}��L��]X|���o
�4mb�pC�/G�*w������V���T�/8nS�yZk��,v���%�i��Y���v�O�p���b�@-�IW��'4��_�CsOUepp\�����&���Uc��Sn����Z�P�]��.`�D�:S'B�_1.i�־^{��+����7)*�#Aн�OgQ|Z �u+7��ݴd}�E�� �/��c�)���I�Օ���V24��_�:��/;����s%���w&I|Lx.aQӤ��p��e�;�!Ei.�A�kL�a97{SArx��Y��KlM.�[A�u!�l�h�C�E���Np�9��Ր�$�9���`����Q�')Y�(o	k:�oܧE���! ���T�ׄ6҄�����k(�1wqɂ�RtHk����$�Vw�G�Y�B2+*�nY�m��6��S�`3�':�dc*u��u�>R��  �W�'	�����"���ظ��i%am��nh��O&s}��iE���n�TK ���h)��ZpG�� ^��!��&'o�4�>sԏ%MF���r���T�n�ͽ%�K�QYnN

��&�"	�4�� ���W�O��;�t��7��TX� �%ubϻ^�'�.,��/Œ�P��\�IN_��QĨ2EE�^�o�|w�o�LA�%�o�,*�J|���^�ܩ���o��&�1�T�;x���P����_J`�� 	s�����Tf=������X�cm2��Ge�j؀��ӌ'��?�F1�xE�#��1�j27��xu��*�����s3����	m��vR�HZ"�� C�B&,��Q}ɶ&d�͗�N�AD����&���YH��*7��e���3�c�:�)IF���gzd1�B��lN��@�7�Ŷ��a�qA��v�1� 7�(��Q~��Q�|L�d�P�W��?���� ��Hl,Df����&�.CK�N�7[���BmX�k̶\%�q�����rï��3��zfuGoJ�q�`:��$7K����qz�*�7��؄�2��M[�̄s��0��y!�1e����Ȍ���1Ί����5�?7"�q�*lC��)����jn/�$�$�8����̯��%)�Wa�i���ҹWEL��R%�R���^���!�\�uXE�Y!���0�rwL����<e�����w˖���gM�h��$�m�l7��������ֳ��)��:�j*l�n�C�2�)E���� ]
p�%�9�ʮ�F���������+�
����1�6	u���7���f^M�R2':�30��-�́卅g_�سӗ8/ �&(����^Q
|�U�Ka�����۔񫝰ȨNF���V���V�2Az��ܙx/�3H�+����de��@��� /[ؙ���Ǧ��=2���.��y�E���^��gDe�H�tL�{�R�?e%���쓋�|k������	z�#پZm_U�?=�g'Q�䆋0?G��n�-I�3�6�۹{{��*��Ư�0��M�`����79f�2���'3⦣4o�V3ų*Y�1r�����
���@G��S�'<�P;�6�����R�����U5�n���7��ͨK��������F���Ƒ� ��z��?:`�z������6kG��T+]�}���6�u���qe�ºh��*�0��������uJ�I�z4���čuk� 封J�yUu]����P��C�\�����X�.�؍84s*6�����T6�7ս2�RB,�7�N��1����w|3����iw4���a8�X�C����p���йFM�%:Y���o�=e�a�n�9��������it��zH�Bcs=ӿ�J���I,Φ�M�c��|���7S�龛�>9dn&L��!iJ9�&�'�=�k�����=�ku�K��,
�G��^�7@����΋Z��Xu���?bfr�͎�>��:>���]��~k+EZ�R�iK�V�#�$��6��9�4��R��%�`e�J��6�Wܽ�®Jg9·�kvDӏ�֗��݅�����f�� �x|}�Տ�U��At|����`܎]�Bs��&s�h鸹��@��-�l�"�2�c�����|��MҘ�z,��ު𒝤��j;4:+7�f��xIJ]��skYP�I��K�x��tųT�bx%���1WR���r��%X��|����}�-���R,m���8, ?Pm�; �j���;0ۊ4�m����$eqb�y�>$n�͈���I��څR/C�֛�j��K!���
�*�b���������%���)�!9|���/��;�^���֚Z�,[����F��� ���B݀xXԣ��Z�$��F4��-���R��6�V�b�6Y̫�ܤp�o_#&9����ͬy:w�$;��4d6S�x����<4lo�<��Ծ�I��>f��r
�Z+Ġ)�|&륕�p|��G=d��p���<���)��I ݘ�ꈾn���1��4	�d��T1�I��Ĉ-�#�����0�#��p���C�1έ�ۆϫ�=���8��x<G�mܼ�k�V<B�Ύ�{�\$*O)9Q���tls�$�p��M2��oy*?N��׋�x�(���'��D�53$[!�:���m �����n'�6c*^%z�k���|%=�{��^��,|||S�8��X��}�u'� G��8鄔��Hj�S��	ΰ;����d�T��^F��)O|:湛�YRQ�ɸ��H�y�n(���X0��%L<�$���:�u�jڏ�4��l%_BI���7��v��`�H�=� ���gq���W�n�XΌ,B[�ث%�"!*O��e׺�Fki�|��Z���%���#B�V�������^y�ܿ��쟐�����S�.)'��ꠁ�K;�@�xK�c�0�h��܌f0?8�^Ta8+zJ,�x'�`Q�t�,�]�~l�E�}
�����7l.������*�˗Y����ze�?�ப��}�/7�/c��i��\�m��3���1@B(�������J�<^]3�0��?7�vK�De.�N0=�i燩�J�8b��#���4X��A�lbJ�`�p�8�e{�\M�>�nu{!C�O�(�4F���f�lF�� i���	��,��T/��I��r�zkv��J4����`y�a��̻�ʘ0B<����D&���pif�=�H�ÞSݸQl�QP��1�bQC�P �Jo7WAu����p�vZp~�5�=_�+�| 7�e�7=��%��#:f7s�