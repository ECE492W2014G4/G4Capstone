��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P��v�"<ߞ��&'��k%P碶�R�ӣ�sĞ������FY&[~x��Zg��_� ��Q?�^#E��w��]�ǭ��|�ǢGe��/�1���C,��%�.ipjh�3� m?�C��<HW��@�
�\�@�q�����6���`p{s߾:�8)J9O:/�P*���Y�S�q�F`1E�L���0�<)�e������&߷�Tې]8:]�r��{0Z�^�¢���v��٧�������/5��ӚU�G�_��@�]��������`W�Q.���'�������Dͮ�?�#��dF#���T���h]:nc`�ϴ���o�j�Ҏi�?w��|��2�hs�7��ҥ��>�u��y��|R[S��*bd6(=0�d$e�m���vm?"^e�7]a��p9K����2�&07�a\��'BF��*(���/�V=;t
pQ�x!�5�N�C��Z�CK:Ȧy��x��[��zZ�nyLR���|����2�C���/r�aN��V���]��06#�����_9n隩֗j�9��t�A��! �ʛ`���&�� n���p|�q��]v̿�ݤ�f!۔���￝o/LT��s��k_l��q�k�rNv���ȳ~��Om����~����Hi��[���L��n�J���#:B�j� �J��<�s��ﵛ�I�Ә���?7�R�<�i�M��{�����_��%�eHPۓݲ��~f`B������T»��J9^�nDזM���!"�!�/��m���lC��*I�\��q���ȭeo�%A6�|�k7�a�����睟C��Ò"�\tj���u��z���hs�?P��w�n�&���h�]v�o,�r�������<�����*�I�7�.�0������[G��ЫID��fҁ�9M��Ć��T0[B-���%�E��tU��O�6��1WČ�]��3�U�J�;~v7�dHrQ#��xm-�����k��?�j��%W,;L��	�fT��a�wW�A��BX�q����;�PNO���"F�a䤰u���o�ۚ���������|���{��nh�:.��ʜ��w	�mW�j옜
��ܻf��Ģ����U����)�I�f�jt�����CM�)��Ƈ��s����g��k�;�c��Q��AU'"qzx��E�K_5'�%�O��b���/�dTŭ�?f��C�1v���M7�E<|)dᷢ�}�s�ix�d�0�t���G̡E2���6+dk/�\�:/G)�˃�q�'-�F/�=g{ E�Eqt9 U�c��@c��f�J�<�?_���w����;~;��)B�4�D@�	@��t��ˡV��d�s��~.gM6-�N��x�L��Ռ��1L�7��鷶c2�3R 2���$4��t j%J�T�����q�i*�3-S�A�z�$���A)ԍ�Ey���z��}ۄ��(Ƚ��ܵ�Yb��K��f��v- �<�MX�s'�	3s� �Ic�k{�ٱ��Eِ�B�(GO>7D���_ch�vԼ�9�O�i����������\)��-B�k���1.����L�r�]Eob�~��G&BW����}������ԯ!<�iHk��+1y���m�/Qf�U�}�!ֻ����o2��Z�P��'^#bN̡��Ռc�cΤ�ý�/� 7tH�l`�D}!��y'Lę������BCF�{���I�g��{�+�=��&�6/B�!y�m�P�
�&G���i�1�zD[���Gb(�z��M��Bb��;?�:�KZse�����eY 6��	���i�Q�Z�N+�|Rx6���(Y�~�L�i��X�nU���"�V�Hrx_�uH�v��/���H�ZFUì]�:E�2n�O/� �ֽL葼�����fg��{{����L�nې��an��%�����ny���A�� ��