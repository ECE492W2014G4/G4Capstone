��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P��v�"<ߞ��&'��k%P碶�R�ӣ�sĞ������FY&ƓhҠ��?���{�??��F�ʭ'�Z����c�VH3�g:�P��vEn`ĥX{�n���V��1r�jft|,�pX��Jҧ������>E�7�H��z{�쏪���pO/��2����9���8���@x-̾n���[���[ݑ�Jl<�@�F1����Z��JjP%%��@�H��%\]̑�>
E�M�="��ֶ�g��,�֗�_�l3U)l�à�	И�����ZB6��^Fy<������AIб?���r
X˽����:^�dW~�\������m�Vg����u�'�ˎcD؋>����y�y!HUF��Tk�Y��Y������T3j�|�xYO���4O�8e��rȫ�u�(	hZ#�ZP���s�0(.:�vc����Vp�)u[$����&?�﹫(a)��D(���D-�{�Ϋ�2�f}$\���p�U�V��ޅM���z��ċ�H�����2��D�����E���ٯ�����k�cd^�V�$��t4���R󉼠3Y������*m�ʼ�%�7B0��B�>I��U���Sč�^���C,W�z��=�,!�Cu�PC��Ѱ+���]�o��jϢ-U��Q�H�2�{]vUa*���0�:�'��&e��"X��_�Ҁ �<��Yb>����،�����|�MhG�UǪY5X��;��kj��R���iRi�d�1�-��y� �Ё�d*E^iu�¿�(3�()t��|Z��vM�g�^��z���/�*���1]�wm� (���v�ܾ�YCE˶�ߦ:�n�P��'A�~^g�<nx�B� �T�s�{���j��Ѻ��\D���!���A��82�6X���x�L��Q���j���T
805·�HP6X1�X��:�0��X�����QԨ��v�=s���7(%�h��V�1���(�'��F�;���Z/���SԦ��d�P�i���"_��5cu}��S�vq}&򈙴[|�L�T�a}l����L��m	J�"Y�e�B��)�	"���u��y��BǮ ��00 i�^n���X�ڠc�N�u��lV^��Kn�z��7���u��|��e�"҂�2&39��Z��� Z���Ĝ�eh�z;��Cw�=Z�C����u�J����nsɴ����p�ᰋ:��`����q�_ϟ%��� bS�v�=����i*S�<U�B�Z��K�$��Z/�`}0'AJ����<Ӎ�NZ��[�I2 Y���rP��Ky�C�Ϟ;�ʙQ\p���X��T�0�>H�Ȳ�_�۩pb*$��Z�֟#�5d?�;�R��lD�9�Fe��b�\&����SG~Ig����lPx��m�?�{n,Ȱ_�\6�d�,��P��-�� ̓贆js�7����:�{%��� �����C�g��9�t{]|�q�Q�F���I�!�����I@�^�J�e6=����R
}l�)�!=�47�b�9(�w�ϧ����3�]�HBb{V����@���ݷ�l�����w���\�!�9���S�k��9��rGȅ�{�j���� �g��/�u7
�>����( xRb����#I�˴NA6����q\$�#HZ���Q3�.�$�g�`�g>��@��m��U���#e�=pq|5��yW��D�Q�}S�
?�m�]?�e�e��2
�g���5@y���h�-�VV� ��1��B3
͗�;�mئ.�^^�W�f}V@���d��̚��qz߂ע5.l�6��͵��� �׃V�����g�ٲm�f7OWޚ\���;�P_|x�p`� BJ�@}H�d��6\�J�����1�"N����M�U9u��%�u�5G>�<Z(f�����������$v�|�ߒE``��ۻoU%�����Q��4�Z���W���w�I|.�ш�S��d6��H�x��'"�vA����c�1Om�Q%�����;���:K�-��%��"��O^�;`�)B��+�:�g��^�-����{Jt���U����Dͳ�R#L�7��Suhq1�*^�b��ׄ`0V�_M�,��p��'���a�n�W=�~ݓ��P��g�^_Z�����@V�V1�'wU�D3�w��*��������xZ�������?1؏��R�_��h2u8\��6���X�ot��l�k��7�K��l
Y�'�&kDohv������6�#�n����ɍ��y�{}��
4��1F�]�v��K���P��H��f�,�5��D���O�$dJ����#2�r��CH-���������G���}��rr�a;���b��NAD�O~�8���AC֩<���D�#�Q����bTo����`���IQ�v�A���,�W�N���J5R�n�=
9�=-#�kL<ą��Z��7yi���T�W��������|f4{�>�8�U����/k�<X��E���ys� �R:�UtF�u��PL�M��	��e�K�4ݘ�X�3c0@J���ڮ�Pq�1����N�=c��U�T�+Aj�^m��¶���be{t���K�v���^���E�L�v��>�[��!���t]^��/	����}�"�9(OB�P���~e�H� �~��o��T��2��ޥ.(���LFt{�샪�gJe8�
�Ct�r�H]|Ƕ���.O�j"Gs�-sD�B�������%��Q���V"��u�+!�d��+ų$��Q��~���~�C�4k�U�>lUd!>CY%�S����Y��!�<��WO:�X�K@���a���=� ��ZU�c/�B,&�n�P�����-%��$�qF�=C^Պ�o�!�� �>m�'�wR?��?2�R�\Ќv�����
�Mw����8�g~̢�-ed-g#�,]��e��aה�_j}1M,Z�Q��H��+"�%L���/��y��6Qͭ��b�?�2� ��T��kt��K�9�K�g��h���e�鉢�F��%�z�]����x��q!_0������UJ�S8�:�J&�i��r���fT�7� S!ÖR���v[ݙ����5�㨌�7B��Ve�e�S3�sx�D��7�xіP�hD��Ȉ�Q.�Wa���Z.�����@�y��rߩ�}�}�j������"�;+���.R����V*Lx�T�h��X������U*a%G�G!O�ڡҸ��XBq�&����dM&�2�~3��<_YF��_�˂es��>�N�So��̖9���pbK�e��U'_{���v�)���:*��s���V����n�`���]��-�:V����z�v�X�v��֖��c���^j����!}��ɇ�8~�$�������#��}�@��]��`�7����")[qN0'(LB""�d|پ�#�ih��8㟦U�>31�v��_S�X�zp&j �3p�gf�����F
=��^(�Ud@$d߃O��ǹ�Gi��&Vn������[�%��Xe.0������A@�}���s���)KKb� �M��������ή�%aM��M�������Sdk'i�2s���3����<7,r����xH0���l
%����V��[A�1e}!I��;�=b��[Ћ����U�`zwX��G��DL�Hh&N�p~<jQSSR�D6��D^�_�B����Z������Q7JI�P)-~Q�G�����>�>B؝b[li�Ά&vt�B�e"V� �">�mu"`�ت��кN��O��c�%�1�q�̺u[4�u��3��}oԯ$X�+ޢgr�����W!�j�?޿C� '�v��wq���u�T�rA���\���vz�]�hBm�6{���9EKA7ˇ5�*7�pD����D.Rd�~ES
J��쭗�";��;W�C����{��oU5�6�>��o4϶������鿤H���t��P����n�5i��zN�֒u8��\w���y4Yl���l}�Ʒ�:�������~#�S��3��H�^4f=��mX1�m��%��챽��:Z!�1f���P��[Y@PW�#�z{L�����j"��	N42��?B!r�?�h �$L��Y�Xm G$�����lH'�Hi�y�s��)�R>.[�y�7ޜ'q �uA����ʙ��:��@!�آ/<?��m�������M-�?
��U�AP����O��X��ſ�+�N��سK[2$�[��K�[l-#�#?H$ƨ�[bH6Ô�,��#�fˣ�^޹d��=Sk>"�����UUT�M�%V2��^��Z�ਗ�E#�t�0$��ga�1
S�T%\Rݍ�eat��:@.49�^����%����C����6"Fn}���B����H���[~I�L�U�>��E�3��7{��VOD%pG$�*�6�:��6"�:4L[DO_ɬ��-��!Q-&�����˄_^�s�Dܢp�zH���Y�SJt��eCt3��8�dQ@��~���ۀ�����Z�T�e Z"�e�OW�?�?��4k��·5q���K9f��(�NZ�'�u
'"LQv�	F8Q�X���-#�(W�eн�	1��,�=sS?����nZ/��t/
H%��N]�hb�{��c.�?ʎ�/&���p������ED��\ k[���#��{�)�<��<�|p�g���=Nn�����#Wɿsaĕ�����Ozf���A3����@VΠlh����K��hq���
c��tJ��G�����*���=C�PEM	�Zn�h�EΩ��e�A+�?%�ځ�ΥMv�2nֱ�MÄ�U�=�5��Ty�'$PC2C�ZXx�4N�{R��N��Œjl���P�M1�@{�HR9�.O4 �ݢ�v-K��k �+v�(��C�F��?����D�඘��/*��E=������+�;m�Aʪ��Y��Up�G/�>���?���؟8|�\&��/TN��K���M��!�����ս`��,���aB��K��cp/�j��R"l@36�d����/:H��7�xL1|�����#�c˴~�`�ݖ���u��>+|�����u���������\
�fh^G ZPT�A2"Q@m��lS���S�a��@4-6�"*����#�iSi��z|�/��֠]�{�q�E��0>%���C�uYWX�!�$�I6To����PW�p�'�g�sG�hic8P��·;�2�ip�ێvL��\�>���RB�$�E�sFj&ǎ�f?6��I��/�4�4�)8B�!��ܯil������xX��dI&�xL��tY�B��J��T��#�ƥ�p�0�&���o*�-�񮽐ppas8+�/��P*db��پ�ނd`�=��q�@���,����+�5K1�|�|�uq�_4�ur�7q�KY���ӌ��M �'m�S\[�i,�n�"���bO�c̨C�ā�f�6;/��'��J
��m���ǕR)�����2 �$��6嫧�]r�fT{����G����, �����P�%�o3h��XV`q���WG���Ob��b�_��?c�~�0��Vv�UZדZ�:>�Y���P:H�d�w��\��bm�k������%����)���d��b�[�n�P��s�q�/�������ʽ��fT���g���:X��Q-�h�*���A
�S&[_}�F#?���L��hd�lb����%�S�P�=7�O��d#uv�~h�v��"����;+��W��v�l�
@�K�ߕƯ>�TgrG*/�4�t<Y�S�GG5��.*?�Ю��1?y�`�D��,xBI@�JG��*J#��]���_^y�����*_���\l��TCLf�z�48�ڸ�8S�T�ړs���B�b���a�WM����=e��ݾ;�'[�n�q�sFU�vDj�*�7O�Ǜ���={��y�@zj�����2�5�i}�Ό�<Ys)��&s��I��aM�����Z�		�Lȳ .<���C8��ڮ6�
-��K0���=w��	�H�8n�i��x'o�R��JP�'@�a�юc\yxB�b%�}�쉪�o|Y��Kds��1�H����%؈xF��~��dj�H�Fv�h�������EB��|�1;���L6%�����u�ml-��
Q�䚿�S�X0����%��TT��PQn�1�d���X(�޾�3���������'��k�څoA���uܚ�Ѿ��I�5<�I����sw�؄@TF�?�|k-����h��_89��S�e���xvn���2W�-[+�v�_�A��8��_�g0s'0����A�c"B{vj�����^���~I��G�g
zX��.��L�kB2t��I��|'g>�ΐ�1?@\7ڷ��3���:]5�9��Ȥm���ݘt�@ h�*
����G�ʟL�V���ض�f$"8[h����R����=	A�x�}ؠ�N) R���XA��]ƫ��G�s	�d��NMǾMvz�ʜC��M��E�_(q�eޣ&��k���3B/�h���} ӎS32�u���70�"9�q��=�zS��+�:oV���C���Ґ �JK�{��B]q��4�<��o����T[��h+'	gإsl�9��~�X9��L��ɓBF2%oIq}P���w�>�lj=mէ���Q6~��+����s�+��Bݽ �c�v�,|�2�#�OL��ݡӤ($ŀ��4+3f�����J����mWW��!^v��������8�G�Qm�y&�S�����^kTʉ?J&R��Z��(�a��zJ�6]�,;$��M�e��ɣIq{�K�$�?U�x�r:��D*����^.ْ[Mt��(5�]�^���J���%��t�K��T[jݡ���fO�e��K��h: ;��,o+�%\��#�ե�d������q-��JU��,�!{~w�r}��.M�9���Oc҅�0v򓦀b�N41��*:�F�T���?��<�/�4ϒa��b�`��Dq�NBġ�w�I��=Y�D�o�_w����J�gj��,��C�~g>Y��T]�_V9���J7�ʚ�׮��y�ڥ�6�5��2J3����RES!��C��Rmջ3?�G�Y��Gy!���A����#�N�%���˩����`�i y�/B1�`��HB�S�=�T��d���ǝ��˓�S�o�3לn&o;Ď;�\>1�[���$�V����k��'���v�v
���M".M�nV>i��߫���?"�J��)�vM�_&u�����A�DT��]$4׳T;"q7Kξ���i�7���#M���ʋ0�d�"K��%���Ѽ�D��|V|�P�i�	a�e��uF�xc�w���z9"^'�%|5�ZRԛ���r=Я
�B��G~�����
b'y�}�0�7�p��\�9�I��
3�є�:9V}A�~��p3�xre\
��&:�0��8�ϵ��$�}���g`��o�
s�������$��4Z�vAz���;��E�Ӿ�
�����Qc�O��ԍ��E�CC5�����.�����뎯�~̴�V̛� ���jN4��������vN��$Y`�3�����4`�;����k�w�-�F��bL���Cwo�� �H�d�Z'��j7�/���-�M˫!���ێ����`��,��J�`u�z+��ޖzb�򪳂���Jd#Av�9�Ӫ�r��
�ʗ2xֈ�VOx��f����_�*�������2�':J���a9L�O��z�c��p��zp�<ٳ��z��xY�;W?}�2>�����!f���T�����n�Jt"�4�Dױ\r���7�ͺiښA��	@&C�q�V�^.�W
�k/��\����7fJe/BRSJ-L��o.4
���X�>��	u�[����T�T +�5	��a�@�oy}�2�*���$��H�����K>&C �b���
o8��"�	I�4<��B��i( �,��n����*3(��a����\L~����`<���K/����B��56}g�Wb��F�������V ׃d&��U=v�����̈́s������.�>�!�آ�_+�:iu�eFg��8c���A�q�j�!KZ��!~� q�fI|V�
oɓ��!�j��xͽ9�vB��lw�A5�~(�D���l8�L#�<'>�w���9Q �]k R~��v����c��ԛ����M/��mע�t
:_Ra�9C�$ J��dA.�3�w2�y�ţ�ixY�r�E���]�=�MgR��Í����0�9�v�?��O 5&�o],Vd�Jl��؂�-��b,�v�T_�Z�bvW���M��̓�(��+ ����'�尃�z�ɸe	]ZI��Ar�cDz�����.� f1��qM�HJ��Z_e�R �<˔��!Zk$>�(���h�ڠ=Ĥ�@�?�'�[Cb�E� 6Qx��%0�ߝ2�P0�-��y?�qքw�~��2�1d��85lF�ETV��/K�3&0���Coõc�z� %���������$��!�W�0,�oݵݸ�ʔ�VʻKQʊg'�O��?�M���9�gw��@X'�Ʌ�h0�o�Y��N�P'���������-9��6��X�~0�Pb�dx�hn��� ~�>}�g��e5�Y�t�c�ܛ�ɂ;1���F͏��w.�}�J��<�Q,�6�@%j�i �/��8j
	#'��3M��%��ck���2�f��0���}E���$ѥN���?��4~~k|�_{�6=� �dh}��2j�׵V�AGF#�1r�l���\:���BZU(�zR4C�\�!�6Ž��Vo��%b��x�C���Ƃcd���]�: {��ݫ��0�H�͖�!c\�oR��	z% ��l@R�7���$�qY�^_)u��p�ZP��&8h�h,rDBD��w���1��Է�28�ϲ��$����j������$?��H�3�SZ��{#+Qc�⷟)_�ʝ�{�����_���%�� ����7观��B���w��t3h*`|�]�D�s��+Ob��s+���/^uʻkE;r̓����8I5����]�r�Q��mb?���%U�`��q�~ �<"9�]��h[�9.��)��1tq�H9Q�?q��#���0D��!P4pF�΄�I�n�et�9�*�6�TN}�W�p4�PзM�΂+�^(1�\�%���BVڼo��)R.;�1RL�)֠�F�|��?���v�5;��^��m���*�>���J�k#�� �h�){Iv���`���s�E,��) �%tӓ�Cd�M�6T�FzHj��̰��&�hSk�>"ک�)xQ��p	��-΋`c��F�ƥDev��Y��A[;��WP%�bC�E��ნ��e� �c�Ț�Xv͆���f�r�3��K3���pc�ވ��щ�УS��M��FS�j[d��3p�����+@U�±�G�;�n{�fF�i���4�%˲����n1��؝G8E��ر��CKTT\�F�-M'Aơ½�t�� �o��p�-�nu}�A�O�����;�B���q\/��b�g�;SKf�߳v�M������]�g����'<i���c��IpS�8�`)W*�*P��&Wy��2h��5Q�s�襾���� |WF�"����N�3��Y�F-�&�ف�)�=X�:�gZ��uH{}���>=>Jؐ!x 4�7�����"$�JeM<�FS�=��p1�����s��~����Q@bi�{j��N���R�������T��6�)� dظ�ن������}c�X*��w�}�ȟG�F�y2z~��&{����U;�/,y'�2��3�5�v�4�?9c�� |���#{Ǫy�;2�����Nxӈ����`�J�gZ~��N�j�P?�
�ǉ�P����Vڮ[ӱ�z%�i�Z� d���ܺ��m���37�����RFdi��K�9W@���ՠљ�KT庢G/���Z���z��4$1���f]�9�bqQ�����ߍ��r���Z�G�e�h}8]�_��155�0��D���TŁ뺮nr`[���.�����g��xHgt�~��\�͌��v�ւ��[���hoNc;�j%����sǔ��o`r�R*����L	+b}S�7,+{}
 n<\wR��?"�)[r6���Rmή���Ie���qI�"yI{���Uab<��'�R~�7��f.c
ʪԈ�8�#ld�@�5R9S2�4����P�h잝4k~�P@s�4��	y ,��R��JH���Ar��o(
4�}�R�D�nZ�� ���$�u�|�'����Ag�P� ���Ԏ�����I'÷���1��M{fad����F�=��:�2��@��x�WT.��������)n�󣇬f6�r�TGB^D�%@�y�+8y:��o�_����Ar�9���86���i�(T< ������ �։f	1�������:��q*�AY�
�� yù` �12
2-e��,H��Q�592EnCM\���&;<S���OáW����5���2��s�P�F�[��TZ�u�m�Z�����x��\��
l��-;!,���#�Ά��h�f�b��f�?��Q+�10�M\O��{EeXF��@~W�ܡ�r�a���m��3G�%C�)��.�LE���~pz����~�:0�q�M���Q-P�?e:�JL�/�X��2<��dY/"*�G0�Fb�Q���r��<���}_[^T�����p��}N:�����_pe��~��%k���,&ki�<đ��.�� �Hj����c�������%����������П��8kQ��91 �Q�6�hF��#���j�T�nW��+v�ȕ��h�����q�	Ɩ�����Q�͖\� �UIh�B%Ň����ꇤ�ۻ0��Y�����Ko�+f^2��ad1�QXUe��.::���-9��匤�+˘+��ȽZ�rHv�e�ئ�6w�r��OF\��q��qD�����7k��w��ӫ��E���[�G������i�=)���K����~)�ӂ#�߾z&3�$�?��H�}nA�d��bO���q�d�E&�H�*G;�'H�[*��i�>X�a�:�ڪ�{�M��6�d�5YF�Ø���/���!a���Ő��,`��z>��ȥ{X�6�o4����p�\���nlh�����1_t��4&,�EC�䩒U��5c^�~�BL44�9�{�����G���g?�5+�1pFƨ`�t��s��������ezQ�s!Bu/Ys=���ߡw>(83�ʂҶI9%��2�"^��e���ՐM�mv�r����}V�p�c�y\"�9G�.ƌϪt���J;����Cl����(�AݳԹ�o��j�Jx�*%���OQ�83'MK�1��o�E�8�����w�����C�U�r#��r2L��m�5#� �?�	�ap�Y�op��ق��)�`F+}�@��D;�B�G�̨1���]	��E-"`E��o&�~�0�o���j�N��p򬉓Yq��	�|���4˂��FN�c�t��m�Fמ �p�>B �z���Wcp�>��J�{���u��6ؐ¶�T�V��I��\XYg�i���L�� ��6D��`G��5��j�x��U4����I�����:��9l��v:�7u�2����.dkR�dz�j8C9��nW��ck��HfT�=�����xQ���M�٩������F�ݟ�WumqV�-f���J͡(PÎ��3�����XR�)�'΂������Cp|u��w��m_�A/	*�翇<�Y������>��iB��G��u����^	ɑ�H�Ľ4"�/��K��ʹ�- z�kBs��:��f־��7�{ϰ4G�6���R	J�.T�?�pD�3�T;$�6|������V�������������@�c�R��׏���A0v+"�rQ�^'�U'���~�ҪE7�@آ{�	��q3w!A���ln\��5>=..D�!�;&��=���&O�;�6�w"߸�j���.*��]mepʑ�k;�1�Ԝ�[aȃ=��"=���T{]K�u
4� ��Ew3-a�D\����������h��Ý��XV��6j��Qގ�K����K(t�SĈ�-,��,N-���EU�:���f ���wVcyy���X���Wp9����#� =>)��
��3��l<�~�gJō�i7}��|�EU�+��2v�	�ȋ��>���ZH�-y3�_%��b��6<>�Oz���|�S�
�����,�@��4����Cgg��:i5X8��J?g3�����a�V�Mr;�P�,����9ӱ5�E%G2ޟHU��ֳ�a��=���JC�tA 4ŧ�.���i�|3��,�`�������o0�
L�b������mʹz�J��й�`C/�Ͱ����U�u&�4�(lWȠp���PX\�W}=���B菂��r�uwdۃ�|�f^>��O�gÌy�P���)��w��e~>�&� ��;�On��~Rpؤ�>3rѐ.�]cs,O�����$x��$�����Ŭ-�&A�NrǗ��
l���O7!��~\�9��g�Son��99�����$�;����q�����V?��',3���EkSe�l͌��tB^Z����e����9�Qě�N.�i��*I	1��Y��k&��
��� �p�k�%�:�X�~b�~�Yв�P#Sl2�3{���.�'�#��dN-I0:�D]8֣�U�v�3p�L$�ϟ%��c�t{���W��W��,:gq�:��8�K�Qз�BZ��s�K��fj-�5���kf�8H����]ͮn�_������b��?��+ G�zT��|��[�����xȁ~ʻS�l<K�U�-f�.�����������k ��i���>�������Ӫ"0�����KP�����R��$�k�V':���oB���y'�	�?A�p�����J���d�jF��r�CB� T4H�ԅjf��̎˪k�OYr:��/*���t�_-&��ç2�ٿ8b�=��?�
C>c߽9�"n�H<��3���5˅g����)�w!7K�n�ܐ�����O�Ö/��:�G,#��Kݩ]n��t"+����|A���C*r��⧲.����+A�����Z<���ˌ�FA��.Ϙ�
�
%\�J4��l�.�.�D�m4�y�n�8�T(�N'�������G,CX��%�7�yT�a�8D�%��&��&��<T�
�Y@�p�Z��W�茺l%	o��������w��:�^U�EԕE��KdY��,���@@wtr�loG+-M�L~_R���2G�df�c0x
N�oWQ��r��,ĉ��{p.��Z<��KT;=�S�e�i��$܂�I�&ʊI	@(��W��.o�o\5,�dI��Ѐ�oE��g�<~"Ͼ���tÕ-�`U��낞�#�0}-��[6|��w�:�)Ld��!U��jx�W�I ud�!�>r������	�3!!�p��}�dg��zvY�ߒ�K��kVC�R���K �J^��O���`6F�8ڢ��*b"��f�Q��W��m���m��O�AU�a�{֟x�LQ�%}�#�"�F�Ym�Kxu?�.���*���yu���@���c���7�VwC������<������A7�34p����@�:^�>����Y�d�):�����0���4����@6��K���.3�;0�4�:���k�o�{���r�6�b,-_Zx�V]\�W<⟜��L
��$�@L��%�IF03,�M�!G�,�~Q����xg^��N1��	�Y���&W��w�-^2�'�g�c��i�Hj?aJ�5Úp��I���AHr���ޣ��\x�����H�K(#@8��1���ml��`�>���D�s`[ʟ�6aC��t#�ֆ)��7�۔�{}'�f^�B�}md��UpS([@x��c�3xd�JӁ�T[h��t ����eḥ�?���r�~��@&��	�w�TU��[��鹭7�*�!�$&��n�n�K�	C0�
M�E�/�m
�_�@�E�������a��֤pD�A�D��C�[��Y?x0*J%�
�=hO}!j��-�|$�`�	���R&s,���Z~���1��wk�=�+�e�-7�0���~��D��b�S��?���22���s8��A�4�U�,�\�
��	��Goer45�ّ��e����ϰa�[uG�q"�=*cx�M����Z�E���V�o�9�f@�n��~��(� �J��R(���q����Uht��/�n�q�����aP�٩���EW�������ڦ�*X����<neyכJq�P���sEK��J^)*v�w��6;1�;W�&9�_T�ғ@�:��X�kb���Pm��;�;oR�uef ׵#��>��RV�fp/��8�������(ih�Rϖ�&@Sq�R>�~��H�π6NΞp�n{ҫ�-#�zƏ]����X�&o���:O�����X��z-$Z���I����枵��0M��j�h8^����A^�u�N�@��2xDח��֍�.�ۈKq�}4o�Kh>�Nʇ㉬��-&�|̆��Q�������,A���6Nm�lsm��\�Q�3'��� �ρXG�{��ٝy�����&���f�n)wx�� ���Je�tş#"\ⰸ`h<��r����2����M�/�������1 �0R���}�'!�|k�3��=܍��oYq�ƪוB|�sT�׾Z@_��Z)	A�P	��2#ѐjoܿ�u7
�{�]��${_X��h���H�l���j Ks�k�7J���ԙ��ق�!�'R+Ǹ^��9;@Cއ�6$u��T�i��a�`v����|U�p�N��Z����A��t������QRI�W��>
-�P/���H��B�)V�G��忛���j1�W�63�D�~	��-a��/*L.o7Fr��T�p�B���������L�D'�4[�
��%C��^��E����8�6N]�샗�p��\f�HQ�o�K\�O'B$ i��N,�2hk�Z.�P���$��H�������W�k�u�"�*�?�q��f)ޙO��P�t�[�1��&(�4�����='��k���żac;���yv���p��:��Ø2LU<�T_�������7�/��y��z� d�E��-L/��(����LT�=�Q�%�8� 6��I]����;D;�X�ƷA���hq��㔺9&Ɲ�f/n��O�vfƮ�_#����z��m�L�	�uw˜}|����=qeZ���9c>��QI����CK�f�]�Z>;����&�X�� '��547z�+���J���B�3�x�x��gIʂ��!�Z�l��M��<b<�Q{ғ �P �0L��)̨�/�9�2�⻍y�y|}.a����>�E��&����H]�'�r�����=LiD&���ֱƼH��}�|1�c���x��~ �.H3��;X-�3�J���d�YW���<^��`��;�J=a��n��>���5y@�����c��,��J��!��\��C]��5��J�Ā�`?�`��	e����E���>i�16����1h�<q@\�E�:k�"��ٶ����|yy[^�7� n���|�ܝlO�9��_�@�#���K2�.���#{WKN����-d[$�v.��ǀqK�nLZ8涚J�������-�Y
�Q��*'� �,/�1 U�	fRh��m@\��_�U��}$R3���NP�Q��lV��!4Q��ࣙ���;���ߠ	Ϙ!� ���^`0�T�a��I����db�!PyP�� �t!�0�H�\q%�=M���g��_��GO�Z���zZ�I�f�	�,����Rg��%��Ջ'u���,�0j����͇f���O�8S�VZD�i��yB���ry3�ֳg���m�gtϽ�a8̾�Z�'�-�y�,����Jr$|����k�5��X�#R%/�`��j��ͫ�)>�B""��X�x0'�E���`-&�T��� >�#�G/Y)����	5-(��u��v��������>0�/�R�^�����{A��;D\u�*	�!8��"�Ŷ��?4�;��]|��6�(�
�`�`��nȩ�e=%�w��s�~�h�����5���W��m�ҢO�$��_9E8o*xŦ���{�|K󵬌���#7j5��(�=�w��`�n�;�=����w#��G��B��E�#}����P��d|~��.�����}�c�}	2�~/��`��|ݩ�.0��{õ�r)�g��~-T�fhե�8���z��!Ԯ3��]�d4��%���K0T��6������z&~���H�I�^i��ȘZZ8�����Ƀ%�����O��)��/�5qT���gۖ]6t�4���
d26��P�is#�U:�����e��y���!!����w�i��1�?���V8�|�_ڢk
၀��]��O1V��?z�ʰ����xǽo�1?�N|cs�/�K�e�Bը.�{���{K#itt��!�2..�+��gD������w���oW�5|��od�������f�K�q�>�2�^R��f��J)�j/T�Ĳ�,�����xz=!�:��� A���/������u� YH�;f��4�6�;"!����ׯ��Ĵ�K�W޷��*��)i:�W��W5�hY�����n���5���hLP��/(/��i�9�`�u�%�(*��fzO�z:k�nݑ8���}qS�E)Č�/$T�o_�4����5�Ek\����pr������Ȫ#��@PK��P"7�f��<2gbX�z�ЬU�~�`���~��4�z��\���mY>��ߝ����n�3�8�����.B���Բ�k7�QԵ��v��P��_іFPh��Ty�@��T�֓��[��mY�S8�ʑL�fXa�/�9ɴ��Vat��j'�l>	7�N;��"�|:��bk��e��ۂ, ��ɸ���\9�e);�vB��0L�i���P1��P/XgA�#��D�9g��v/����h߀�]pA������,��nN��Л�c��̨$//�h	�o� 醟��]cjca�+��a� �K�$������s-sc@D&�*��j�B����l�\��x^S7����m�����5��sD�XdwMH�=}�f������HY��D����$��]�=�'�_�b�ƴ��Wg����I0�V<\"V�C�f�d��FU�&i�8S����'�c�.�E�ٲ�nC�$�޻��¿��T���؍B|��ۓZqO�T���z��<S�6��,��釦y�+����>�
O�ɬ`6�G��ٝ����� 9,�!2���S72���]�"xe��s*[�a�/�g��G�VP�����O ��sĊ#���3����̅��#��	Ai�0�ݘBd>uc�P��դ�f`?�E�!0��n�,��d5n���.�S��qV��A�}mN5H���6v�{i"�*&�*���y�ƈH ��Y�����ď�8l$���]�:
���NK�[�v�9�x[�(�#�?����3���o�f�b�+>��1��m����C�H*��a��R��h3f��'�8�9���-<��Or	�U#�&|z���s;��y�k��1����ӊp��E�]J����� ޗ�?���hL�J7 `�����
��I���&�~[S�u�Jf��[��n#�)�J���Ԝ�dp�'84���PF��Ȁ�^(��^��w�KӿXUO̧y�d��,:�f 4(���n�@\B D����-��̦� ��~ѣl��<s.Ч���#KD���LCFE?�X���u�ʬC��-�����j�]��9j��+�NvL;�sΉ���_}ҹ��,�=Y���Y�.�y�C]8���a�jN�L���a G�:j�`P-x�VRyJ�j���Рm��7F��g��	2�g/|���f����G4��mb�	�H� PD����@�9����BӒ�@1���n%���������bQ!�D��ϸ�lʋ��Ge5�u�]�8kV����bDK�r�U�6��h�����E�s�Ԟ�7�h�|�u�@-�\Xq0�s ⢴��
�T����'�.�q
�6�?��7��$؁� ��=���	���u �&��F
�X	 ?Q��)1u����c�!�V):g�Ũ���>�[���M������JJb�� Z���?Bu��C�8�������RԈ�����L	ԴD��4�#~��}����NP����-E��G�798�n���4X˻is�0O�FrW|��K�aXl	���,RpR>��������	MIT�c{1+_%C����͟q�#-����I��#r!5O��\Fy�IԷA��� �Ƽi��@5ft&.tj܇0	���i��H$
�el�y�$	fc��w���n��DE�#:���N��N��c����ސ�# ͵�i	9�vp���6�mLH݁E�d~E�d���jI�Yq��d���V���ߝ�߯e���`������"g�|��+�����͚�!�c1֡�&5�/�(sph&Ht��[�
���j|`Kf��Ȝ�Ķ�~2�qD���$���L�s�i���Z�VƁ:�X�Pqʹ+��&�Jƀ2q��{��D]4����w��2��rz�7˙	��{gG�J@M$��O�8~�|o��?��%�
�A�Z��0���b:���P3��8d�>�!
���bi��8a���7ҿ����*d�@)إ5�
X�<n\��#F[�O(+[���F��ۦf�u��#\���DnU$��>� �g-3�-�t����I��.��۳x�#���v5�ԩ1�����`[���=絛8�
*J����K�0���n���o�{�k��?��m��hj	̶��[����|͢i���)N�� P�f�?!4��Z�٧�e��*��o����E7a;�!���)��娉51|�b�	�����3�o����N���}B���V}�7��>�b�uQĪ��{U��a.��O}T��Lq�5�SA�ْ%����\��Ӗ�ч�u|���]7|!�t�z�5G%�SY�Ě\E�.3����e��|��%���B�2�&Vg$��w�с���Hs`G�i�fNG b���¹ѕa�v���q��� ��١�$ �3ODF��+�ԑ�	F�t.PaNg<�-�=v�K��6[Hni�u�̾��z;�m���҂8"{���ɢ���*}Č�Wdk��7B�����3�L�Uv���a_��B�)��k�0si]�LΥ������=��Tj�@�zH�Q�n'id3�Ĳ���'���K�q�v�$�����>C q*M.R�75�jx{��!G���i���>��u�ə��i��Q�\'s�GR�Z�:��[��K�m+bb�M��o�Cn�)x��ѵ��[Ժ��{g�1�`��15� ��|Y��;�O2� �Z����0c�cA�Yn��0����\E�Jh
��vJ����?���3�x�yEfD�T�3Gx�ە���D�]����6]o3�q'��*J�d�}�P�v�vxd�n�ݺ`,p��/�?|"/��<�mQ��qR{.�r�m����z[a�z����`����ה��j�g��`x3�����k�[
B���,�]]@x����bc���/a����o�)��mz��A���5���B��&;ܩ� �p���Z
�(���Ձ��G]&{�@de�y���je�%B���,�Զ��e-����9zc,�3_F�VD��jA������̄���������mU����9GW��c@~��Nk>˖&:�5��*�D�����y(ҥd�[�Pʒy#�l�jj��������#VݱخoY�c�0R�U��*�p.��#������勃��^��<�Nk%VP�����P�9uؕ�tg���qªj�5t�}V�Df�O��y��%
��[����ZJ���=%8�2�Fq�ct�/�҇h^D��9�ͻ���s��돲]}r���� ы4p)�rE+��%�$j�VOJ}1���ڬs$-�C2Q�K����'h��N�����]��[����WϸJ���n>��I�'k>�}{���d6q�6����qma?�Eؐ{��?��-&��mT�����oŘ��y�Fwdܤ���,�m`F�}��C�9B��޳����^C�R�V��Ct����阻��.�\���4�d�^��Ua�ɚ`�r�d�pj��Ț�.�s�g���n��}�j�DE�&<�Ł�$jx���qj�����V�ޢ�`D #�Tk��1X�c���7��R� ����yA�)(��u�RC����8�S�r�� �!=�9�J�#E��~.lſ^��Ing�����k7��Mb�ӫ����.���]��bq�[�ɥ
�D�#��9��l���gE�!Z�V!6pH���X��Z��m��M�~�>�Eí��ρڭ�:�cH�/����a��[��J�d�"�p��:�.zH���P���ܞ+�6"=6X*�A���w��Ʒ�#Ci���UѭY#����'���*��Vp;^!ڙJ3Ŋ
��^�`d}ewR>+k��I�9:��i,��^ȅ��o4Z i�#S_����(�I7��:`?�f]�ͻ[1.���͈��������7����}������D���7VI��~iVH� -�������S�]qZL�3PA��s���Eb���!�|$а�2��Z���k���?,����V���ó�^�eAC�%Bϡ�o��whi|v�ع�ELKrRQ��.¤�j�9l�pF����=.4�yOD()�#��%h������ՙe��I�7���-fR�QOC�&.o�,L�ӧ.�|�@9�j��y��#�P-Q�A
R�^nv���o�u����p���(��y�8��>l����[^�`GT�@k]�zu6��� ݉	�:�W���V
�6����а�p�J��<,a���a�j7a�;_��Wm�`�,VG�;�X��r�Ie3�oS��b�sV�I�t�T-����Z��AwKg/�8�la�;H:�%���r'���&��E�[q϶e����Xܴ�i-W��YT���-p��;�;`���sy#�-�?�ͤk��ؼ��<��a8�M���,��q�<8f+ݽZ�����I���T�ÃlԖ�������=5V��J�A=~0����p�J����kE{BϜZ֖��1w��xz�<4���T�y�ܓ\���!X�)-��}� ��-Ν�CH��,��4�߳�W�RO*����R�ORX #������F�#��~ӿPk�"m���7j:|w�
+�%�Kd��4�%�x���O����z�cM�A0|�.�d�����tM]�'p��y)[Lo�����ڠ/��2����s2y�cKxB�Pz�ƴ�7p���gʕ����>s3x�զ^��̼�D�EjЗ��IFJ���!���o{5��%S-�6$�P����d��ICF����m��]cL������2��O՚�!��S�d�Md���m�qe��0�S'�Y:�.��O��_�;�������v�"��m��ɼ~Q"pЋo16(��n���8����0��ܴ ���e����%��O��l����Ii*��S2o�&�����c3�+��UCnm����_-�_S�F,��l�!�*A���4��9�v�ʌH�2��Dtڽ���~K��xz�N��,(&�}_����$��)�0��W��-	g�����:`@�ǀq-�f��tX�H!�Sg41�5Ea5�{#M�xm�t����8L��Ʌ�r��"-���� ���1���u�ϭ.��63^Ȭ��&! k=e��R����*¯v�K���\_��"��?{N"%�;/��|�m�K��v����]�dV���r�@84@F�a�F
ץ�.e�%�j���ִ雰ZϤ:8��N$��2�m�:뎶�R|�l*V -�q�x*x<p�؋k�6x�\��koO"Zp�b��Ti�˪��Mu3�'r)�2LӇ�(?�3�w��IV�T�c�d�:����m��˰$��%ûP��)�?�bv����~�c�s�o�<g&�/��Fႛ�Q'JA�n�};J�D	�~�rb?Rf1?^��%V$ωn0B�B�t��Y��V�n���~w�K�<�]S��w�=�`��M|�������1]e�j-P�S��<7t�a	�g?�\�0� �
�e,���#?�����/e��DWK�v���T�>�oNe�2���Z��5*��<�'ȧ�f` ���\�18���xT����>%�6�4�]	�f�ӽ�O�4�������W����^���_�\Qu�c���fA���,��Q�����2�
K&ƴ#�e���>J�%胀����iC�O3����|�lƗ|��T.�m>+`>�}T��6e/���e& �)��d/�}��Ħ�3ΰS[�u�[�m\�c��_��v?5M�C�-��JAAc����q����!FC� ��=�Θ;�H��iU�ۿ᯲���M�>b���X	Q��yXdg5������:A�}��ì��V�+{<��Fo��q}!<#]7�[h�0焄a���혥����(��iK7eeYTO��UN��	�J>�E����*5!C�I8�pd�)��(�w>�7Y��\���^�S �	�C��6_q��(jr��U�!�vjҁ^��{�1�X`#F.w���������Zi��v\�H�jX�"�o(.��2�Ėh�љ�N�k�2�H�~�2�wzC�{h�����yY�(e�Y�M�S����u>����ȂC�;[#b�A�����q>9�$܋6��LA�H���6�<�2�D�x'���^���Mo����+�_>R�	> aC�x)nx@�m�)�Ȩ��O���7��=��jz�e}
|e.�`�%k��e��?�S�^M��E=Kd��6Y_�1.�?�%d�E��AJά38�b�ٿ���X걤��A>�?�k�3K׼l�z��8*HY�i�.V�!��� t%�����(�w�q����y�"�����!}�`t&"x
�����[�h�6V�@�?�u�u��CP #ѧJ�3��%B�-���-ڡc��7��<����z򫦚Ӯ���o<wp��=g�R���`;�
x�-��"�s�j3�s�P�rA �����啼_4/G��͊��}5(�ҭqp�<k�8�+O�N�!5CWE�L LT���vH�[n#ž��ҋ7X�}8T�T���b��v�5KB�-�����te�$��"?9]0�GXI���{,��B�Vl�d#;�⃁��0?�]X����@���Ԩt�g�)���
ב���qw��rA�XnYcU��< x�JE����ޭAzX��&)�z�&�]6߲u��!��ݢ�����Fb�%˳Hp?Cُ~\xfǱ��l��擡Lr l��'�!Xk\f.��l���k�4~!b�m}��7��Q9�满���_�׊7��x�*��c%���6�
��$o�k��	;Ye�Cy6b�輑�(I6�ג��'���s������z��-P
G�S[�?d���<��v%����!+KF�	H����V/㼊s#���X@C�v��N���+��֝K��h%�R_�[�
Z���z�3><a�U2ϑ�D��H=
�Q" �����j��n�~��g�j�b9�;0Љ��>���N�d_��8��Sa��ͽ��Ru���`n�*��wP�3��g�|�I���!
�}�gU�i�Pז|�Dqq�y�	�vh�0Z.�ҡ+���-V��|��^��cH�n�9P��|��bȑp���geR&�`x�Ϋ0�2�+�#n~̂epr�>�ɾ�q�"��\0���Nb4i�(�g|�á�H�����(����_2(ɸ�z�Y"ợ*���Ds9��b�ъ�Tx֚1��)�s-�
Ex�����ޘ����
��g��t`��m�r�?��!6�o`f�E�?s#Yآ)U��K}�d�ݕk9�
�f4]zh���-b���3�=u��KG�/un�wN��Qd5?��$`Q�'G�5�d��7
���K��4���c � [��(���V��m@η�����9�(��J��!�=Tv�;ZgٓQ������(J:���.QaG��l���D�Xk�9��2	](�)����aN�@PUF�ګkM��cQYW6�y�� �1B{�>��~�0Fҝ���;�����
�[w�b�n���R࠷�E�`���ӻ��B�� ��iE�6G�X��[�r�LFz��
���n�56��h;�|�"..�o�A���m�~�gl�w��	8£�m-�ǌ^�w��u�VS�?�동%��TNIi��b@����6*����ǖmO���h#�^��o�X�c�@cK�9���{�Q�;�ȱ�����n�s9o��!�)WG��Ë7������Y%�;�8I�/^Nu�׈�����A2-��νTδ�1V��a���p�]'+��K
��0L��	f!�Iw[�����n�NHa�T%n�K�G8�r�<���K��N��b�����}��[�j��� �'j����"x�3!ФV#���}����׃��c�J/=ĵg�;@�<��z.ʒ���s��k���,�JH*XzA�6[��8k�x.d��9�}�|���ʣ,Y*Fxw��kL����5�K�i��I4��/g����lH�wK+�j�|Ts�̊�5�q��ᯞK�;�Ι���P>*�`mh��6��y'�y����_������_e��u@q5,���R�f��g�- D
!�M�!lS�/@��.S~���M��6�ީ��� K� Y򻆲j�'�`��9k�n��;<Q�$R�/���e��-#�M�`ϏTKN���oL�
��S^�	��B=�L�`v��J<Y(��7骓��z1|^����ڈ���5T�B�����ʻ���4��!~�E�U�i�؍���h'����>@�sF�A�����-�`r�;�"��½��5��(�)�!=$�����u���uje��$Zi�ע�-(b������TP���N���Ũ����<0�@�Z@Y�����R�W@��@-���_w�ϩ|���3�g �#�L���������p��<�IJ1T��+rrJ�Fx���Q��T�:PBH�}o`�w�C�|�����@Y~��*w��-��).�IY���9�}�o�����΢zL:��Rv�_	�ε�L�p|0��pS3[ӕb�.H�:�? Fg�N��o9a���1���C�*$L�Eϡ�!s�]S1�F�ƨ?�e�m���a��R�KE7W�ي�I�_�e�pЫ�6���`�����h��V���9&0w�=*r4<c'����â	-�@jP���AG�0���c����=h���Q%���Г9����~7���'ç��L3�J""��)E#)itm�O���C�F�[����ou}���~)�<�"�a���e� `hqR�}��x`�8G�wq��(4pNK"q�|���^Uf�Z��%�D�7<b��r�pΨ��r��Ϥ�~Y�Mo�:��[������'5�,�������|�A��fH�ׁ�L��*��Z..���^�f�zn�{9�/�N8�K"|E��I�O��������dC��- f����s�>n�x\T5�J�~�3%'�(SU�nşs]�H�x<B�sV{jO�M��Z8<�2J�c�bm �GDx��vL���t>u٪�즺�-Tj�vA��*c ���#P��ٹևe4���_�p�ǃ��x���.듰�<'�vVr&���o�#q�D�<��.��/���	�y%O��}�A�W�_m)0�JDAv~���W���t�A�`�z�`T+�ؗ�&�]�;,?g�+?�EO��Bl��2��N 10cC"1 �I$�� �5�Զ8������ڼ`��"��2/� X�Yq;���1�HD����Zaӵ� �Aro���/�l����`A�;�'��c�Cx�ь�ϒ�!�Fc�PQ/�MN#�u�������!�����D��gx���7p9�{2~L3�kdZ��[Q.A�S��ڐN�!��s+��=l�6��5_��C�Y��I2�YZi���KG�R4�x�T���⛊a�ħ�U��'�����d�	%�i`_����_��YK7��+�k��g�s�)�CT�����;+8&Y.p��nP��%Ft�8��0~4="��IK�*;@:�l�ʈ.$D�D��4(*��4����9�!��(��:yƋ����7>�L߂�O3�E�����v��5�����d�R��Qי�(rØ���{y׫ؽ�a�D9�@�R�n� i�G��F��e�T��� ��{!;@_ҥU�`��8�z�=bݼ��U�0�0uO��J���UP�U�$��v���XW�9�T�m`��.���RM�/uBK%����w魳�~�Y5i����G��È��@L��u�d�4J�^n:�E��wkp0B<���zD���C7o��"B�Ƀ�߄w������;^�6Z,B�v����W�`]��/Sl|~
��n^�$֎مZ��%"+xӇd:8H��ߺ�*i�m�Ⱦ<���_���'0$�!+l&fh4Q��C���}��>r�:y9��ӗ8�K�@>��m��� ƣԓ�ݮ��_k��o�Y�{�YT�<~R;7c�/r�U��W~�����mEѹ���BfM��T�qT\�!�b�/HY1����	<9����B��S�@+���W@U
��T�%�VKq���"���BL/���M50�D�����A�,�b�9���05�/ݕ�ot��A�2q�z�p��s�>s�UF},n�O�K�j��-��v�1�Ux���#�!z"��"�nɥ�A	�*�0�ރ|;E6�8�ZY!I.�W%��ߕ�z\�t���dXD� �wf�\�]�z�j�Mpk������gd�;j�Eԃ��/�;c���%vE �W3�4����-�T��|_�1��/�zp��Z;� !и�7afaj���[.�ow�Z��֣ZwR�4��w8&��{���V\�c�0�Ua��>k���$�IƩ��Z�:�XH���G�9��z��(KC���~U1�v1I=|�Τ(_IwM� �B;�8���>�wѧ(C�P,���QuH�k����6���+�c;��X(�J����4���K��ޝ\K����F����QY���T��Ɩ(��)�#������f�v!��	��c�-�W�}������>�H�z'���,�W�ReX���x!�FN�"q�>ڽ�ʳ��̻�_�����7�RВ��|��4*Z�T*	6�����Y]¸:�*�6��Z�%7�%�v�2P0��	���4 �ȈA�
�iy��V:�|�������$[龠[L������l���vM�bur�/�?H=Sz���fɩ��զ��"ؙ �WzBО��؛l�_=����_n],��Q$)IAuF<�l�X���8�5�iN3�=�2�iTИbb��&"�3�0޺��ʉ>��b�[3}��d��&"��5�V{P(s�0�Dzv�V�p�l��Ax����iؔ =�r�0��rbEu;��ކq��W�H��T��#�q���]��?��O����C���#���?�l���5m}�Q��o�N�rCe6F��s��&��~͍g�)�4�0�O'�X�VcM!���}V@�4'���y�w��r��}��BS�Q_�*ݟ^��H
`~`UZ��Y�2���J"$�B9�.��a�o[�梮ʀ[�Pik�j���V�"��U\�V��;�Ih*�r�%נ��4K�߾dI)��$�߲�� H������v��'X�u&F@���ԣI�+3F����vf��S�y1o+^M�#zw+�э�����#��
EgW冷��`D�"�x�~��������I��J&;�.ڒ���́���R�x����XH�i�^K�1�+�B�G�[����G{CdT�����xF�e��2'�0�\�$�"��R�C��8�
���7-O���\�'�����.R��F���j�,!�:� m�u�v��e�����l���bm�ШCj��I^���^��}ap��:�-����t�P���Ǩ�p�q��
pӦ��+����:)<-�����s�͏,	���g�����������MG ��~wW;�:����|�&��� l�B��PB�*{�u��ݞ�*r�M`)���){���5��3e��]���v#$L���z�7Y+�B�G*����$��ل��܉�Cѫ+�p�R�ń����A��X��s�@�Q���̈́��W;nU �Lډo�g?;��<*S�3p^���B�]PAJx��+?Tk��
�� A�+�9w�������f 4Bx15���(^=�c�@�4eU�me�Sod��[�e�xzM��+:n������Ƶ��\"P��'Ȣ~�f�����hԌf�iC�k#}�竵��-�D�c,�<����7)?9�J�9	�}A��b\�7�����J �7���->��!$/�L�'�4t��a��$��v&`n�;tfG�Xݜ�2OL�l�����9�._�x�)�h9#Cay�.h��$�Tq֝r`��v����x�
<������?���sLЄ3��zvV�� 
���W=��a���ӱ̣[ȁm�=g	M�~K�ɥ�.��m�]�x|�
���Ր
��/��,x]xl5!����b�E[� )XT�Q�A@�p�k�s����E��֫:��}���AA�4U.��Q��SH9{L�{�يƌ{b@|����2��$�jڟ���[��.]���ÌgX"y�"���Wo�r��/�^GE����P�A3�l���h�3���0W|s��\%�]��|�Q���4hDrT[I�U�Ѐ���M�ړ��C�l�$H[L4ju\���6m�C��!_襪B� i�oiV�U���m!�$�*�RV�hY'4|��� ����Z&����ڭ{�%H��L�7^綼<�b��&FBB��)ߖ¼٥2�";a�v__�k'��'9%�����2>:���GK��.���b�P�`�.T&V����7]���FT������ɸnr���A��^�Y~�j�7���ތ< ��Bf�c��P6�������I��,1���g~G^�qծ6|��C�	�8��)>��Y�Z�*�	:_
;i�ydšg6��A�1�jJ�M�7��0%�\���@6\Mk_sW4r~ˁ��ar�U�DX���c0�A�*۝]��]���Uaq��m�0�A��3�4�-r��� ���f��9C��;�v�w�'��Cs� yM���3酣k��.�O�F�9d�l�z�P�X�F�U`<����� 59�D�5�%H	�!�4
c"����,N�]5���BY�3�DsD� 82�s�$��ɒ���5�6j
8��������/���f��j/~���>E�y��~m����#��h2Sp�ߵ"��Y�=MsW1`����IMc�ś�{D�l�L���t��}��	�墜�-Qh�=���l|H��B��)�I8�19��ο��U��V��A]{u���2�5�!fs�)U�k�ld��T!I�e= �^��{S�s�y7�Ѭu�B����3}rxo�Xs����ĳ�L��WI�8�/3����l�1I����`l_�x.M��!M[�A/���X���ym���{_�`��?
�6�M�m��N;as�qJ�@��	�2}AXF���ڶV�s�7?=��V"�d#c��T5��?to>sFT����X1�(���y7:�1�՚`C��\�'l����ÓE�34'������:8� �M�`�'��B�@��;9���p�-��e�1`n�?W�-�*l$��ڮ��Z#��̧��v`н8��V��3W��Ao%&�F��l&�f`��-��c{B��V�x:�rc�@s��C�������I�������cD�g����I���@��C�&~�=cū><k���Hو�OEJ�|zczn���dZ�b3:���A�n�Pv��4�s�S%�"Q2Ȅˈ:�Bx��8���^�{�Q;J�4��pH1īK	���a�Alr)V�)| ���GF;����O�);Ͷ��_)�}e.��U��z�P�E�;6���zg1F6Ț�ȃe����Bgf<��Q;�\o��zSl'H�"[4���2,M��J-%;�I����pH��M�2��)b9+P�e	��pA�XS�7���|�������LU�5����|�ۻ�&�N����\Y�i���6ö9���j׸ �Ϙ���`t��o)��~��^1�b�
�'�qʐ/-'D�t\h���]�`�16���qz6?����9�%\�%���CNd̤ߨ� ����vo>ZOq��ϸX�]��W���/�������މ���e8�e����������^�U�H���輣�"h�^�e6��l&1`Ap�����C�)��{k�K���Gې�j
���e:~��5���ցiYs�:��Y?�8p��:�;�����6{���Rv�;(��K�'���
a�����8�g }_7GSy)�.Ӹ�m��Lb��Bk���ג��9�?�yw�9������G�o�D���J݉�9��h΍v�%�I�1YܕfFŰ'�oŝ�V6�g�^Ț�
}uf�(����*�L_�w��5U�'�Rp7#}��3�+�j�xP��z��BK���y>�ɏq1h>�F��Uυ���k���̡�ݑ�z�X-��{Wҧ]�g��O]���c!��""*���e6vC?�L�g�G)���C�H����f)P���F����2��jjϳ�t׸�%{��ѵ?�@�)�?5�i�^mV퉞ƶLBFԮ�CQα�h��ЖM�&�|�Di���`��J��D�9N��&ͫ�ב�%�����ˉwW���c�ׁ��u^�5ўl��wѾ�~�smmF� Dr�R?�J�W��H;>��&Z����!�bg����� NT���;ܼēzls8$6���T���z�Ц��(U��ꁎі�^\��p�G}-l2-oZ8���I�$&�0O�4�X]�}Ut��\����)�`�?,paR"v&���sV�Du�䆲z��"Qo�H	;cq�(����N<������I����:WK��h[���L{u�s1�����|E�r�\*̊_��+��S�^�~������@5Ur�h���ҪW&�T$�&��0�H��YG�XҶ6t�'FId�r'�Mi6����g_� (`�G�Z20p����27N�;�Ό:=�5��G%:���5�=��+A?!ZV�?���1a�xY�u[X����_�}��v����;)L8��Īpί����:��#���<D��q�LO�U�̷_�D��}~��EBv���)��-=ev����_�꼢�X���m)�ψ��8�m�AVKō����� r�>�%��C[�\��P$�^8M}��q�`�����K��No�;�v�6~,��$E��I��;��;��2C{t����$|I%w�њ�^0�]�Ʉ)����� ɑ����$\3t|�-��0/��+�bUt�-&��ܤs�[�D�-��囂��o<��Ň*z�ByO���s3s �A:=Y�ze����g�ߙ$��U��{�,�W�:KjW�ƫ�عpo$P?��p�U~<r��N��"io<��M�2���A>5� �6;"�ߘ�(�4P��^~`*���{g��������J�w���%�L�yj�&�n�BdHw�ߕu���N�;����`課���M=n'LK���n����a��S�dnV�-�n�6��=c���2WNx�4��$�г'�nn�Di��UR)DMĠ���G�U�}7>%-��%�{ɻ�=���z[xIҜ���,����02�'E���pnPS����5��"�Z��ylL|ĭYSkr�,�,�&Oo�"	#��Lihը����a��� mm���)}���-�(ō-�.��K@d/���v��H☷aQoKN��ԃ�����[!j��$�c�������<D��*w[Y��/�¸o��]y�~�	�T0J�sI�q�g���S"\Q��J��囂�r:	��LӃ��h[ g���<{�ao�_���-��o5.P�<Dڴ��#��.Jtsx�4��;��̓��b���p.���u�w�f�`��_bf=�^�E������k:)Gh�� Ѡng���}���W&gE(MiB�#������MwN���P�eCӥR0h7B+ʴkq����(����w��B��d�_VB>�+��d�I/F,�5D
�2ë���I��м��%VbVxM�E���T�Ь���D2'm�@�,�\%�!FP���`��E�Dv�-:I�x�R`�0�����@��LT���
�~\��kkg���">�`LM��q�
".������-ܲDwh��U�l}(Q1��/��3ĮK�yb�|7�k�����`ǚ���՚��+�f��@,��|�f�\��E���� ���8����@i]��FAJ�ܗ��Di9}�˘��Vv�H)�D��)��,6�� �U~m'(Q���É��(�%�1$�]�hgG�~8������R��J��o8|�;S�#��Ge�~��qP�;��%�����S>��Jo�9�P��pE��\�e�HhE�S}�1?M�˹<�<���\-'���l�����z�o�2�Ԭ���<���=Z@������V���H��I�y�q1�fޡ�?,�j��J&��O-ts^2_�	�{.�D���A�: ���=`����0�5�b$�Ⴍr}��xM�R��o8n:@��L9A[J��C�F���߄�����#&J�	�H[��dc|Tu<
N?}ϯڇTB���[L�{Xo��� ������̞���v�zϝ���#Vd�ʞ����%iq�ۘ�[�y��?'�D�W��_~OpaǦ���P>_��Vs�t^0@� "����GҜ����`|~X?�p%�!g.a�ݏ��Dϴ��f�:�� ���l���>��پn����?g뎸f\b�F�]����3���m4�ϕ!��8���J�(�_{��j����0���I�mB$�x�?b9=y�J/��;���p\ߕ�c�ZL�O4�J�H��)��<p��ЄM.�d%u�=�W������0�wj�����<��F'�)!1��HH����5��[�I�b̦]�N� <Ώ>�>ʗ��%�uF�^h8J��#�׸n��v�۰D�D� ����z�>O�=�	X���`�	ljP��u�n��<�f���5�z�	ЫjI���,A�p$T++6�F�~�?����J|y	M��
�H��Pʗb$����΀!�p==/������j�D�x"�\:L@��@K��Hn���ф�V� h�.mdE�����$22���9�#�@ǃ�V"'x㯇�I�|dטR��w;��@�)���ts�ǻ�V|�u�q�\�N劧���A2���vs֏�i��\f�@,�Y0e�����؏U4���׬n-�Ne����L�q�[]T22�(	�d��c�)���X�
�w�G�2�i���$��A�U��ӭ�23�'��{�mf,z��Q�,0������7�I�@M�;M�zuY1�՟<�Gt䮘C�$;�$��t>&��A\D��H��;�j���6�q{��|�0|u>4�P���w[4��,�E�S�bh:��t��$y���)��Q,pM������[��F����[�깚�Xy(�L�����9���cP�����R��@���~��Ƈ
�i��"n�p������;K-��i�U�6��9s���/�l��eb���HFvӤ�.3��C��*�t�$$�K�C6B�0f�CJ=�o����)�\�|���hy���8�E�O/<y�/3M���s]=';��ۃ�>'��~�[�Ac:��_�
[\V[;��U&C�ޟN3n���@t��.&��H��lb�Uxu#�S�������E��S�_u?̨I�?�^ ��%�V�I5�n�A������9���l�*5���̬QA�N��R��l����� �%h�W��2��e�K}z���8\���%v�5�ʎ�b�TO�l xJfg&�����5v j��s�m�b`�V�����y /�v��?D��&�iԽfX'!!�d<��S͎\�����j���-���J����E�EX��g�	8��	-�W(�6旨��{يS��#�DQ�c�I��,�k�}�n�EYN�g�0&<6y�BL�k9TY��������mư+��Pv*��_�]Rʪ5���T�>^	;���ǆ�4��=V~M{@�9�~�C�QF�0�MܿH� J	m��h�ƕ�t�սk�@���xb�vW|�OhP%81����^������%��7Cݼ�!���z�<���$-��-��5%�뿌�`K*IF�*�JSR��J�x�\��k���^��&����^�w!H�����]����@~�W���@�_p#k�8�������4cs�����~�tW��j/��,�5��V�q��L�����B�П�ͦ&�pf�D�B%�.��V���	��#q����=� �fr9{�B�Y?��E��/�����r/頃F�	bSL,�_�tx"��,��"|Ͽ��m�ҳ-���&E����������СK�\(�>��{ڊ���F쐮,�} $ףA��ح��O�����|-�76��N�{�}�FI(��K�>��l��!��"���~&3;��(�皇��&��7�B��$�My��{���BP֫�@�������>�rQ�2��Gq8���b4ô����W���E�߶!Y���D��"%�T���c���5kzG�):	K�ք�T�@/�Uk���_vp����15^�v�-��RL��{�%X�ք��宆�M��g�~4��L��cq��}6�<��,�8�d9��k:��9|(D�Lo�7�vhJ<�z������gESE,��E�t�v����La�'�R:Cm8��^"�=�9c5?����v�c~���lFs^9���#�qv����]]M���sX���H�÷d&�>"�����L^�2��I|���3x�|���S�����2��q �Q��\z���z[�������`՗e7x.��92�����:45~[�2�W]g��v�������pݏg��sS�-,����;�ڧe�I�4�4�>#�x�s�	��m-�j����h�{L�#���3�9��S����0E���Z�_д�0�q�\��Х��쉢_����ԈF�p�A�m"��@7�i ���{-m^:~�
'����Z�Xk6Z��I�����9��Ҝ4xC�Ɵ�i��ӽ0omaB-}Y�Q�+
�8���Ka��ɽ ���28㵹�ʃ]fwF�*HyE:�P�9R�����;�^5Y���7�v@����.Q.za��p`�8!�Qw`Z6��a^��
�<��.���7�� �pu���`�����Zၥذ�fOL�Q���VH;|�����. Q@Ξ�9�\�*,�_�� �y�5��!L/�("�,m�懤���z��
Oy�oU���NpH-�D58�A�.��!��.��'D���:0`"�B��up9Q���T��b�_���Ԇ�g�.f7�T�C�w�3��ɔctzg����20�k�?zci��ʷ�r�w4B��rڟE *jז�w�saZv��U܃��(Vi��n��sޢ��$�	�K�+ �=�ꄪ�!:'�"����lZ���`��j>g�n�k�=`�r�T�� ���#_ �Y��;��:F%y��0w�@�q
�{�:�%�/�M����Q�=7L������IJ.�!ϽU���R��eO��v�+-*Lŭ#�)��3Gh-�����p1}�܋�᱁}UC�˪7�]����RBFR,9�xq��)��H��΄^������pK��H���h7-{��lkz�!�|�O!���I�%9�6"�y�RǟЁ	�\ ��2�A���t�����֙ݬ��A�K�a;}�#��ִ��R ��t�_5۶^Ź����P3?�z17�������AE�rŘN��|ݮ��:p�t1�D%�=H�b��>���T�(������<z�!P�J%��0W&e�V���)0ۛkf�~!�.3&+���a��v���؏Ή�mS�����yޛ��s2(o��!	! r�-���[�Ώ��Q�f�
y���ٸw�&`A bl)�42�O����Z�]0G�Q	}x��2`��؈#��gb�~��W8�+*�t�
������xz�_�b_:,
,c�P��@P��^搅��9���p��C~ �|�ᘹ��6%*ꔏ��p�9E��L7�{���*Ɩj�b�������a��ѷ�F�G�L�����1���`�_]���C��s�g��3�k��K0v5ʚ�X�~�F[�`ѧ����}������%��B
�p�w�q�)|���)ɭ�g������܄-98("�5�dhZg;2;�L�K�d�9n��Uu8����Г��y��@�S�D�v��[\�*`F�h���/�ŗ��<�\�	��{��9&����[V���V�g�2q�ߑ<G{�-��?��q�2�*�T_'%�6��ZK��di��1 �j,�a&'eh�Ra.wHH�;$����s�!X��U`a:�	���Td��Q�\������@0�G{-�K�\|�.��,r�a�Q�=���i���l���p��A��@�0�z�K�k��U� YD��q�r������o��x�Wߝ���8?o��y^877�>�7V�5<�WPu�M�f�EP:�:x��4>���\�u�t�)��l�~k�SC�ኧ�͌Dn|��
���N>�_tG>��g_r=$�
�I��b_:��&��k�5\�������~a(!4���1�-aJ>i��8 ��͍-Jm
-�>���N؋�Feu*x �';��4�/�^b!Y!�����c��(*����=���� � Ϗ��nk��?ޣ�ζ��m�� �E�� �]UamT�hׯ� �$�H�j+=1 ��`n�BE�l4��>x����n��2\���K��>H�������\1|����׍�h��7�߷�b����DD�����12/b��x���쇣���9W��0�/��{�au�?�X��*����7_������n?�����y
��<��|�I�1O����[x&��2��oq�K�lp��esA�`��OJ�H��!�f|~@ -x�<�=�յ7�#�J?���ܦhAe��wXBeV�����n\����R�B�B����QG]���'���/��k�?��n"�usW������.	�1�m���C�6>�K/����rY������̍Arqmu5<�FL��'�����F�	��<�^c`sW�A���p^DF(mF��#�$��������"�|���[�%�Y�р���ud�[�����|T��cpakj�W�ޮ,W~_?��'�~�ٻ���3
2(�~��]���K(�Pv&��ɠ�Z1���"|��a��_8��|�#����v=i^� #��Zomj?<�i�X��%���I5���rKꖇ�� �߻��TL��-��5���.�Mz!���L,���
v�?�G�y��З��?��N�H,�yX��P�NZhh��H��%���W��I9�CB �����璿�-������[�����ƺ�bchiݕ$�z)­R2��Γ4���c�u8�Bi`l����o���Gi�
����ߒ:����[�*����Pz�^�����Hf��V�`��7��:�q�W��X���:���
E���Ob�t
#x^GW��l_F��U#��]k���_�YLlUh �������,��aW���7�N7��a�k�.Vk�f}���`[�V(ڛ�8$8�򈈻{��\"6�jL2f��4Xxo�šerpq�
4���	��-�p�Qq��8��ݣ��l��5v�%�&Lδ5���1K0��q����g1���Qn��B���Ғ1�0�{Mz۲��W
6�m�?-.������A{��+a��́�}�_f;��[ձ�/�4�W�VV��<pLz���teē��BN��ևw��\	c�8F)@z�![Ud��V#�6�c(��*�s��GXq�����H�7�Z=�zZ�'}�RQ�S>나{�J��Ԉ]��=�A�ԵQ�ɛ�Xx�xyɿG!2�L�ߴ��p���*�������/䜸WI�6��}/,��~I��OB{݌,��|����C�&���C���~�\���|>�X	XZ��9X��{#�I�x"��~�8�j�H
1���$�k�L��B�8PS쇱ؔ��(�IP��A_=�zJ���`b��97�� �o��EW���.�TK���)���H*��ȭ��O���d�P�M2��Ԃ��5���x�^�:@�f��ɿ�n1� �����
�A*��5�߂b�nz��j���X�I�F�Aڙ��"����� ��[@��b��Ȳs��}�axn���^ �K[�#Q����%��Ɣ�Pi�q���%��i��'��k[
�T��Ȥ�sf9 �N�]���*�=�8����Y^���Z�Q��a�|��������[��k�rP���>n��Øt�U���������}���DW�H!#�а�nʦs�Eoi��E�,��8���&�D�@�'D2����v�Ղ��;��gQ��zj��	��D=�8E���u4{x����cs����ҮH��w����`�л�l���~����z��dB��Y�)I3�á��B�g�6�hoQң]���\(޻!b�%��͝�ݭ
����3��c�w_�?Չ�G�s�����u��b��G� �=ǘBކ
��yjK��)d�<7����ׂ��p>�66�r˿��zV6k�+��央��Xٗ���k��2�{b���>Ƨ��9�b`zVʋ�+G�1�k��)�
LE��>�!��m���Y��m��,z3��ݤujf�H���%A�^�F������Oj�J�T�95$�B��'_��J˸�3$�w�y�/�~
�ؿ��]�������7(�'�E�ҡ�kI�mw�ퟺ��@
I@O��zp����������S�C��֜}.�ku��Z3@�a��p��~�9#GX�V�B+��w�J��5{©�w�c�����Ll��E����$�X�9�K���ԧlc�
Bx$]�0r�!!}Pȶz-(���R
��ִt��ig,�m�H�b�����l�@�z�1h�6��F���#�9��=�a�d�bw��@��gIw���^����#��� :�����0��;i�E�p��Y�2�(=�b��3���(1�ˉа~C����}��6�@LnTϠMV�D�!6/��� ���:a���:�Z��n�p3��6��Cw�/���ŧ?�2$X~_/�������c�hu-ܨ��9YŐ���xPi��!�#�G��ʹٛ<$,��2���й�C~R�Z�db-����ī~g��m�:L�ĝ�E�c_�b��\�k��)-	��Q֔�����^����yd���Y��(���,x�pԪӧ*��p?K�*�>g�$�`��}Ә�I���5�}"�?u!��q%�������ڔ��#�A|��c!~2����
�5��C�ͼ[U��S��_���[o��y�+}&�׍H�9ٝ��U^Y�z�r�:���G�������K[�F^�]��)T���$z����j�����,��
x���X�gB�as_}J�,��R�n���O��M�qb��H([͊$u��*0���9�ց7G�Pi�h6�L_
��qS��}��X�b-j�m+
�5fL�p�M_�-���G�h/6� ϯ��&��<tEɍY�1o-��/W00��;�d �s��ŀ�9w�c�6�jc�O
_��E�8����F��C ����F�<��V��܎&j��1�0���CK�׭��}�U�]w��b'[y�����X
L��<�1���I8����3Z�,�$�E{���Ц��ŁL��s1�3r�/��%Xү�e�t1z6~���^U��3x��2�f7[4�*[���U�m�?���we���ǎ|7�E�;�)s{�?%b����w;ࠏJ�8)e����Qy���ހ�v�3�ڮ��\9v-M;�mdEۂ0�N9����
�aV�]^��D����]�뇔�Ú��B}�v
h3�t��J��gԋ�N�0Ь7~p����X8 ��I�v���{�x7�4��l�ܯe>އ�u�
ך{���o��[��,���K�5��S��,I�,��#f�%��#�}r�D	�Q�.��N�R�!\��_��L�	�8�m��P+e{�3a	��&)��YA�����R����lY<���^d��*�.s�`(�i ���Xs^����o��v_U���U���
�!z>��l6�[�2}��o�N�t���f���ؠ���ք��e�^��t-���H�<�˛��f��Uge��hK�Ya��!)�1`i>ǥ��%�<�%ɻ����md�Ta�=�*&�m�Ƈ�sٹ��lZ�a��~'0�%�!q���k���1�ۺd����$^��F����1��GI��K�?�ga�f,�D�.�{�=�n���e�T(�,/��^�0������m�C�I��/yu����+�m�;/8dm^�#����b��^�|G�6y�#�E�7N���-�A�:���VԤ��d�;����]r��2a�a�ˏ�C=�SB,n@���'��+�����R��*���S��?��1 ����s��/��r�~��H��������Pށ��!9������mWܑ}�����?iIGp��x"o3��	3��YſOqڒ'n�Ŝ�/�j��%l]�,��|��ɠ�`�ˤ�h�8��3I��5J�<²h	�\Nӝ2E&���N;C>���������Z1+_CN�̟����v�>|�y�Ӎ�;�6�}���*;@����~p�f�J�yS
�|0�y%*44�֬�ϗ p�Ν��1m�5����s��]U���>�!z��F�h{�tc�bb\�H$C��Y��H=[�|U�,+�����̚���]��B!=0B�vv/��\�m�:cD�u1�1y�x V�*D Ni O�E�D��e��Wn��rZ�c�-,fo]�N:�!*��L�벸�{�o�Tj.\����:X�|C����jei=bM)Sk�%Nl4�3���s�����ס�e�<�qAB̶X�պ�� �����ƅ�ţ��p�)��v�9��$f�A�7x�鼻0�����U�}3G���0�a9���Oܻw�a���X�	��
�x�][U喅.�`QEiq!��а����k�u��W[�C,�.�#�a�c~���>�����=�Bkz�Н�ƚz���	��663�N���?��
�s5�D��!<�J@�7��ʖx��z%,�u�-��Q�p�� m���4��Σ��r@��]�h�i�dd6�#~BZ6�[Cǜ��#���I�_O�N�����u'��xi���F�ř��*���ß4!��/������+���͸����UԜ6�˞�v����Зk�IG@g/�:#0c �M��U@�SH/���3٭���Y�fm��7q�Dr7c�@>u��x!x^��;����\���(%$��9V���p��
�sf.��@��+���^K�zh>�	/��/�{�ksݟ�Y�P��$�G��( ��L�.�M�2��fCp2 ��NF��[I�����	-Y��A�\��i��/���X�b���՜[��\��z0���n]s��X�=�S������A��p�	�+Z]��%p�/A0%��]����ਂ��	��Ҭ ��*ɡq���5v�!۔�v㽱ǵP�|C0E=�a�=�~�����������M4*�w��\ӂ(�o��p�nBe��>���z�o�u�c�]2.fX�WKj	��2�׺�������"(!A��Z���f�N�f��_��KƦ?q#{��$K:M�WP�`{%f����	�J4��K��[S��F�?�z�T�a�}0�~ҍ;��B�����"��,��k'L��垌����{����_f��d��#��+9j� �/;�y�|M��h�&M�����Xs�K�䪞���R*0.�:���4�6\I�p��V��ftL�6Y��r﹧KR(#��7��a���ɰ���m��*P|�ıV� jɪ��\�h��+��d�6F�����K��͛E�E=}��X�c/����6dG�crhn�}L��M��ceD�@U�d�wX%a	�ߗ�M�SJ���p%i$�G[HFZ����#I�m�ϲS��4HMa�j���'f�ף��)O~-��'�`W��*�(�^A͋�Ɗ�>�X��`Dj��bo Ȼ�0�O,=�>H^�񀹁���:#bB�k�~0���0xUG3޵�a>&$�)�H&ͰӼ��X�%Q��������z�6�W���ޯ���Po�F�e%:��GH��}�lҨV�w��N~#�Q�vkT�lU��j�G�� Z��/#��5h߯H讓F*G�X6�yQ�o�PfO�#dcixn�0j� �o��_ES�(�^��_hk�6G8�[
��@�2�M�|丒񼟩!�<�=-�c�l	����/b��JMR�[�Vb�m�;t~�E� !�T��S��
��|D8�c}	u.*�=�SL�f��`��@�1�G߿Ol���LC��'֯�� ��w
�j�,8����t m��B��1�ova�"4 |�:M]�mGMcvƯ��\��ék�@ee��Y�ˌB�Q�p�SX��y�A����tP�g
�Yl�J��$�/����YHoG����}s5�H��0�s#��4]�H��h�� �ߢ��ߕB�Gt�t��.(&o�ڪ�c Z�j	o�����dŌ����ƶu��UHde���u^�?�	:�;��<��=���H�,K���Z@�THڸL��{��ǯ\�	Y,nu��|�gc��e�H�b�F�K��@��#�~{RVw��s�؝Gu:|'as�E�����l�n�h���g�a2B{������L��lE}t]־6�Mo��R���݂=�lu(SakQ�o�e�����������Y0T��Oj�r��CFzi<J�nq����{i_�}w�RL�aK@y{���;9�k4�9���Y~��]ЎA��\KE��D�pZtȫ���Q�)T�(�O��Ζí��~���#���M���i2��N��XØT���+[@Z����'��V�_֜�<K@Lm
V�O�n��Y|�̸#�
�U�gb�	3`}<�)D�L���P��MA�&�@q�|q)�c.�L�3��/L�����Ɍ�T�
���'ΰ��	-AK�}Ԝ!�n�/�A/���qnc֔jnX�"Y;̐s�9,Bp���#�T�C�' �(4~�ķJe��N�WG�E�R�bY^�e��.�o��oC�[������mܸ�\�D8��yN�
�K�.�{qji��-{}֕	ucvs����#W�2�E��9c�v$ɐ���d����f'�h�+}�]l�mЖ	�є! 6o\�Oo���	ɉ-�A3�Im
(��3˻~*�+�#�{������]�ě-*��� l�c�O�`����.-)����jQ�B��}�?E���ۅ���(�Ŋu�*�f�Y�k�S�͗Hpg�@��rsx*�UvCwI�R 	�^���E{+�����s���a����[�\y
���#ةYpk�;�|��z3Wd�vW���E[�ӣ�'��"�ܥ����A����n�S���C�θ�mҸ�J`���B~�����a�?�g{?E���㛛�
=	\�.��i䦎�#�}o�l6���Y�;�B�hP�(��r����k'^0��' �w��*a�sʓZuL�8sG��}.���,|�<;n���I��GrE�����j� ��BL��t���ư�(�����y����m�b�� �5)0���]��!o���C$T�p�-\�:4��m��(�o��{�<�����c�ߎW-�
>�}Y@:����m�݀W1ZF|,d������е�/uݟ���G[<w�,gi�R��s�p?�(�OB����i@��N��tW <E���+\E_=����u0H��V-���Eq\v���u0�� ����x��y��iW��9�AއV@�6n��� B�1l���y��
�����Y�<T*��������a��3m�;
�c��Qqz�O��tȾ�c�I<E�1�j�O�r��H;��G��
�B3V�L%���m�T͘(?���F�l�9���,V��@��������۬t�KͰm��Ex^��jŖ4S�r.�~ i�ٸxn����#�C�;���ܚ����ԋ���e��R��r>��݄:M�RB���
��&ЃPn3��0-"���.��ٰ2EȀX���2���k�&͓5 j]-K��z1�0Ϻ?8�*��_��޷�Z���i��P���O�ʒԋXC/�|�����)��V�2��:4T��k��JH ��T4��xl1RX���%���S���B;h���9�&-gp�Q��!K��1}��w�em��0LU��p|��
�k��.�@l�k^9�R#���A9��_
�\n)�#��l�P*�r%�'t��x�nK�<�;���F	����������P�-�v�"-2��	um� � ���/I��f�w�5ZG�P�rI:���+��7!wL�b'�p��a��W�B�l�$'{�j��{�bW��:�/gjm��@$�_>���וf��s���j�
�*�Q8#�`�+��ܪ_��K�Ҁ*u�{x��܇W�_6=�YsH�B0��nyl}�9��-�˦��^hd5s�
�hI��r騷[[�F��S������N����A�N���,WHH&��#��geH{3�w��fGg��o	&�R[wL��pL��<��	�{���6��Y{�h(�k9�λU�v�u�"8�t�ږ�3�%媎`��K˸�rIAs��:b��vx�3�Ț�z!$7�V�D�e=T����n��Ti3��෈J_�7n.�[boS�M�g�$9�`US�?w��R-k!sW�e�f�;�L�NT:�|Cu�
�1���+�M�,P���ē�D����F��X(����� �/�����ҿ(6��)��z-S��L݈�� ���4��e����ET~��o�{rLRɫ������f��9�
����y.�L�n���HHR.������5����ޠ���q�Xy�c
��ѲU��9s͆�d8�܎�C��Rdu#h9�%԰5x�OR.F�|�}l�ߋd���2�n`{�.����$ޠ��nv��3�(�����-Im�3�3�8ʫ��F�yX�#w��O�d��s ;�*��Mm;��oZ���nl5A���^��|�]C�X+�$�m���OLt} �t��4�@�5��s��࣠똅��v�S�Sxb���Fy�8T����Q4�[y���ݶ�M2�2�`���0bC���:�,#�jv͸'=�#������0�S%M������z�LJcB[?`�$�#2j��7�~J��̝�/���J�]��������%l5��|��۠�X&�D?o�T ��ZZ�%��	�wH��)$9mk�y�J��]��<��_�>�,0��aC	є��^I�
������hJk�h�ʂޔ)N�a��2�n����Q̈�Οu*�厨�>j��%=��Q4��[�Ѻ�׀**1�3���<�A1D't7�������Z�q�5飭
�������w �DպH���~@0��?�)�~5�$^�Pe1�D�h���C-�U�)��U�k\e�C[5p3a�M�L���C���8��A��{�U-�U��l~��	����eS>�35@��N��j�[	G���lCɐ~q6Q@'�4��ɫT�4�S��+���[�<���rY�X��9տa�斚��9�hsB����-`y6��}������3�ֽV�K��ػ�rݡ�4u���O�&�Md���a���NQ�qV*f��$�Q��5��N����sO�(�s8OD�Z;�Oos�H��v#���:��v� �W9�qo{]N�Z��\B�[7'�r�!�A�%���*(L��ըAo'�WcHC|��� Se�L�HD=��m:�	�u����� 3�k�j8�R>���Y:g��ڨ�!�C�T��	��B��
Y<5��JJ�����j�u��� �R9�#5	v�-��� �"Sh�s�^���t��<�0\�_��:�)R�������x���Gf�WZ'[t�zЭX��t{5����"��,rn�%I�M��f�@���Rh��Ц�FP�$�w�tӝ�tp��|C��H���s���Αdȩ�T�/���q��Q$��A�z�QL�Y�E��2�����R�G�]�S��;���$IHK���ZşR��X��(��ڎG�)c��O��U,rR�lT�YL^�'8]��XA�U��30 g6���/��v�e;�!ݴ���m������oN���H��rI�Nҝ0��k둈|�.�����&^͜�zUC.�ǷPF؍$�����y3@����� �D�U��:��YĂ�]�y�z��@������yoQ!����N�Z=��gP7�hO;��:�t�JA�߿U���|t��*���r�]Uȿ�#��y/���-H��7w�1�yr��n�}�5��]߫��8�2��v�)��M	̦ _��Vu�P�Qzn�7��D������A�K�Q^4�� fQ#`�{��د,t�< wBθ4s�ĝO�DB�X����h`��CZ8������K)��w99=�v)ok���^����@��-&[�W%�@���~U���z��hf�u�����K\0m����OS�w�5#ݯ	NZ��$��$ż�	��yTK��m��p%�9��'�rg�+#�|��:-�����Q���^B�R���ӕ�ϘJ��[Ҏ��ki+�-�=�Y�=:��TsK��;~�5������Oٸ�_r<�V'���bz<���v ���D��"[��p���"�����'�����j�'?�b�$iJ ߰�@o�R*:)|���@)�;tX�ʾ�Ϸ��_�t~�<����K<غ�[2�g���>����n��q���!#�t6s����sZ���6�#nCYEj�{8#�B���v=��Hz��Z_h��"�}�0jV�5*�PŶ�K���%����b)s�z����i0l�j��yJ�4��=�W�;�K,Ru�|P��[tS�D���̡�M�[�T�Kx�M��p�K�aq!D['2Sd0��m;���o��Y��˨�`��)`�pp����.�Ƌ����6F ��n_�����4��/߼�蒻PR�M���,@��<���|��Վ#�o�&ᎅ{�\���I�D�)ڹ�X��h_(砢Po��qT;; 2��^���{�H�2c$hs�u�a��;�ۢj�1ɪ<k�b�ĸ��I�^*r'��D��-����� ����4���9}��H��
�O	g��B}�-d6m.��zi�6}�&PB�(q��/h|�$����Ν'��Y�H7��M��{�� �>P�
�@rq�	�MHPJ��ӓ)�S��L��sZ���s3�$��_[TnGƝN7s�F�}���Rc�n�P�>��Z��2�3>H/�OR�Nb '����g^TO핐��Ԇ�T��<X8��7�Y��t��Gs�Z�|���������ڮ�TC�6���a��c��E�%G��a*9\�N���؀��v����f�e%P�g$�-y���4��>�*,�T��}����@��4�9!�	���Ⱥ4��&��G`�!GVܢ2�B����)�$���2�ň(��h�U�I{��m�@��G�N�TJa���;^hBo�@��MN�������x��7A���x]�p����8��BR�.� ���0���C�P�S��{�����h�8[4��I޶G����jv��`
?$ҵX_�I����o�Wi��ϏWf��k̒G.�[���!6޶Fk>wFm��)6��rk���Di<�I���k�Gr��^͍�`>/j�3��a�W�����+o	�M��������$���4���(�S�����̹k�MH��Ż�&ٸ,�2��`�!����t�5A3s 2�i|��Qn�,B(�xo�O\pL��E���� ߿"Bl�^ �Ym�)�׵���!��uf0�'��-{��"��,x��0gk΁G��%.ړ��<����,��~1�48�˾޼_�l �M�IVV@@�����b�Q2ܩD�5�A~����%��ne��h���5&�A ~_��lf<���%�<y^>e' �.��q�R?	*<���#�Y����#���/Z�ab7��n�Lf����&@c�!�hW�"�{6���Km��������YݸU�v�Z��l�/��㓿S �h~�����ӑ�W�D1=	�D��͕W�1����`"���Qj��}a!Z�	`~ �G?�ψ���(��RB��j�Y]T�]�Q������r�q���@��RQ��1���f��4�T�-�Ӏ-4^�v�|o����]��;��ĢN�A�Zqܓ9��Mx��Y	/.��@�1�����~�d��Y�\{6�ƃ�ª���l��~��@\�����X�
�_���ۆ�� ����{G�3�p6u�"q��Sʵ_��J�
��\�~+x|6Pŵ����)y��bZ�x�b��r1���`�f�m�~-S(� w���&�b��a�T��{p�G$C�(�����s'qe������|���U)%(��������iXR�I��=��u�̞��ɔŐo���OdҖ>�]ӄ�b�+A0M��|-�_Y$��P�|W��4�B�!I�EQ�Gg�ك����e^gH�m}���u�R�Y�s�����鴷� � �l4�:˵IIJ�(�}*���'k�6�Fd��A��\�gn�Y|����د��gp���L��uCWx��
��e ��dF(Sq�*.��촡��p�أn
��m��=���؉��+R@�Q4�� ��?�h���5��������1ۜ7��Hꂦ"鼠� �3u�5�05�t����@AZ�i�p�)��H��ҮG�����&�Q�ӛ��4�J9u��Y�#�8�]-~�tr7]ȋĆ��cG�vK�vo��R�@�d�yz��#��\5��<
ʪ][͐\J"�~��\
�=9�zd��30>K����ڸ�e"�Ʉc	4v�l���4���U�"b��4X�u�`Y�s��4�����j���ӌܱ�¨����*�nuP�
J�ũ�^h�{7.����Y�k��J�4wr�7��&(q�9Ro�bѬdF�-�;����t��6H�������ZGɻD�����ZI��1ҍQ�f��E��aw��܍��$Z"��H}�Q�3Tٔ�;JR����,va,�<����-���I �k<��#ۈ) )�}�u"���ʷ��&�(E�'U�>EP#��,�2���x#$��?4�Ο_n��¯���y*c�p%ŕ�尪-�]�e۷�f<�����A�����f��6�fM�����HO4�?�v�hJ�6d*��?Y��Ũ&G�q8�M=�����{�Ѕ2-���;��FMV�x7��{�������wkk�^��#4��hk�"dw̳҈p���1F���ق�������J���>������18w]QѰ�
�Z���C8r��IaK�����,}����羙8�/��z}�;��5��@�ⵊ���N��ל�ٗ��IB�Q�e"���pm��jFI]�i���m�������OW}$�I�1�VN��#��Qz��]��."]�k3ַ[��F�x'9�X%����GFD�a��SSf����|���9��vv�y��'|����0~L�H�Q�T
:Q|G{t88�!�@F��Y-�)�mdn�i��1�ߒO�p��Zɕ�e|���6�P�N��hz��:�˃��w�ll<`"� ��
�|XpTJpm�0}���7�J.ij;����O '�ys���~q�Y]����+�*���a�4��#W�j� �b��G?�ceAmm��m�����O�
Yǥ'�l�H~������C�Ь'�5�^̤�]bg!ל!l�`���|���b�M�7MB�$��TQ@��v���N9f��L�[�����] ���ZFa@�B��F^�XUօ�Oz�m���p]/��89���m���w��0�F��@�!���E��gH���x��R�=��
	'�q�e�d�J�I� %����)�ӕ0|�R+t�4� ܨ/��`���[���a���l�*h;q�g~RE�ﭩ)+1�$�=���[�S����W��/��j&Ə�[��v+�x�HYl�~���;gǛ�Q���P�0�c�Ԛ/�P��9p���`b��eE��"��/<�����F��8j�������I�v"�2Ig���.+
Gq�k��MG�D�J����n�h�iP��& ��2���L�0��ʹ�3WCz�
�t���C�����ý3�w)�c��_��he��f�����Nis�Q ����.��9����P����3�s��\Ue���b�H=e=_�UrdA}��I~"]��4��^z?��C9�"J�f
iv�aط�a�o���7MP��&����Y����S�"�C\AS�/�|D�_���N@
����0\'PA�ʨl">�=X�;z��2j�p	� �)݀9����֝��*���s����8vS2�Y�mY�#;�XhE͏�H���e��mUV��_���2>�e���i4W� /:���5��<ڌHj����j}|ݷF�FkAg��Ӧ��#�rI���;}0<ܙ��jA�Y���arg ��M
H��A��m��"�c,���c��5�<]E��3�+�@��B	��B��N��H�gn8į
}`kU��]:�h��px��#]�.k"�� G�Qk\���~&��v�za�js�4�<n��mZh�"�J:���V��Y�](��`Z\�W�?p�L3��ҋv��5�~^�o������*`0���|[��4i�����џق�W,�3F��~^Y^:��*m{D6Q��-�eQ����G��ak���g�KmS���6#�-��Û�|�ǂ�,�����M�����$?
q߳���enF��j�9��g�3��B>$�In�<#��c�P��7\wy��SF�
��ͯ�fDĘ�CA q�S���+��ig���~�	dj-s�SK��F >�pe��3�k�A'�3\��������n�}S�=9�W��
�)�+����T�sb?"O�/5���n�����
u�6��dKm��|��;3%|(��j"��!�J+��s��%���7Ƭo������Vj��X�.�!U2�#�7��򼄭=t��'�=��Kpo^_AJ3��йi����,{��n�w�f�dލ�h��޳��DѨur���w(+9W��k�?�hj�6D���_��P�!��v�7H�����8�4e���v�\_?%��2�T��-M�����567M���3�J�$J�v���0E��˱�w�bt� ��R��g���!�>��t;��$m�U�JU�n)a�=f��n*�s���V�=��,�J�J`�����j����Lm��_�s�*�&;18��|/2�>~)�|��Q;k}��2u7����e�����`�F��ĸ� ��z�1H�lIJ�����e�g*�"~��mc �j��JS}�go;;-;����Ӗ���ڄ���v@�`�˔�¢��:��++�
-~�ͅ�V����m�[a���Y~��6u�b:�܀�J��K$<V��,��T';��󗵓^x�H�/���5c�A��"�EL�T`��ƴ�y�
�p'�l�s�=/���:��FUt�����Pq�������g����w��J"o&@���Xi~=��S.����m�������<�O馃��������}�����6dw�7+��bj#�?t��u���x]Gc����`��Y9_��'}��H�B#eR�,���`V�Q_�B�I�A�/be�w�C�	���a��.�a����z�������3KM�B�?�B�Ѥ��^�
��)�i�W��	���7���L�^p{(�
u�8R'�9�r1���g�g>	7h�����|.�T�(H��"[A��t�`u.��4+��7~���=��9(�x�[�!^�DaBF�ݦRP��!/H~�#Ӆ�1���'���9#�Dq� 
Dm�%�vw�8mɜ�{��G*�)��q�p���-\�+����`�L6wfc��@�D����Q{�$�v���^�NT���nd�SL9MO�ԝ�æ�u�	DOe�L�)x�9��/!"S|��~��D0�p���T�2
98 Q���w��_T�:�E3�"�1Ҧ� B�B
E0�^��n�)j˷���Kh�_�?�y\�{�)��z�!?�_`t��?d��!o�-'�.��$Z�K��Ҏ�O�MaTw4��ުꆕc���훩ǸnO�f#�y��ڦJ	�d�So��R�S�q��!_��Ǟ�Ox��3�fmQT���_s������`< ޳�q{AI�������4�C����s�]:R�����^Q�`DL�K�B&��T�kS}杔`������!��F.�8t��_�L�_�MQpͭv����՘nRRxi�BTUIkw�D&	��[6�}J�/R��ޟ��oa|Er<M�v�����O����ջQ�4�G�='�WP0P�Ĕ�	u��/hp�R������?VN�ˆ�<LjA����+���.)-�*�w�, ��M@9X�CH+*�������>S�[Ȯ��g\[�/�x�?�ۜ,�1��f]���PNU;e:�Oͣ�� ��X���L���ϵl��"�媽���J�A�䑫��;�p�]���,]�A��ӝ)
���Lh�|���%+�����qahU�x3բ_�j��rL�!4_ОEi'ԸF8ӝQzx�CU/�'��S2�j�~yt2>r!Qo�7����OB(ޛ(���T�]P�A�)ד-p����+�V&_c1�f�ԵB��Gn�c��O#�k�@`�}<�'Wզj�Ugc
 ;{q�;�����2'��%͢tf�K-�\����C6�����Fo�QdF�[��L�/�L����E.[4s~M�7�7��g���V�V*�u��� ��Cqݐv_��x!���e%��P~u�|�DAo1��{V�8�i��m�}ٜK��C³Ҋ�hA�y�߂ϒ����E,��:1$m͘�����ɇ02�U�+�F�
�?Z��Q�������U!|,kuq�f��3�{�t����[�3$���t��Hv�����ۄ � �f^i�?a�)c��l��r����_� �P�������jt��ƅ���w�z�K|�����	�V���,s{ACዾǚ7	��8��o�_�]���g��6"1ׄ�2i�L��AH�<2��Hy�A��\H\�g�Q0Kϖ<�@����ED�ual\ԟGz(�R$]��X�>��v�CW���
l��$��Q���~6x*ˎUN��T�GUp?3T�n���}*p�l�-tmq��ݣ��?Z�[��^4��.�o��4�^�#o*8¬�����:1��wۿ����䦎��Q��Q�*��թ�\�K���.?M#�}���a���+��A����B���#�U���E��Y˄�O�`�.�4���L�\�o�x{d�f��n	Y�z�^
��{�#�}��cB���?� �Cwk���\�o��[F�&9�U���_�,�7{�9�Ϩ���=O�/��,��K`�#�<��w�r�=�a��p͵� e	����TvD���	�+ɽd�*�,�!��)5����������v�`�^+��QRDvIm����l�z[��O��.:��'-������w��n@�l�g�R��l�T���|��x���dF�=�F!��������'G�Ai)�Q�~ U	�y`�x^���|5�[_�Ճ�$r� ����H���4	�?Pb�0����IF��'�j{D)UYŴ�v<fD<l����c��hx�ȧ����Ķ�]`RU���#�B-�q���h�o��*q9F�a�yW<��OH�\��9�. ��g]��Gv*H�|M�z.jM%~QUqm�	w�R[��k����vH;�[�����^��3Y��u�wa�s�%��: %\b>�v���9=�l;�z_@�i�
L:±3�䗐�-��m$y�Ơ��\���/D�}S_+���d��b*��"�#��7�PiwK13��C�a�ϤB����aV����ei>��p�i'�Ў�L.@�k��:�������h_7��T�S��u���uYd�)�LX��_��T����j>�Rʚӫ3�kH�)�-].�H�X[������}�r����/��2b��::�"�7��A�x�0ͺ���b�l疯#�w"�I5������l�o. ݐ��mA��w@i� IA,٧J���Dk�ȃP�Iq�� ��2Gͺ	�Tn��)б���j�U�
�\04��O��)�Y9O��6�y���d&J�m�Ý9�rW�Rj%���^"�6��W��js��Ĉ��.��υ�d���I��n��BK�+2s8��{ޟ���p�Z�2AKߖBYK�U��*\IK���}�Ę\����i����O��[K�+�B<�{h��6	Z�Yָ;����}�=A{y�\|(�����������E}��+V
]�������Ջ��ϼ���O˔��
>悝�ꁿ�@7��B��\�d�7^d�K��h�M�>�	H&�\�,*@ΊF	���O��X��mQ �}d$���Jߋ*+�0Y�������LQ�1����T$%E�D�X��}���ۧ�ꫣ��8��43�|�uqx�/�X�z�D~F��Q�I�@.zT��b�{l	�^Io5�B��#U?���ۉ���]���,.>v��kR�cm�L�����Ku�k�����j�	J�X�ގ`y@q���_}A�sC���}�}t6�H7K,v���7���'�:���W�n��%��$����n�R��c����O�L��H���&E�4S;r�x�����;�`O�x��xw㪷9?�B�J��&wA�^��;,Ŭ�IC���N����g��Kߥ馏U�W@
����Z��ƒ[�\�ᔕ6@2�a}Qei�#��N�����Y�����"� Y�%�J�V8��R���jW��+4>��+m��IR���J�y|����{�?3���Jz 㭋 ��&��g�;�Fn��PKZ�xL:@�X	5���kF^#��>f�g: ��u�J`Po>Q�$�[�p�P�E��a�5�(����dH�3��FR�/X��z�b)�Z~�^�[�`t<��>tu|�W3]���`��V�fo�Lx��8܁q?2OZ�� �Ӌ�]i��nb�w��sw���QZj�&��y���R��QQɅ��qNI�"�W�	X|��_ܯ\Ug�IV��n;ūb�E���nTژiX4T�0YZE��~ϳ���"��]��� �9�L���Y��� �Ù�m2f��@
�����H��x`�xQ�]לz����f���Y�6��ѣY'�Ũ[V���o-5K����r+��1Y�����x�~B�؃�uO����c39�v<|FAlI�Pa�KaS�dE*p�i�QZ�/�	�"s��N��ؿ�$��L�}��j8�?�:���hl#;��l/����a��)HaVU%+w!�Л�X�±���ׄ�����.�|a��7��m:�FT�!%Ϡ����G04G4]F��������}v�S����S-ai������&�Ǡ�9��LiY'|��h�(0����E҅x��)�WL�����]D�UPTwi��jb�3#��{z�]P��?GT2��H~E�3�^��B��s��un����@���X��'#x��%��P����i���5g�1O��>�݀��,A�._��*��z�G�����ۄA���������xp//��_E���_$�Z��.�:H1�^q��k$�h��V^�[�@��@]j<��^g�a��
�ېs�P ��`$�<)9�([JC��'���)=?�% {n۵@�;%ǐJ��HG;�=ʨ{�I��$_�̻��d����ش���T4�~��u��Ѝ`��B}�p�'`�����D��CgCM�!�ԡ���uHC�;f���ؘ'z�
��A�I��ڻ�5*D�ێ�� Vn+�%�*=re��OW�*2�\Cf,�g��>�`}����iF�M=�r9GΡ�9T��6��b_ӕ��'��ƽ2�W^G ��T��L��Š�Qѕ�[írO�B�7S�9'�C���R����rw�Aξ0���"R��όg�Ȝ%�XW�t�O���z$����h;�k[���iHe��8/*���S�%����'��*ZUf2�8$��վ�E��(闡|R�%�Aݳ�#�}�ٸ�D�q@��]��f=�B��]��}����g�+�YyR���|� �Y�	!��Y:~aU����v�qJ,q�N���o��SnqT̊��~��.�Ki%Ve �p0�r�#�p���L*�4��Y*��W���������d.�/�K�&�.����]UΎ�ӎ�$�?�y��w�R�Ӭ�|Ń%�1P������F���"��̶g����0g	��o���f�TeG�6��X�F1�-޳��� �h-ZZ�$����2��1���'�I�����f7t9�o��f5�W���}4#�F��FZ�f�<߶6� ӷY�*D��	5��͊�t򞿥;�� j|O�D�;
aM�_N�{e���M��T��h[�V	|l\W�����q��H�i�	���Ŋ�-����J�~xlCU�%#��A�yB��;�_���NW������]�����XĤ���]�^=ꢙ���ۙT�%���Y��*4��?n��c��?�l%�
�*�n���<i�]���'�\L«�\��M���G�`9�A׻O&�V�D��a�\??<��O@��mg?����r���枚��U��)�w"�Q}Z��ݯU7x�����6�OQk���(� �jL�qH�l�j
��2&�����{��M�S=�e���)2�I�CѱBҁ���M��e`�\r��M��m

�x|)k9�7�_��Ԋ���1�U}�_Z��?� ��bi)Ư�d�1o/Ѱvs��(bRE���_��)w�`L>2t��l�/>�s^U)�	�Z7f�&�Ш�G�1�x;���tX��A��̑NQ ��,wZ���䳁�?v�������9Ww>��/g�7����(=@}6�q��apD&I�N3�Zڌ(׍�x'�x�r9A|q^�:^
���'G�Q��c��U�jc�Z��K	��E[�똙��^�=@STN�$ەW5^��2#��*����>�V0`^Gv����&�H�Q�lT��TY���R�+([jC/z��$#�b%�YmO/���dGo��<���A"�����6�*���q��xR�K)%����`���e�Aw;9�zz��hC��Dt��k�CC��̭�36P������A��`���(�H��U��_n��}��ۘ�7[�4�ʥ|6���C��T��X��@��fElq�<��%����|Jص�Ęy��V+E�^<A�(��)�D^h��S^
�/������<dl��DB;�-M��+$��e�ɞ\䶨5�隙�Ta��}�v;|��Ap��/^�пx&��v�.�~xy*\�i����n�,�������+^}���J�!�2�z�؏]� L�4����ij��&k�AC�?�L ����a����9�h:�Y!ha�4����U�a���Ư��ç�&���%;���U��̻m�@�6�C�6+ܾ�5@�S������� �w�r(xG�i�� b�Q��(�s_��e�>��~"�������A�B�=O���0����v��6]��e�U�������0������ω5���KL�#8���l���8db�/w\p(��QL2�@o�{�)X��ʨ3���Ө�ͣ^�>��A��r�/�p-E\����D�" �Q�=�8���r8J6@�'@ #?ý�� 
9|�ϋ�̞��	�BN'�)N��0�B�����D���S׌�s�Dmj�Ʈ�ڇ5S�х;���=Ł�EŔݙN��go�I��(5�!�������+l1�<��Ai)>�5���}آ��l+f���N�Q�I�2O�9��L ����� �&Ceh�4�3v��.0�)��`�q��m$�$����n�@�t��wN+4�It������D�C4u�zO�N^��������<�K+��y�?�%Nx�"�  �=�3_�؂��pu8邖-:a$�H�
S>�G4U��7�� �BWS����(�z��̲Nt~B��������ǜ��`>��Q�+v��#�kg�Y�15M}µT}�2 llO# N�lA<dF;J/�X9��<ּ���p{�	��t��%E:��4���o ���%�_5��X1��`�� Cl���,Z�s�H��Vy�Y����;�R��6�u���P? /�1��C�@��I�JM���.��KfEtq\�r�`�3�I�Ğ}}b�2�^}�>L��i����詺͟w�o��l��V���r��sP�H��;A��@���|�ۖ|h��rK�TWh�М6{���.V4�A�`ٴ�s0��j#㵘ƑB`�!E�����kH�`w��XzA~�&�3ɃD��tN�]~D.�zIx	��
�����F$}� ��8�nkB^P�'
�,U�}����TqA�۵HAq�K�t�/Q#,�����)fAl��U�ś:pG�Kt��,�>H�g��N�r<m�c�M�g��^��/�"�#��[x�]c+)�ɶ�;�~����T�c7U�W|z�"�rˬm���B��>���"m >���iM������Nj����P'���\}�!���7ff��s���?K�6�����P�1|UHPmD�H�q�f�F$-���s�����z��KdqŰJ^c��j�� i	�f�/�Z�7��=�J*Ă�lҚ�$+��k�͈���r(����ėACQkܚ�=����j��P�tR��MF	y����u��Ԓ^;���V��q�v�[J҅�	�
��MP�U-�;�Q��?�gt�������RԷ)�CF�L���¿�#p��F�o0��[C�$��$�A�ElǀZ��u.ӹo�b�������S.X�v�G���nC�lw�l�b+�ai���i��h����ҵ$=$$)G�z@�|H�;m30�'�:	'�}��.������ȵj����2�� �wz���{ψ�M�Ba�ĭܳ^�,�%Y�n�Q�!��<��䫾8�B�kc�v1�U��t�g5����I&R��,V�_��1���}��}���r���:��NM��"��%�-~�ꚋ�!����	�,�Dү ��Q��2#����t������@�In���]aL�0�'��]W㐃�׈����6��O��삺��C�+~s�[���h�����Rvђ�i�Osn�l/�N;F��%$����N�T3$�dӾ!����W��
�L𰟑�1�c��aa=v�-�DJ�F��9��&��.���E�v,����L�g�J�C3��Ō-��J����\�����duEl3�h����F� �TWC: 	.��V�U1�6�һ\���Ш�9'�!�wrhc�zHL��
l���d	�[�m�?�����$����������q筂$�� Ng
��>,5�L�X��_�JOjw?f,a>j>������M�g����a�K��_f�)���w��5�<�]BzWfJ��=I���p4���X����PH҉�����|�E�uŷȆ4=��bN����#���ʍyc6+!�j�X�~r��qXp��RU_�x��t����ƅ�Hѕ
�V�ݸi�������b[{�5oY�攲�0��ӟ?��zʶJ뛟cUҀ��&Հsh��AJ2ҊR���C[9�v��8'N�8Z�v��+a�|#)��ޅ�R�R�RxN���w�Tg��������x}M(�MX,�E���'J2��m�|���z�#���c���������o
|+�*���'��F����4IY�}AU���A�ҋ��m6��z����N���m�C����ܟ��o��t��+���8-~����;�Wd���:{�t���Ԫ
@kPE��`�y�"o��P�1i����R|�ɲC_G(��>G�[]��ׄN?���t]�BL|tۙ��a7��|߉�쒅vE�(kAMäb�΅�-alىZn��wg����^�`���1P�t�%��.�u���?�L:��w���o��xYV�r䪲(q#z�X���B!z,8���ِ��.Ή��U:����� 2�r����ph*{V3+�SZ���6z���[�W�k��il|~�x��I(��g���mW����3���bj�F,Ì�Wð��w�Gy���g�[���I�(Aܚ#���T�8n�
�a��m ФU�F�d0fl���	ʑ��P��}��:�aU`���`F� �/4�v"j }w������M�[�J�۫��>o�CRK��P��u�(ĵZ��Ő,���7al��R;��j���3Rj�������54���p���-(�KM ;4h���a,�9�Ym��.4�ZrMI�E "����B���i��K��W#���k��I�!@��b��邭�qH9>�P��dݹJ�:>�ᩙL��_�sY��w�ؖѬ-;�����+�N�@Yp$�ұ���Yo3�
Ms�p���/V v�Ʋ��f���҅�W��ǰ�hͤ�b���og�+�K�'�l[�C���HW�-��0h]��
ͧ��tHkw�X�М(��"ō�tW�I�zx�G�V!���%��2��Jg����8SJ�f���!ﰻ�:=uF�o��a��y�	��@����*��Pp���&+����l�18iJ�~�:��N��WRƁz��z=!����|~9�sg܆v�B�Ɖs�!��*h�T�����ȃj����h�<�*���kr��O|[�٫�M�$)Vg](d�BǮV�$�D���5�ELG�D�>��n��R}�l>S������!TY�/���y�.�% 6[Lq��S���2E��XW��3�����kê�r�ٷf����)j"�ѿ��w5�2�[g�&n#�p�{������@TD���}�n��t�PBX�_�j�i*�3=�*qj�bP��p��S���rʵ��v��]���sN-��Z�E���N�/8�V��>�$s�y�*�[+���o��EXߋ�P(���NvS�va/�8�X�F���T����5�ۤL�xIgl��(�E�0 h�uFa�J�o㛵���5�^�SX� ]D_	��*�-���I���2�1v=;̚�w�k<�N\��I����N�d�' �_ea�vG�&l��¯��t��XUs[W̘V��=��l��0E��sؙEf�%�K
T��^Ue~^;ND�9�iHn�С|b��:�%�Ȣ+U�jcՙ��1e��h�F.�����Vp�h��[#Q��ȶ�L�0)d���z
%�Qh������y��v����<��F�J�D�["��@��03�B�qYz�\(�r��w���񥋷U��^�E2�9\�}���!���6�&^��=��w|��<�H��E�O����m��@��艣m�Tq�o�[�5�TO��W:g�s܅|^�{E��p��NqgՉ�m;e�!���rs~0�� <>���I�FFuLE�3a�<���p��5u�/h�����,����7�M� �r�F�ŝ6�7�>��Y��z|�x�,�?/*��o
��K�oI���L�Wg���fG���dY�%�*�Yg�R���rM\����P\�H���V*u���=�zAH��i��܆�������6���2ND�ּP��Y|�A辔!�&_>��֔w-~�N�٢�^Ĵ�%����;�n�yUy[�L/�[��j{) rg�d�u�@�^sVM-}2�����v�M[���l"V��T8�v��5��n��^f�b�՘G��MA
�_�^#y�����*v�ҍ,�X�Ɋ(������)$���H*U_CH������L���˒g���F7i�� q7����&��Gb]!�2'ZG��!����Vl��QSA�3)��]�ޯt�/��G&LWL�29�zwE.9]�q���ꅱߕ5�LH5*"ݽ�v�s�|2f�)�4��i�JoH�z��?~]�U[�����xu��L��V�
�9�w {�Z����x��ƲF��|=qq��\Uqc�		�]�(K�?��XLf�d�9�=l��W9��/�2�o�YX�/z�.��T5�u���n`rԎCZZ��z�Q�{�߳���E��>6J�r��F��ƽ�J�b�m��삘�f^]2�ɂ|C��!`�i}hm����.M5FG��Y��U$�cEk��ѲX<�rT7gm`���#1����[��@�ٜ,�CT���jLm:��7���]�b;A��U'͠G-���n��\u����eƖ��
�(C٩x�$�PbE{���c���Ќ
���vY�8z�K'7'�F�c��j�V�1�.C�>�XN^c˸��%�X���S�1�0N�cl��̃\s���S��O1�?{��9J��'�E���ol�ץb�R����vt֝NT$�ԋe�R�E���E1;��1H�p.W�n�^8N�aq7p˺�������w5S��Su�
~��
�����p����ɴ�����L���?g~��o�ȏ< �4��OT�́��*E�vf3MtC
<W�<y(ś�`�+�DJ��9S\�;8��z�ZL2���<�&��{���5��ˇ΍��̙P�7|�[��YN%��os}[�	���"�DAjX����lbJ�i���\�	6�	��W���T�2m��G�9<Q�8��E
�(��O�D�̯	�Q��� ��VLd�L+��� ��is�t	��������,yƂ��	�{��Lԍ}�+��ӗ����M�
?�)+�anl�8$��ցѻ����Z���M�1�$R�w�7O�fw�k�~w��c������3q�f�]`+��K���	�������f�%{(�1%O�a\5P}[�\~G�9R��Y�0��>K� ��83k�wq��v��J�) V\�1�x�rT�V5��vn�"-�����$���]1�.�$���:7*w�oJ�J?b����agQr_(L�3U�3̇�e����c�n�_4�����5�@�4������m�7;W�n�*ر�+�����jI�:�@�� #q����>ue��NC�d#Ə�B�=�]����w��4�v�f���7�Y��ʳ�K��%B��}KR<���ߑ��뷘�C ��1P�"�0���;릴(-Ai�L�q~|52�}ZD���������qWЪ��q�"�uA*�f9>Х;�V�U�a�r�ox�\?�o^� ;]����=]��A�x���AAeX܄�1B���I��$��PF��ɚE�X��|d��@'S;�X� ���M	~��z���S�)?����j��r��_8Z[ꍿ����O��J�6� ^���|��:��`lf���{�P�?%f���ڳr���ɴ@�E���pM�k]���0�8���E���[=��[�a���zo��J�o�Z�m��L)
�#��c*�?�\5n�J�� Oț�S�	^�����!�A��X��k���KfM÷�n�������YU�� -b8"�hw�-�M>����~��Pi�>����n��{l���k�@n4L�-�ʪLG~(mj	�e���M�9���;�7T��v�F��RaU��N�@�Qr�s{E��rWH˞�N�҅�*j�5j��Y��P��}32�}���7eJ�b���9`�䶥�D����]���"SAS(M��&��'����_��kZ��q�|k��n���H$Л!yg	̛�2�6�`$d���Z��j
H���.��Kj���E�"��iH���I�0�1�j�bV�5��8Ka�o��N��^P�D4��E]b��N�FR�j��v�\�Z��ӗWL���2Ѿ�n'�6!������I4�{a��͍��*��椿[�0�)�H��\����ɾv�@�T������pR�P[�<T���,��]�&@2 �|]fs��-��%n9N#���V Ml�����F�p�/'�M���	F���3� 7���̆/2�`�5��cF�T���#����Ԑ�����]pM�8��:�\�1(b]A��""�Qd�[[^6ɱ1�ym�\�ō��-�-�(D���5|`!Z�oO�q�hP�l�/o��%&k��-0hS�ൠ��>�� ����1;χko��O:x���퀲�6v�z蚳��.�U3���p��~6�����h�v�M@�}��'�w�-���߷�i*�vET��Յ	 ���D�϶|��-�����P����K۱w�[�|~ORZ΃
�[��Y�Q<�=?��ՑP��u�o�x�*�P2�O�� ���di���oԋp4S�,5�p.9��t�~�\)�F؛6���C�|,�]���4�!�AV�L	?�Gis�ID�"�.+U�iF��pZ�%\�t(�fϗ�)�)i����y恝�}���o7�aC*\bd��]��T �׻9}�-U��~}����#�?�~t�O'�b$�����j�,���̜����K��pH��E�*.�����j��{[@�@��"#�vhمP\�s(��3�6�����2w��5)��I�nu]�o;��~�z�7]ʆ�/�ص�QB^��T*�K�hW'��tt�J)��t��j�o[����f!J\���p����x�#�#�c�:{9�l�xc�N	9����W�1�q��%l�Gp}��e�I�)����r�B1g_���
֑�ʶk%C6����]�,�����6Y�q�I�X̥7��Po�(��w����s\�'��|F����l�V�?q �A�v�k+A+�Дz��4Y6dX��q0k�&�S7���f m�{b
�m}�ht�����#��b��8~.m���EP&Z-\�Ż�����9�� �1��ȍ���|�$9y0��[,�����&%�͑$+�¡�yX/�6 &��^���Ju*k����w=���]�9T]�t�X����E�+��bR/��`c���`)n�i�J�:߼&q�����NS>n��"��QǢ@K����'����s�;���E�g�Pr��������e���X�( e��W#���=�HF�h9�_��0��)�)���^(!�^�F*�V�s~X|@ѩ@��_��	��3.n�Ӈ^}�
�A� qE~�v/�� L^*��Z�x&4�:1l/k���'�`畊D����ٞ;�,�S�!��m��%��8�������|�Z�
+K�� `Ͻ����銸Pĉ��qu��&I(�B�o�V��j������RTg��a
�V�p�rZ;A���,�%�!��������qq�!`����1�N��1�gf�gt/t��;�P�r�
B�C�"(J�G�u{h��8R�bay��{O��A��`�a���bA��b8K�Wf7HId�
"��	�����v�s@�R���<Yi`��L^{��]O+,ZR����X	��Ƌ��Oсk�缁H41�t�������R�[���R��)�$sָN�u+�
�����R���Uf%L��|��fFk!���T`e�0f<D��O˼�Y��6s�GG�z̫W&
+�H�<��6C���JImp�8���`s�˗�r���{�қ>>P�R��T��4;�ɍ:�,���e��Tb�x�18u���������j����b��;=�K���򦋄+��`&�������"̍A|����R�t��'�'e��̩*a'�ŀ�>����Z�C���-��u!�нraӮ�����x�40��|R�_j��	 8x~P<�����S�T{�����l'ق��%�2�s��	��d��!���6c���yUuĮ��t��x�0ץ6��j��k���^�;�-P�+���;{�[o��%�l��\'��7z]��'�~��!}�h�>(ػh�K��_�f�K��{�%O(�,'��}e7���g���&���ik�x����N=s����oSS�˄r�qGPʻ��K+��T�>)$��&vO�|��)����d�	��hԀ F�)ڌ�L$��Qbʆ�2��ZOS�2z�Hu���٣ϛ՝��A���LF���#�L��:��[���R���-۶�.�P�QL��x��FW(�I��y)a�sY�'�ȳ$��Rѻ�dv�!@,�� 9{�{-�~�]��ZiɑG�DnJ�o�Q���GR�Quyvb����A�k���ѳ�c�Ǿgj�	J(8�G�\�څ�C�T~�;������*�?	"����t2����5	b$�Am���'�@��Ї%�/h�辨林���r��E`��5�N��Lh�#�Y�����x�_P�3���%PQ����g���T�S�%S�B?�]��E����U���Ԃ'��͂�v��Bn��B���B������ko~9����pZօ�q3��<�ָ�[n����y��f�B2����eX`�I����sJW�'=��m�Q�������ДV��tdJ�N����al�E� G��%B�8��-Z��X ���M�3sS��-E�
J��sPRG��p�Y�&]�C�����D�ţ�
l��@�&	wW閙1�����f=��UP	b�k<������J�!kx��˹b�ϸT�)�%���y��NU�.����[߾O�*�FRÑ��@w���j�Ճ%X�e�o�;��`M}ۂ��dgݬ�<�G�!�4������}Ui�ŵ�ul���;xj�"՝H��ެ�:|���]�i�9��2Ъ��oI��m=�ڔN�^=i�^rayJ��!�����vQ���U���K�����)��RA������~�s��;Ǌ����h[��P�4^�Xt:���F�r��̵߈���O�_��b�ҝ��o�w�#������Y<l�%�!�|T;�Q�=/�U �[5i��)��vg�����U�`��]W��J퇟5YГ��S-&۵�Q)\���#-0:!�F<�G��0��G��xT|w�Q@��0ey�dQFBu����<_i]l�܊E�x6�G:���7w�ѱf��,7�j���C�WUB����������(Ӛ^u�~G?6��ys3��[���-��	��Ҏa���9�zPE�;�@6��)?�ѐ	�y�ܝeH�(W��IM �G��7�D�U�(!���y�Hp���{J��L?�u���*��E%fEgC������*ˀj�2�:�[����#���'�Z� �>�B�p�3�������w*+�N��Bм�-���DD�?�'!�qC��7iK��u��	����0�6AF��9*"X�ȃ5` 
�aD�H� �5`�PX�����9�x��pS��XK��q�a�G�y�a��^�6{��`fR���j�bt�/yAC���i�$b�j�]��:b0�6_ա�`.���x��Q�G��nsa���j�������8jy�he�����*�g�/�,x$ܳ�A2r���m����9bt3K)�^�����ڛX��ĥV�%�����9�^���tH� �,�V�� �@}��/�P����r��~ٔO0R�Ͽ�gw��{���)f���5��cd�5'ۇ�����f�:��"|��ye���[�S��\��2�W�FL� y2�p��E�;S����,�V𲵨qs��a�����z4z���j�A�t2�4�K�甆��Z? =��]R�G\����Q�������'+��3�������o�?�:�^�/�����҂����~�G�\����ٻ��Gj:�pV<|��q���I�7��z����#X��K�5.��O:^��K+��p�ցM9ϝT�x0�4�\G����9���rϒ.q��t�:�!%�"j������L�5+���V�`�_I�w������Ŧ� L�TV)w4a�$��=�T�M�|�%M/,�!U���0D�
I�\�Qv��}H� ���K���=�-��?s��dN��H���`R���ؘ���� ~�@4c��'����hh��O��%~��آtȰ��e���'�z�KQ�w1:"���X�/�;���{���f)՚�9M�e�&��݅¼u1�*���G�����N�>z��ؑ���#��FtΌ9G f�G��O�F���1��'�ME�5S��A���/��2�$���w����	+c@�p3H�[Z�'%$ߦbZ�7�y�v��w���9�E���gi��_E���Z��p�w	���u��u����N�]ۀUB�E}S���*��D�`��jkm�p��?�m	����NZ���A���ʐ�i�\�ώ����ɝ��W�`;�����LN��2u¶�?q�x34�A�T����ش����}.a~_fYz �� X�:�>��$�����B��:��h�����!��k�.��7%��ۡN���nT��/P7Ӎ�Ȧ���8���c� �G���J��C��"��A!JN9���z��]�!�ٜ�����\���ǂ��}�Q�cI��+���{�_�|�96�6E9*���?�ƻct���T_��M��v�z�#9��f�2v���*�Ds�N
��)AD�}5��e&V|��{�cXq�1�L72���a�0�{ܢS��c38p���R�SF3����.�������ў����U��vb*��$�l�(�~��zlw�?}�6�EP�g��^[Z(�@C��&}�4�d@�?H�7I\+��%��ڪ�#��R�3B���E��V�@�|7�]����.��=����ëf��ܗ�_`	��mW��ƕ�N��${m�b�+�z9���d�+��k:��l�[�{h��;j�s؈g3m�
��J! d�<�Y�>�<��N������-q��uL'@�W+-Cu&��@�9iO�i��p�  ƞ�#F;���8���g���ǈ��Q�<�Rq��������|u�Fu!��p8~YE��jG���Jr�YYQa;e
�eK���Vy�v�5
gx�^Z���m]~.�X�0忽mx���P��Hs�w�X��Z�ߘ��JR�O9b0�#����-�7����ߙI]��Ybݴ�#�+�\��o���zo=���DJt��ŧ�w Z���0�F1�횡���&��9r�֓�����5�����ߚ�!�h���Lz���jx ��d�1�s{?8����-ё�xE��s���8��Q���3�����g~qJKn��鷲�7k2�wt�����%k)Թ�Y���CM�9?n�i�R�[�}4D l;��GLgQ�m^Zß-H�{�oݬD���IG$u�Z��e���N�M-�[�A�i�D�jYP���|g�_/��c�����	��*iQRO(i����V�iOZh6�F�v�Q�,�*�����$lyM�W��s-��=eK��T�<�0 jR�/\��`I5R�e�0D]���Zj�u���D6Y��^��l6���&�-U���:F�fm�,i�ч�(q�JSU֧�;��p���qѯi )1{&?����#ض�(�B���Gڷy�B��0Y�qsW���)��m/���j��)]TJ���P΁H:��c����\�h�%\nuA{W����V Gw>���`1��	u&�#��|���Э��`��]�ނ��-������k����' 7�,*{3^I���4|�m���{h�K�n`�FnW-����%TĨ��j�>����?�<��k��'�JS�џ5+9i-��.<E�6S�8$�P����`:���O�ڗ0�x�r�xu�>@��A�0}{U43�����|fg�Ɩ%s��"�G�c��u◐�N�5��Yt��L�TEM3=<��*.:/�f��@���_���w�7�=%H��a���o��G�SΊ*C�}Ҋm�-s%�٠)(|5�яnt�]��9�#���A�xp>�-񥨯�T"��2�`�*�@F �j����{e�d����>���^��N� ����������j���+ŃY��OF���3���ߩ���S���K������3߽�Vu�Y$&�D�f���!�`1��W�P[�<���Bt�h�v3�'z��?Y�~��' <��M�r���I��j?�o�%>֮fB_�i% -�T�|�\�A^=��p��X������4�h���P�<�Ř��l%�ranf�W�@������վ�2찼���=$�o�~�$ɜzF7�?�wK��!��:��)�3H�o	q:�����P�u �s�0�2��y�'q��Zk���c��wR����CH����}0
a���D��g�	|����L䩂��_�!3��>lmǣ�f��g�Jm�99�3#s��ph��Uw���D��6`���#��K�J]W�7Xs����$��|AF@�3+40���8��c��q�KP�c��K�I͞����ψ����j�X����q�:��6�h-�G��g�������n(��8 �Hr��W��jϹ��w����p39f5���PJG�JK7�3k��}"EF�5�Ә�,1�1�S,E��3<��{�{84K�Q �hj�@+?�k�:���jRժ�i&�~jGJa<q����L}`�V�yAF������'R�ht^�O�i,�N����WWX�H��z.���RM�jW *9��0��iw@k�(�C���D���|=�2��ܟ�S'����+V�zS�r7�*@�~�h�ˆ�}�C7[
QU��!U��Ei����t,�Cu���wii�>bA���VCN*XU��PǤ��
ADM�E�J�jV4����\�[�1E�4������Xʑ�E�9	(����tD��[�%�3�3�L�<�T`&2o��᭦��>��XQ@r�}�Gޑ43lu�l&ݰ`d={�|�y��I�6��%98ؾH�d���x,	]������ C���K���h�# �� �+q��X'>E
x(��+ֈ�tv?�.N��`#!�!��"���r�b���� ���5x�����C�n��`�S~���;-��^�����#���O����T2��a�\��x��R٥�]�Y��+ڍ�C�hkz;B�yo<]\5.��DGԋ�ݹ��eUx��r�(�p���д�OW���Ha`��t��.�c�OGsۉ8n��N����U��9xP
-�1���Q�y1��B^]~|{+-�X���g���v� q�[=8%%�!����0�T��s���!'���&��� bR]e����fs3w���l`z'ao(@�i8����d�.�l|��I��]�|����>Ke���5L6�|T���vT���LH���{Ӏ$�d�x��D�P�$c���M]t�>uq�Nn���dR���O�e ��j!��Ҿe@>K:��i��]�)ǡjZv�['�H�<���[�МԬ��2�<Cr��@�����Em���cZY�F���W �����096��⹞ƣR��PV2ih��5�(�`�����#��)�-,�Q�׳,�O��13<�c����*��	zE"�?m����|=��'��H����Ļw��϶��NX� ���8���� ^k�&m���态��q5_7�j�H����	��z_{0���Ul�J�+#P	ϻ=�nI#>�!���
���~c/�z������]4Jr��X�)�r�����9��N�"��i�E��+�6JBF!����1q�q��L�8Q^eN�ȝH���w.��M~��҃[��O�#���;��D��Q�st���w	�;6r_�h�d/��Ť����h�¬���h<YF�N'�v�I��Qad�k,�����.I����G,�P��o؇�Jv2;ro�	�:���S���Y�:A^�>�XG�\�����]�̅�^ �<��ۦ|������ty�C�e��)���ԍ�C�{�W��k��'�EP]=X�T2�3'9�ȹ
�!�4kټ5�5����%��� �����(����H���*�Q�&���י1����kC!��=5������A��s-__��4v��đ�� ss�Nܞ�z����+��o�hIfq�z�1N���g%!�o����+�)�uᝎ�Y���(��&���'��VBq{Ħp)�d�N�(w2շq��`L0��k��z�t+�J�1��(''Fd��e�֬MU���3�XC���� k��z�+�V�#���������f�w�����6+�_��6���Ǧ��<Л�X�b��#�&O���P���_%aN�ȵ0�ǎN�O	8�V���G߼���f��?e ��KJC���:�� N�.�jJ�0����,����N�3��:-�>��.{Zߖ�����քV�ȟIƺ;Žʠ�^���rq6F,��݈��zr%�Du��R�j���F#�f��e֨�1���f֌�D��Ȗ�bO3r8�|"�38�{�s��!V�&t#y$5J���`M��a`B���q>2ט#����8:g�2�ta�5� �Ӳq�h=�y~���a����͙9X����G��Zt��#M�6�"�ݮ��Ƀ� oU��Y�Vv�^>1�\�9��3fƃ��6/���l�/�4l�h|��x����w�=��<�÷5%^i
���"���(n�)e޼��#� ��{p<��"@ŊJ7������ek�5J�|9���/�C��c��Ed._�����lb�� �ַ׶ߥ^��<+������"�A��A����"�P!���*�wX�WZ�b���n�?��"ߊ�y�D�������Y�`Q\<��B͑+��?B\P�
����j����vD��S�i�m�59h�Z��YBo`G��$�pb��9r��jɍ�+�u.Zx=���Z&���Q������WӴ=�eW�N �üd���p!Z���~=��� ���'�O'^~��4_d�U�9���U`����w�SDI�}K4���צoF�w��U�ÌEc5.����to�>t��Z��-��U�[���KHź��]&��=$?7�l,������&�����<�hT��`��k��:��K��э9�b>$n�̙!���و<� #㩘'[ 78�Y�3�n&�o�uj謯
���u��-�G�슐D~*�j��K5�m��}���D�V��'�9TA,��Y��wL1��w�D�?˱�ԟ��N��g��:�	,��ͱl*�%�H^���
P�W ���/YM��acK�9��Z=��J�MB�� `�0��,E Ce�Yr��n����o����%�_�FfR5������}��v8Шn��[��|*�7�S��;3��
��תh�q��/ڟ����xai6z��[{�	C�~K9�C�5�k�j@En���Yʀ�&�fF�]F��a��N�*Nγ��kK�Mi%�`� .���!Q�����S"nh$�Ot6��.�hm��䨩��A�7�P�M3�#C��P�ϸ��}��Ō�U�&�R*�ĸmai��E���R�]�θ�nV�1�� �%6-M������Y��w��0+
O��G��
7��7��tC��WUt��ظF�B�z����{c��%�7?��X׬Z�pP�9W��}�Ѕ��i�a�#�[w��� l?�π�b��,�4��J�;�򙊢j��>�֖ew�+{A�2&��N��S��b �k��o.+��+;���̴��u�.���T(�C@!�|%rJ�k9儕x����Kv�GO�$^� �\�1NQ�mU�n_KT��Hq�*�w��c�cۆ�]�ي� m��^����lވ������տZ��Ǔ�D%��2�٭�G�� ��o�� G�f�
�P�E�&@m���B:,��.q홉���.6ن���<�{%��Ve�ۣ���`ƽ�'��q"2�*t0����n�T]� ���J�H9�H�
�~G�KOʙ�"���]�;T�l�Ź{����V��ّK8�%�w̼�~/�������ƿd���n���|ݰn��5P(_�wٻ���
���D�r �R:�����������<��qګ��w�zS4�r�o�_U�[�8���lW�<5��ը� ~�s"y�wb��t'�)��ب�bY?���c�|�I���"+T�����$� �&ߓ�|�׃NL� 6`8���}�� �B�W\��n�·�d��ؾ��a�����l�tn*�,��C8���Zf��鼲˺L�����.Dad����4R�L�:ʳu5@�R�
�C�n���3���^���d=Ff��xݱo�+PʥK�ڭ�i�FQ(��geQ����Mh��\���x�S�	�;���x"��+8<f�g���-��J��Yy�C������*�=/؜��[�u��ަ�*�B�j�:`Ǡ��;S��H��$�WbW���	��/�Z�^�6���DYS�cS�S��n(�;-f�T��3�>�A��9JX�5��yq��^��1�0��6�PSv�<�<S��y����6|�P��0tNy� ҭ���V+�`׆�%U��Q��j�B�)%Z�=-�(��� ��r\6�c���4l�<>)���r���W7����ϐ���ZZ�G/<sx|T��5�������س8��F�(��r��Ѐ������/Lq��8�Q�������f8�r����Q\��1��9jRoU+*���nrT���{k�;�Sb_�Ij���5U/)�!?�j���~j�&I�t�,��p�I�y^�`_���\7�²�=N��{��\��A��Q|G�?��;q:f�p))v�1��������b�P��<륈�	���YF�/��h^��*ODNf���c�)7
s�,�,JA��'<[XtEIu*J������ku���o�O�*�5Wɧ��}��z��j/i��7Src��!�"��i�����f��R�S��j�똲p<�Ċ��z�~?�����6}$���	^���U0/��-�ov��W���t��Cn�:=��ZBId�DE5��W[ι��!B����0'$p�U'(*[�U~�� ��+R��	�:<f��m|b��؍�g�J�Pl)��)���oJ�����KK^������;1�T0~��y��p{��, Hϫ�� J!b����c�S̵}F
��@/6���]D�mF�o�)$y�t�8B,�9���ĩ�ժ���z�r�;i�^g6����`�S�Mx��`��p��fwXa�����U�x����V��O���2�b�'7�[�p�.;�;2�/ȯZ�"ߥ=<���f�����N o�T��Ԍ�p��)�c���_G����`љ�4�b��G=���X=�	�:���U[i��Y�&����:�AxD�f��nO���C��8/u���V�Þ��U��]ꑍ�`
��������a��}����e1�jb���j{H��_`j�n��k�;%��&�^�g0	�lϔ�$^�6��\[h���h�,�-D��
�jzcui�pD���J_ ��=66>���q����"�o����f��� t˸ײ�D�ۭ����V���Bڷ��O�qNTN�
����cd'�	�|�IT�@s~!9
�U !qd!P�}rV�`���f ��i���W���wu���y�Z�u}��ҝ�K�S�嚆��j�ZZ�8����|�2 �?��A��5�=f!r�~@��jŕ�m?�X-��+Z��u�k�v����E��
6���o���Z%�А��ƺ�J���j�*��OQ/��iŠ��.����{q��3#]�m��\L��S�xk�׶hU�1V�=���j���\� �c�.�\�̦��GĈ ��CvS���G:iS��O9��ۮc0�h��
���km�Q���x~�ж�_��A'[�n<��HH0�3��~���b�}af���t��%���+y���~��ߌ�f�\X�~@_�.ȫ����*�ܵN�/���-;��b�٠�PkfW��K��\�n7֩[Ǝ��5-�`p􋋻w�2���ݱ�8���||��AUJ�6Yώ!��h?\�-���\y�6~�Sk%�0�̦�\�r�mJs5�I��l"	��vN��e���ξ�bqʧZ}�x�v�w��~2�qK�*f��:&tU^~Ys>�k=���C|�ANsVV�K��t\$�0eTO�o`�<M�{�*��y��ٶ�s&:�_���[աS���Zp]�n*
�x���K^
�iv��0�w�/�9�|�v37�A&�W��g=�]!۪�W�kE��<�����F�E�st������Z� �>�y�I��T�凁����5��pU�<	4���o�6�f�.� szt����v;��v�lZ巾K�]�2}DT�t���h�"u��M>�"g�����G��Pջ��A��!�)���X�0�D��� Ə�ՙE�M���jt�{����aΒ���y1M$���)���o�:�f�^���fO	��J:#�����=?�u� ��'zՀO�';�G�М*=�E�ԍ/1�~?>{ܸ}#B߬�=���fI�hH�R{x��j��;2���c�8ɔ^n��"�=;�����/�
Aq�I	d���~$�ƎA�E7����?�M
�FAѿ>&1�N��k�Q-�׈A0Sc��N�� 7 �5����0�+)��.�8ɡ��|!Zgۜ$�=��n��V9_�J[�������WI���=垩����<�8��J� �Xf^��l�����[$L�'#�=�\��%�O�z����.vK&͞J�h �l �gݜ%�"��]i\$-y]�Yl�Jz�A6[�b��V�&_û����,�"�WiZF(����p<4rxV��t���ز�s�/q� ���2�D:����|�a������ax���82����D7��n˥Zx��T�ϕF��}5���c0ф��c�&Ƚ����Z��/,�*/�p�(oD��D!��ãs���V��%��Ͼm}����uTyS�m6��F��⯸/���ʑ��
�sd7�fٓ�]qO�R4ʃU(-�J��Iډ������#��云�}�e}��ꦐ?-ND�K�V.e:�[s�h��vr]�0E2U-(;�|N�4C��hљ����U�zH�.���&��o�K"ܖ��
��
~>~G��[��8lԡc�^��wt�`�eBÊ�2~IVo����c�>�:�p@Q���"���(��;M�	�X��7']N)[�E�88)�/p�Gh���9w`�I�XP��E��4�!�w1\��ɏ*<ԐɏEHI��~����`t0��%��@�ɷ��-�i�C�
���N]h��w��������J,prpQ��u������V)�p�:S�D�����Ԙ��֛�<�gR���YOEEX���խ���
Rm�DĆ��q��@���ZU)h���e����d�f��m+ކi�?D��sꄦ�Oِ��{*>4��fX�T*5���ܑ��o�an��`poqvs�� }۱�@���,ގ��Wi���
H-�1����Q��J�$�	�/!��Ď�սu^b8�^ҁ�HޫۅH��%0:���x�X�[������?I����зWyw��Zo��S�[��J�럠4��ӏ������E��|)⽭-v)Ը%�7�I������OΥ[5X�J�N�Z����C�:�`Pig�d��1�l���X�m�����wׅ�����Ŋ60*[k�\�دT[|Wx�2]��V�l���X�u��c�eE}���`�"�: hR�W��j�>��|�lЪ���=�|�n��J�}׋���B��}�"O����T�Cy�+�N�š=�=��\�DNY��� �\~I�A䴋��Fg�6C�ܸ4��8�mn�<��s�t��o����{��z�M���]<��������I��a���]�5�b�t�v��Cg���R�Y�?��!���;Cʣ����:���]��C��
�+��Rn�HO=��4|*��+F�߷#h�D]�_�����w�縉g\�O�(���qqa�nV��=;��Ǵ5�^d/3���#t�wv_��I�����p�E�޿3�P�1S ��CkMF��"
ד��N�1A�՜ѿJ�����D�@W{l��,�+���3S��h�΃E3c�7�(�8;Yi�7#�`9k"����r�<��HSe�o�t7G�*���T�[�q�$�9�"Ry5��_��@�0��*N?Z���� ���U��t��`���S�v�n����h�H{�j��U1Ǣ)<��o���Q�,1���)��0�ױo�8Gy�,!-Җ��ʶ���j}�kZ�&�?�d�wa~s����%���ׇ!��/�,����1��Eg����7�yb�>�j"m����0	�*�L h��vk�����z�ջe�%�BUTN}�8��Z?q��+�5F�Xƽ�+�R�z��ָ����=��(��*x��|uZ(g�+7\�k��xk�Q��/�ug��S��H���䆫� }���4OX_���H w��J�)໅�������6}��#�u��$d���B�๜�o�����HT���P�"4�_Ɓ���`)���M���!.��e�
��g�ҩJ�ꪋ��D 9��uV�};X�R�w��@�������Gg�ӂ<��o�1�E �G'\֔e~���>YgL�������/~����U��0�lc�|�mw��9�b������/�|Ay�j.�jM��p�:��jٻ=TL�y���(��U�M����C|I�PN�������g��C��ڥ�/`���ыsE%��<��Zb��{p��]�k�Խ���D��8c��c���=�I��(��2�Oj|kX+R�l�0�e��v���Sy��k�_vtu��ojhe�h�ku���N�����$�g�@6#���(�d�Ip��H�ꯝdx=�ocGN��z�vR�Ǒg�����,�0�i���9yHDG7�˯����7n�w��}��ǅn�`� 
J���S9�8e���ѠA�R8J�0x��A�VR��3^�s�������a,��n1U���:N/�2o�$��Ж]2b���=����y=�1Iq�����.Ua�gDy� �F@�>l���|@s`Ad���8s]�A��S궃�a����̜5���M��v鈸�eo�<�\ctN+p`歺�=�Y`X��MvU	>�!���)F$.����-*�#����4����fw�e|\�~`;"�.}��	���n��B����;-e�pha�J�y�Y�wB��e�2��0ی�D�:�d;���h%"*�I��0��\�u��T���]\�n���J��M���1��F��q/#6���XO���Y�����ך0�燨�i�i�g����S_/jzf�+ ���}���(��u-	���`s� >ɵS���:=|�\����6H�JZ���f�x��hW���al��+DH��S$!��_/Mp0P{�K����SC��]��[���
�J�{��+-���o�#p�P��2�X��T"�(rg�0;ں�tum��� w6Y�
[��)�'2-ր��K����DY����/c�r}��F�lSI��oh�&��%��襎��U��-�#O*��8	����|�wlZQ/`��>��hy��~���}S�F���C�8���]S��c�����-��+	�r���Q�A�}��%IƵ��*-A�\\Q���À}�x����}��I3~�[� !�j�L�=��dj;��c��L��vs�Ҥz��c��%�8�c�j���X�<��\ߙ0�ϳ��Amۺ\-"'\�t(��g�(�n�D����ON{Y��ץ�;fj�\o�O�� X�/p*
O�T�����;��;�K�uN�應�N�"����׫��%����qls�ɜ���"�ʛ��g���<_�`QKXs���B/��0��=�?.loha�-�~˲fq߿����/��]AMM�ZA�pinF]�1���<Ⳝ�\"O����73���R��۾>�V��B����F6�^���zH�fkZQd�{�.�I��᫲f/��!N˒I�Ig�N/�j�O�ߘ�<2�5F���Ԉ�������*XA>R�����W�����}���Ã�m�J��AOճ��T�Į曙�	!�Fg�3p6�b���ȷT��y#��/¨Lx�<��g߆K�t�����6�������(!�B��DL&j- 0l9]Ę����p�!��� ��1���x��U�_{@���	#��ͺ���@��L�� �����`Z>���sc(u�9\>4�p*�"�����4��sj���c��>��O���6.�O`V%ȴK$�GG��:�z_>ZB��F�KZ�d�xP�+d��@���6O�i�ɼxƵ��7H�U�|v���`ԗ�q�`��2�Ր��U�@�W<>���y1��IL 5\���5sAN`�vvFi�>3�[���4��*Lv]�B�3�J9����~��j�ᤔ��-�cJXl���O��LM�B�(� �>^j<ꚲ�%�z�/݂�w���:1�������X䄽�9�on3��ن�	uD�_���7��rg�'�mόh�	+�"��]�O�_c+(xcqm�~����B3>0w��e�B��w��	$���K�={ٍ�^7�g��P��{�V��W^8���)w����÷
�^�(	\�0�wyK�<ڎ�4��AE���I�:Hs90h�+����Ūk6����B��82A"�q&=�t���OZp�6�ff���F`��&�;��:�۫� `,�	�?+X3
�>�=g���^��X��]���y������<ž-RD����h��a��̄�y�\��sth�hL.#�dW��:�֥�!�ߡ!2�P���(������ҕjJ:�F~��K҈��	\�8���ɑ.�W-���A��uQ�|�o��l�����F~�KN="̸����u�.}��p�������3���r��?��@�!��Wװv��oa�H��&Y��� �xpp��94 � Bc��v���0(�|���ֳQ0c����MA��!O��,#9^P�����y�f�$%��6#//�Q��3Oa��w��eYl���n�;Y��� IП������L��QHP�a��[O|$H=Lg��[2�ާ��5�W`��MP�k֬���>6�Q"t�/��w鹥���+"Jf����2]�?�:#h|}F����}aZo"��5������'1Z���P�L�y�c]�i\ ��H��l�)�5'�n~b���0�KC�$�����\"['�dl�1D	�ϡ|%����"�S��?̇�xv~���h3f�u���2������;6���z���.E���~`�L�.���70���D���+�|6��v`Z�)��*4��Zh6[/�<c���+{��N���]��

���.n霃�`�]4ۿ�6g���1C��\Z��Ø@��Ͱ��܌nP�����P�����JS�b��Ƕ����3.>M�޷��NP�P�2Ǎ���&S��_�F��K*��m�����`�&�:���ƒ�g�#X(!Օ�Z�l�+Ɉ-K�7=�G�_�3���Vh,��bpr�iҵ曘+{Aa���e���-���K��]ä���#	���C�/��:|��&ƿ�W�+�F��'�T��%Q�����-�ũۘ�^�5���la:e���Op, �?�j��M��P�FCs��1�)�HP�I���+�ax�!>�<~�~&���R�|nrXr����?Mp�FbFh��1��de����D|&��w>u� ހ�)��y,�w`wGx�t��iָ�_`$ZO(�J_ˬ�DZ�e�����
k�#pJ�8��.�(���	�͔7蟷ޢ��10#$��m�Lq�j�<o��r�2ԍnW[��T:Џb�u��S�a '�â�>'Ӹ�ׁb{9hȈ�	���ߣ?l����6�_HD�o�e�W9�"E
�����,lBl-&��ހ�k�9Ǆ1���4G��䑰���Q��=���qtR.���F�:������R�wCv֢���b�M��W]��f]�QN�}^m��*o|�?�  ��ɻ`4@P��UÊE�
��F�WH���Z'�����
��Y-@�cG �Gß`{xy��J���if,���v^��Z/M�@����Rx"c�L���;�d�U�i��:Yo%�e�5-�S�A����(8��B̿6Њ@�gH��f�bo�����K���wI�;ę^{{�!ڐF���C��U
i'[E�N
2*v�����J��v�]%m�� iR�������А��)[�߹�1h�N�H[9��&�C��+d���0�<�_��gb���,��6u�b�|L�ś�&4�Դ�GPQ`���������r�<l4��c���_��v�Od�eO`3"�����$8hA�$�|��K~��띰��m��K�x ������uN�S�Q�̮P�8�D0���E'ײ@�(��������K뎫�᫰i�r�>nn�����z��d��>{%!#�×�877���j��fC�f:%aA~�\E�w�(T6����(8��ئ9ʷъ���ԏy�R�\���n�8���ذ� ��?U87��ރWE]Rb��Z^u�:ɖ�:h�y]�� ����,.���[R��nJX�k{	�'�`��v�3�/����݊Vhkw�f�GpS5*@�C�c��.v#NB5rlE߆O�6kOj ?m�[".�;8����=���w�ؑLK/Ĝ�{��_����N���=�����Ko�٫1���xϷJx�U�".1���搠��[�8���u����.�	�)A8��J�z ����_�q���u��Ů�UOҏ�E�75��ƒ��?i6�5RRq,Ԧ-�<!�(\��]JNۨ�N�R�����z;�J���[-o���~�J���on�y2`TA2�wclp�Y���`���s�����_��>�l�G���b�4�~�,EE8�LnnԸ��r
����К�g�ɢ Q�$vg��C���󷀗Gr�D��Fɥ�v��c��%
9@�6��-.:��Tn���������݆��T��<|�P�".��y�09��> ^����m�4s�d�<S�k�����므��M�C)��3m|h�M��U��/4!���96R)��,� ����}�]E��n"ݷ�b2�2���k=ek���lrl>���LI9���:���J0�}9SH�$�\�V<5Q=�����q��?��@�������q'&�Tǥ�YVa���������tm�]�@yK�|��^F���=~�];E��z���H�6�����p�p7��I��;��%N�F�_� �*�Hߞ�`S{ί���-�7�L�8v���+Jh���^47���)㷘Sљ�a&��Nw�H��>�~X���K��mRш�����?q՚x����:��Cxރ�g���u���"�7�H��/�S��$��[F�>�>�	�-p˫�7��?�]�
O�KC�bTڽג�J~����O�8�8�6Mdv�\�?�-��+YT28��<���sSOV% ]I��Ϋk�^k�0�@��2�ҵ���nf�	eHxFj��a5~�[�0�p0nR����w<�i@u��Ԉ�`⩥}�GѮ��9n�J�����"��;���e�#㪩�,(8�Ȥ-��������yv�|#4���������8�>��Ѓ�2����L"h�[��0H�ϼ�D�@�cê�ς>@��������1���8�å�"��F��MMǷ�/���L`6O]u��2���1Nq��Ԓ�ŝʍ�yS���v�_b��^�J�Y����c��R�!Bz"��	M�C�8�^����ߪ�r</�q_�0�C��*kB��O�b��	�
�#&�qv�����ZO���d�m�����\�jy�K�hh��x��n����y��l��QF����e��DN�nL�;Ąn�x ���R3�ow��"��Ō�ECo6~��O���a�ޭo��v�ϳ��
��d�a�垓�h��G�8B��D�x��]�Hn��d�+�����sk�b�P�,JV`��4��Y];0�PT�Q�$	|�$�0���K\?�N������u��c�^�
x������l2��
v�W�����G	�� ����r�n�����b���$M�":P�%��i�a貲C���D뮥6rr��NLi�3���T����F�9\X�ޥ���t5�K�}-M�b�+ebau�7[��A�s�p��m�����EÔ$I��u9Gwa�>���%.>D
�_��%=&������/ �E�r8|g���!�!-���e�;9��PG3]�P�=?��;=+k\����˩�u��2E�����׫��43E&�1�x�8��w@�?V�L����!&��:�~M#��\�A3紋��>��ո��"ӝ���Hv�z���߿��RxGjb�]�I&���8Pz ~i�����ج�\n`�nd���&�l~x5(���܀���c��W'��=�!�b,���;�Bb�D�8��9]߯�X���g�v��C�H��5&Nj�>Sn=W(�n^���B�Ŵ�	��vO��h4UG�����%���`��f�!�K�c�W�����G�i��C�Q|��s�#*yD�J���2H,A���V��)Ҹgov!c�[� �~)��r�η�q��Z5���%��D��s���Gn� T�G��[��dL��c�~$T�\�ı�"�^hi?u?��GX�E��w]r�MbÓ��*���� �Vl�'t�7��]>��C�@r�Ƭu0�a޸w:ϲ19�O�~�ތ<_��`��|��]M�.���Z2kN�\C��9Bq��6�`m'E���sA5��pV{�cKǪ�K�+�H9�yL��5�C�R����IJ*ۗ���n��:7H
�z`G3ςS����Bx�!-7�'��	`�\��"3Q�M�B#��;�l��?�{u�$�s���>� jX)��j�����p��{ə�jk�xKkgM�(�����tI5���$'���}���)�j/�T`ˠƵ�29�~�w>���.=�hR&�c�Q�͎�Z�	���1wb+�`���^�#ߚ��ƹ�&�Z����<yZ<S�� 602��"���^�G��y�9�IGP��c�;�5{��9��C8��(�d�׸%i>mF0bnM<�T�ޛ�{�����'Gq�1�,|�RE�hdM	iiT%���^���5T6����\�"�NH��#��ȷ��Z�3�����uI��4ۊ�{
[ִJ�:��dI��O�V��or��s@�E3.�J3τf6gZ�y�.g=��`��PE*�x��.z� ��ơa��(�kyv���}�2��_�D�suO�%=�l�0Q�JO���L_���7l�J�&�W�cY@�y��ԍ3�D�p�CT���+9l��s5���M��ƕ\d�-aR�;���Y�7J����+����2yV�_�+*qi
��S����Ji�"�Ƃw1�TA
�W����?o�L*���m8�{���>��ȆC�̘�ixpQZ���y�o ���26�5���Gb,��Wr���6D�vk%�xOǴ��껶)�tx
�
�h2\��ٴ�wf~Ԑ����N{&Yu���@x�-��cmWk��E�#�/����U-��j� X��ʲ�j�|�g��٪�0Z!b���n�k/�Լ�_lN���ы~]	"�2�Ƕ��'� ��^>�z�y���Њh���f�~�e{�=��df��[)��Zx�X%��j�#k��tK}�I�uQ�}DL��E�d������U��Rx�Nʥ�2M`���9hQM����lv�	\��<�
9��A�:�<��#�M�Y��Y稠 �גr>�胺!y�R
�*����F�G�r_3��Ō�U�������M�i��a���itl�}�~h6D�2������R�����jn\&��9�ڞ����敿*�yҠ2�'�];L��{����90��6��sz���f��;�:^4��%e9*m2��Q��dL,�H��nh����@a����ݚ�Z�y�P�͟�f�0Z?W��3��
P�"4iZ�뽂�Hɤ V��:R��w� ����&}­9S��C��＝��	c��H]\��{f�O>~��72s9�Z��%H���Ȑ"���,Tpق���O=k'��o���5��:�<�~cLu],�]0��Ԩ����)�>����ЮD��{��vw��jf`��d�<��gt#KŉSPX���_#fb���Ho?���L�މ7KW��q���t�������S�p���|@py��̫�]/6p����rj��Rͽ5\��8z��׋�����J��3����t�k ��� *x�r{���q&�������j�u^��C
f/����ݮ:�X/�yiX$]��j�'.]t�@A�_Z
,�1l�5��Q�������>�ƃ��؞�tDY�0��,�o���<aʧ*���)\zK�Q�#�-7�@<g=%���k���%���~޽&'��ev��*i W U��E���f���&S����A;�5;�����f[ �ܬ�+��h@2���0�ĭ�5�-R\٬9A�
8,�Ȇ��O�6�t�<�D4/  ��ܔ����ܝ>(��vw0z���1�g�w���C
�/2��&1A��3?)�OcD�" q��䓶����2����O�������s�������� FTT&G��I%��t�2��Χ}_-_�AU3�^�B���_�5_*'?r��e�Ƈ�1�
:���3�j�J��q#�����lQ&�l+�bGͺ�hGV�a#��m�c~���^�iR��Ѧ��r�zKF�����o�^&��,2��ow�"��\fKE���8aP��y�d�c��`x�� ���I�CB�1��M+�rB�?�z��״�gXe��C��:�XTY"ɏ�6bh�z���L[ �W;3��J����Օ:�{-�
�Rc�"����^e�nm���wq��Y�Y�[f�\��K����^�0�I�90E��U �ԓ|������#υ4��U�q��*�7�x{�z�o,~V� ��`�xyQ%aD� g�B�b�!���5�-c)^!�3�vK9	v�����?`(�u�|��l�3k���/*H����\mL�a���f#Z�.q'��7w���K�4x!w�9P�b���J�Ü+�h�Sd*&ÐYG�i��܅����p�i�Y����w.x����//E��Uԉ<%r5U<"2V�P)�h�˒ W��w7���M�im�M*g��mh&[]S���,�"�����ii��6P�í����U�s��b�+bY��W,Kv���/��ȱE,?����Bf�$��������a�n1PaA�;"�Њf@((nh�F5��x7U����?}?�n��1@*���ޔ��LW	),��g�?%7�(�/Vٺj[~V� /�[�L\�=h�<o��i��5��������}���%c��}P�F��p�v����RP��P��ϕ�a�eH[ܻ�d���؇��2KaQ�?���q��3H��<m����K�k��Ί�S/�M�+��g}F��p�ܲqRT�K�c�ڼg�R/��#^�e�q������/��~���-��{.�����3�����X~U�_nd K�B˼��^VgRn(��f�z�(��00#�U]�u����hV�K�;���9���_���D���E���붫�]��m�bZ���9p�X��z�������I���~�����,s>�$�6�y-P���A<��S��wB���O]1f9�-��2��2�_;+
�����Q�[ 	��0��%�,۰J�\dk�mu'�:u�$
�����UAf����
�u$�<ɮ(�Y[f�tc���$8�o�GM��<O�����'w�4~� �&��R&��R�����M���4�U�>5����j>�����؊��c���*�S��%�Zt��1)�G�(K���j�pUM�F[�E,��*�i����5�*�@~��r���j�To�8��q�xe뵔���I��5'��i*k�����<�4�
�K|T,��%�����+ ~*�sW�1<�Ēe�:�I;�3��z���c)��g�/����oM���k��_�S<��lEN5�n���Q����:8�gJ�*��棲����
�Q�c��»�wԖD���y΋�U�nb�c����)h�Ǎd!s��O=��?y)��B��UL���T���M5��$/�Iy~��%�3N�A��W ��	XI��1������p��\�V�̪f6��n�x�S�3.��'_ݛ��0d�-9�7٠|�� �Ya1�F��Lz$7���V���fHz�zƂ!�Z�ꁀpa�;d��aƷlAy��Q1���z����q-��})R�SI��C1ed	퇔�� ��1W����!=�FZ��Ҫun���彲��&�is�E�4ؿ��1��ᘥ��bI{�?M'����Xӏ��F�!b=���A��\r��]���߲_�iW�LÂ�5�'�_�ӿ�/��P8���P�����|��1r+�8����!�����?�k_�a�Fv��F��:{����,�ɕ�R!��^|�����uς�̂��i&�+X祃�Gaءr��v����=����r��e�(�Zgu ���{��3�W1?��"Nҙ�a��8Ԩ�ſZ�#!}6:H,��i TC���K�":s!�C�V뎊rB�%�l���hg��a^۷O������2�u�1�f�̊����~˰���%��\���g����1��B��2�ء۬j�b��e�y ��bx�%�Ɓ6�O��=R�	��WF���'�B�܄d.�q[�9��x�!k)���tMG{�H����	��P[B��0�����+RN
���"K`��~Fʤe`#wB;���*�[�/\�����w袛<�[z`��ۍ��6d��2�w��KT���$�D����gm���E}��$�����q�J�[�`�q��@����%�w��6��!(kO���EaU�o��6ˮ~-}���N����y�#Y.|o�!t+��k>q���?���)-�pw��_��}8P�~�����&Y���y����R��M�w@� WI�}�|.jc}��D�'v�lj��	�+��0N��&�cq�x���4`e���b�8c��5v�Ȟsώ����vK.���F����Q9�Ѷ��t).�x5�t~��ݽ�%U�*K-�P�.
��X�w|P�O�,9~��j.j����}��/����Q�Y�ʸ�9��5�� K�I���ӁAâ�ĴrĪU�Xl�/�f
ko�iO�����ev���}��8�ħ��X��~��"�:m�ܲUҢ0�+ăT;�Ӟ�$�"�`�i���?3�F�Vˍ����k1�8��`�n�Y�s�ٰ�ң��{�]��R�ϸ�{`9�
W��Tq�䈵\���˾B�j�<�Q�Sy���-��TQ�n�����y��+r��r���ܔV����OӨk�<:z�R�y\�P���F:&^�m_$�%�!cz�'L�9�N��-ۻ�,R5.�d�F�]@��
ɬx��>G!7�4a�����i�
� �T�#n��٠[rð�3�����=�ѯ����cBmUi�`l��q����n,�#ȗˀ�4�����1Dva;�*R�>�1�רi㴽n�2K����e܇���K<�U�2E���.�J�oUA�o�#��ogb� j`it ����j��!����Ք5��'@�Թ�G����G%�3<��倱5�G���D�Ku�jc�^�MϞ�P�w����ǭKa�*���l�`�\����Νm8qJ������V<�Z�� �03���ᔺ̓<^�f�۰��h7{�n{�����{6�&��5��^F'`�r�O�+xƯ"Z����(��*a�����?�v���S�e���^��Mn,k)�/�����8vl	��HŠ����D
���K=����ur��#����୵�mդ/�T�`�
�N/��cښ���mmx��`����*"	ޠX�.��C��nk�sʓù� �(��Iɕk>��Ky�pcj`��ĄJ��PP�ݳ��B-�C(1&JQ�iH�	,� Q�3:D�.��"[A3������phU��w�8L�?D'�=�d���K�������NW�~�OG:��Vi>�5x2LY�J�[�>9#(j�"�ik�	�q� J��]v�IUR���8����/���緧�k$|1����}����pfSA5QB�6��K�-j�����:�ۥT��c~#��U�,�����HY[����?����}Cs�yg{�9�/tӋ,����IU;��JX��A��=�0+�mB�b�U�Jb���9�gc�w�!�'����C<�v�5 ���4�C��������Q�#2@
� |�rEњK��A٦�@}'�QKQ�i!H1z�����ɸV��+��A2Z���� ���0D2���t��AN-'4���(z)�&+*�Qm��)R��W���	S�>���H������A!�����Y9 `쳗M@�8���h1Rq�4�����'�/�.��~H�)/ГH�4����v�`Sȣ�9���Be�����gs�P���lS���LM� ���Yݫ�P_Zw�KM:+|V�@��x�2��"������Ѓ����e��}��o$�v�B��H3#%�tz����s�����E
����~�<��#h=W������LcT���5�)�#��d`q�E;��Q�9E�1IX`�0�eU5���I#��֋����L��8��/g��l"Q�T}G�]<��J"֦�w�Ymۄ���l
�����ҵ�}MQ���!�_���#���y!��x\q�r�9���9�E�G�Q�4sm�_d�r��d�A�Ȥ�[�$��,/qs�eW����b�(eg;^�++���;�$���d�3��]�s�>������FfkMz8�8��w�z�zym44�+A<���D?�O'�����s��]���K�I��W�H㰋��l!]@���d�u��H��ǅ|D�|Į·)�	�nDqf=�(���MI:C}:	��/��{���ҷ�Cj
O����|v��b�`MGK�!��lI�۷%�)r�G�>j�喺�]��{I�y����?�fs�_~p��g��c��os��L����<Kß�b'qb��G�
�uȣ� b�vM�s	�]D?\LU��i>+���e�(�|�0ҏ�O'��R��%Tݟ�A���¥�d/ɬµ���m��,
���������*�X�H(����T���[�i�W�o]jkF%�-��l�bč���D.p��܁����W3g�z��w\MO4b�[���IAB��a��j!�Ox�=4����*@�F�.@X��<���~S�ʤ^%pt߻Ҽ+�i�[0�
Fy���}��
/�h�wq��w���l���C#���}2"w�UlP�e%oHz�u�6{�`��#����;�պޢj�0��1G*{\���5�鱙�l�	�&��^F�! wĹ������͢���jI䍐F�)��	���b��������"�q�,���K�	;E�};?���܍�?K�i;L�y	���V�?�u�7�`َ�dt5���\ƫ�C"�A��n�|�͹��[(D�U��,�3�q 4Es)+��Br��r���1�u�k�Q-à� H4~©����h���i�'��_�'����8`����m���"B���/�#kT����[D$�D�c��6-��Y}'�].di�Y�`�
��c�X���$�Sgy>�����[�6���8��ˮk�-긇gѣ���W��O"�8����{�s^�#+2������,Sp��kN�)�b��g�<(�>����<�q�܃��!_��� =s_B��J!b���&w�9�Mf�F���O�b�C�:Z�e�=	�A�+�GB������T���@�K|5R������F���9'-��W3x��ǒt�fެ�bfLlA�S��� }���O���`U�J�[�W}��05���`��-�&]F�k�t;��0*�����i��n?���5���3�d,1���0��UQ��{���0t���>O+�ş�*J�K������^ޢ]���g��`��Ƨ$}��_���sl`s�a.|7�0��w�7�~m�㥲��pXJ!��cG��KpA8����ߎ���:L/S%��1RK�w�
/����m5�Y;7Y��:��c\F�Ȋ_�3�B�&I��$�����\�v��ƶtN��j����[�-�tv�+z�!�cCB�h^��b2�U�0x��Աݼ�'j�f��4�|0�����M�^��1�#�z�-�<8r���Q<��<�p�"E!��E�2�z)��{G���N�H��>�A��/!�s9��T���&�߀Q&A����7S`�5�k��'�Q�m!/�W�n��:8�O�j��,��g�7����_?��x��:N�i��IhKh�;I���q��l�Mo8ȉ�1׌s��~�p$��@d�Q���q&�/M^����睐��n��nW��T�0A�������nrgR�Ik=���t�
��bf�4<T�F��ug|��WKY�?�3z�)v�^ʟ�]Vsǝ��*���k��[}ˤ7B&�Ru|�s�������f}4g�u��G#��N6ʈ�>��s�J����DHC39�̷Y$���xkn����B7��y/ZA�C�M�$>���{�5И.�4�u�-�+�����a���aa�K~��H�"/����Ff�=���/�O�ǱI��%x/�vMp�q\�!%�9�ԗ�!���΂E;Xp�S�3�V�tf	�BI ���N��3}h���[�t�kֹrC���&�w��F�Ɖ��+�D����A�$!RX{�6�bHXz&+ �k#>�%�~yZ�T�58��b�e�C��ku^���L������t�6D8�`b�A���
𽶷�p��*�6S�2���G��<���N�Ū+�����r�o�«��G��� J����Ҫ���ш�Z)6
\�rShBH�'�k����s�+��[��EAO$	� b许�`Оr9�uc��2�7kw�äf����{Q0G> ��/��Q�#aw����A��DI�3��WOθ(�/ڳRg���䳦ԁ���`ѡ\L�Z�m�&p����%�h��*9D����ZI����|��P�'������H�s_��4��?O"��{� ��}Ϡ7d��)2��=�5`^r�����雑%+�����s0���WL���<H\�X~�"�©ӹr�<�0���+��{�g�?���`*��2t�n68����=tJ�r���vmN��4�<�qa%̬��Yf'�JEz�Z-�-q?L�N�k�\�{��l�����=k�M^�amL<T8ٕ ��������7OpE%W��T�#���v�q�ں�����&�V��՞�D>9C�R��I� �_a�w���[�gJl_� ��hJ	ְ!��E�̛F�������1D��AҎ��=����X����ҿ�l�m4lzбc]��\*4e��Kc��OnF��z+�<�P��e>���W�1�ҋI	5�k�;f�^��Z�B3�c5�h���c	-X�^\�k;�G�s�wK�zǒ��ɲ����������3�9g�8��<T��V�I`)82�֋���˥7I�t���B�6Ҫ�n�B|G��Z&��5H�"�~P�z����wf���!ܯ�]��u��I_�#]���/[@B��j�4�6,#<�b�F�⏽�&8�2o���-���M��ZT1����~�#xbO~�a	��OV�;�I�ب�B�A0�a �9d���n�N���P��1��n�}�TC���� ~�4O8焎��OF�� 1.�񣉎J8AE�J���k]��)�.��H�B�8)����&�O��;�/�惟7���Ev���:,���B�z7�T���.�!�W4���3�����F�v[ '�л$g�BxI2��dmX���ٟZ�n��f׼��A�ȵ�vv���N	��w��s��eRv�R�G�
�p��7���KΚ�C�ٺnF�)���@�2hgY{�&͢]�Y0;	l'גu�KҔ=�9/_���F��0�(?=�6���b� RX�wr