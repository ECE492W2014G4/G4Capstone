��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P��v�"<ߞ��&'��k%P碶�R�ӣ�sĞ������FY&G��n|s���<f79�Q�fLjG��ԓ�H���Hwe������	] ��͔��>�y��;��Z���$dJg�h�_�!q��Oi��Mֺ]�]�� H��
����{GHa�	���[����vb�5�s��`i)-'��N�{�*���4S?����R�#��;ϸ� ����'ʏ�9_�]���X�&�j�mOQ���9
��^�o�v8���RVAW6����&Y�����ұ7���i��d8/��f���KR	c�I0�j�ϲX.�0�nX���E�8�>��^�+�+�1|��J;�:�>���7A��3hr����?�Gp�-n�o�Y�yE躉Cdf�ec7"l��RPEl|�I��g��"�2���5�7ȧ�7'B�Џ�h��փi���|�>��[Zbbop�>��2�ڊ��."�vc�-K7!�t��ӇE���_�S|�U� Da媮���Iy�	�D�_�m�������//��!�ΤC�
��)����> 0���5=�;��� �q��Ә�W�¹TH��H��|H��D3�}�A���I~�;M��@��NOҗ<ܵN6
}� �QzfOVY�3��{))���,��28����Tw�Yďz�u�+��)01A*6��#���̖O:i5��x-X�9�v&0\�h�ձ8�����9*"&G����:U�k��g��8+RmT.�%��j�(�r��=4-��	�S�I:G&e�N�c�p��7�&��/�o҇��-2�x��h���kx��z�s5�eAV���E%��y��0C�W,g����^@�i�`�����O27��x���݋�b��M�uq�$�U`<�>%c{P��F�I�4+�������D��q��WQ��t�5:���Gw.sL5���jijkve�����­(�d���'�ņ���?'�I�4z	K�`MG�J�l�oGH�btn� K�������J�� ��H��%���7�x��/Ҹ|��"7�W%
ځ[���)8Jᡬ�ʹ��";�F>��>Lzc�bA@��q%�|�������Hwl����n�H�J�:�h��S��K�Z��Fm���vU���.$���y����V��Qm^4��By�%d�Э�Fj�k_�B ��ˇ!�)vj�֝E*�����DY�B"��k��86� ��@���p�Y����%?#�w1.�c�ّ`�<��"^�g�����|�;��������9�R]�	c�  ���/rn�����=�j�����a�\�[C�NȑuG���ls�v&����PQ%�Q��Bo;���B��ۑ'������>��e�嚻�^:���3:�������<(LTg���0h���̰_�����⚗`���o�>yr<��"c�8@>�E��d�i-��"��]>��aϦ@�L���klP��|�Df�Xg����;����r�s��BB�Ùg�"O��J<S�~��<J��
4>���Yɣ?���*����c�26'�����m9���1n��:�-d��s�La�C��#!a~Vp�7����1t�/Ȗ��>C���H�~M�h�&�".
�E�V�3$i��E)��j�;��k�f��X�v���2���d&vz�
P�ގy��h|��'
XD![*�i���X^�tŚ��5Z���h^�A�r��]�f���,�|�T!�2��çޟ��ƕ��wDX��}��2�W�>v�_�D>�A��m��>���������?cH���{T����T
�,Yg
�|n�B}�~:>Y�(��2���4J$T�x��a?6>cc���G��i+���1r��х���U��(?��k?lE��Q=]�*�]I��~݇��݇ͳ���cs�*JA�W`��<m(�K�uP����N�&h鏈��35�8ݑ-��`�"����:�9�Ӝj,ӂ�XF��L�*
i�b4��+c�;�I����\�]-)�}���Q� O�!#T2L�d�݉\�1�KҲ��*<?D�&�l��_i |x������$�(}�o�VǶ�ד����V��e�#�����u`�&qz�����]oO�(�D�h� �U��5}�vz��{`��d¥OX��Z�<A���[�hb<�ֻjeE��ojYi��o2F%j����U��3ŞI��}|#H�i ��!ϢsY��?@��A֋��3�n�����]��45iu��Ӆ�%����ۀJ����I���[/��l���*��� )��5��a��������:��"Lŵ7*%�#���0Nt:���w�Tlv<�r&���)� �{�#2k�l�[�a�{�>���J�;QvL̜��&�y�uK��P��/�)(q8�uٱX��)�|X���7���e%��B�y����9�X ������P���(.?"�ޘ֪�q>y�!���)+��Wm��2N]@�l>.
��1,���ԙjϪ��W�
�RD���>4�K���q���P�JVC����l~���C4�����#N;�-�����R�%�k�DAR��V�w�FSse�-����z�于z<��(�N�ķ�t�N�D���şA��:w�.�u�I���0�ە��gKf��'d�G�5�\n0tsbK���#�m���?[��3Z�����[ox�<bK+�6�z��љ��j��Q_������s�Kͬ�O�d�re�DG�v7�P�=K0����R�������@-�]c�̤~u�#H��Es|�mY�@�]��X���QT٘��Ӽ�0P��/�H�T��c��FqOR�/����?��h̵{x/|1�[V�QU6N���6�*�Gy�z@�2��yՑww��i��B��/ѥX����ܪ��t�ji¨`��4�)�����=�dQ�+n�gԥ��~�����[7��W3���#�2�X�`�����*�ԑؙ�8�L�sb!©aRU�.�˲�8'%ъ3	.0\t^����(�9]'7�pJ��vq�����,���F�ȻM�f��ف3�>���ڕ�}ц�@]��_��S����}���T2��W$�-�W����Js�������Wm���]�A���G9d�i��%@�+�4gH(/~8BJȵ1)N��	��*���',R�c-�����&�W��w/[[p�d����An� Tp`@��@"��O"Ҭ�P�;�I^r^����Vf(�i)����k ���@n?A�*)#����:��g���5
��<$F��-��/I�Q*ڟ��5W�{9��|�)5¢�9+oU�p�CFͮ��Ol}� E�%7`3�����S�&�)��N1)����[��	x�/̷���I]����
��SS�{��I�3wd���_{�v��?�z0o���-0���V�ɘ�I����K���|�>"Q��!�#�R����h�4�<��<�-��E�c�2Xſ�w���n�2�ʛ9 �F�g�9�W��6tR�{�f��|��#���hޕj���]���g��ɚ����R�ם�����H�@}�:�[Įb�񋣺�+��RUR�eG�$��]v��0�<gZ�~��Jl��������B�1�|�G݄�5:ǸQ�)3/�#��:<sP���>�Ԏ�p�A��.�X�Z0<R>�"��8n!`u���uMMo	C�ȔZ@&�G��f���A$�8����y�o=�7�5m�-�E"={�����A/sj����3��Ҽ8 �訆��:M�"4��u%�q�u�\]����hV ��xTA��O|�l�3���Fژg}���c�L�8�T
����1�t�;T�*�&�Va��j�A��	98�
)#er��,�7_��9��g7�f>[mI[+�����<B}���Q?����e-@u����%_��i!~�*���N���bqrf3%w�(�K�F��w��s7��3!�(,�d�噱��u��.��r���g;����{��l���Cܹ�sg�`a���x2{hV��ך|�-IE9$s����\saLf	q!����d�)@t��C 6=g��Uw �\k	tC������D����R�	rLe)Ϗ� ά.�����3m����z��ɑ2���#;5T�6��ב���)�o+���%�7ƹ�a8Z_�Ņ�K/�bו�L�����n�<����Au���X�4بw�D�u<���T�?m���~߂�MN������D�_�v�����sل8�s[�o��[���\������_$n��]��t��T���V�������_V%��A{��ac%-�\n����.��!�?�����ݡؕ�5������ d?���~a�U�R��ړ���$��7q��������2X����j�s��l����1nD�׼���x�|X�lG�cG7�����ˠ#��K<�R�{�#�s�C������{N]�����Jp۸���!Y>�n�j��~��>"~���Qt6|Z^�6A4Ψ]xc���es���6��LL���8��"�=^HFW]a�&��|��{J�����X��+2Q�2�w7��0�%����]�]��(]\�2o�]jf�E��k)f�&f1���Z��G��(/�6J���qJ"G���Z�X��gg�U��h'Nz��K�%�<�4]?�]���6���)Nm��#��/!4塬������n��0��X�Ka��eUe����kfO�|'A���&U�s>��#�N�.��-|�<�*]p��:��m߭�?���}l�vָэU�w#
xP���_�©�� ����������v�U� ��GJ��I��ȋ�4ߟ0pd��-��FoJ�9�#�p��(�s��֝lgP-'4��8���"H��yT%|�L��86ܱ��MSJ��O���wN�g�nj]f���&���0�ᲆ�7�T��!B"�B.mU�F�H���� V+���h�V��IrFd���%��,i�����[�Y;���_�}��e� �)z�}�l��x9wIF��3iE������sBM��Y�!w,RR���p��#��wOg
rWgtA����Zqk���{�Gn�| G��w�*�ÖRE�b�� ��U��C�
�~��~e��a��x���6`�
*�Ih��� ���p����{âaR���A��T��UQ�`��� d�c�2��O]V� ֘�[�F~�)�<��/��Si�4�����j^����:e�O�"_	uA��fR[�D�2)"a�JK��/��h�Eb3��]����́���	��x��"/E����ƾ�d���f�f�e_Ka�����t_!L���N�N�<fxM��ݝۉ⹗ZM��%E�������r��:�ޔ�#�׌ u�����1��(��<�CW#����p�ռ$����	chO��H�ȉ��,^��y�.��EkM�Rw����Y�i~�0g��g�u�-��\�lm5xq�Y���b�Q���g7ӄ�b��yn�N���,@�Ee��У�)T&�ň `�Ҵ��a�H<���2!��f��܄E�F&��h:��H���gF1�h�3�ߓ_fN���E#�)�� y������vn�O ����m�9(���(�-Z4 v�%/���b���2���߇����G������U v�
gIJZ{h�D=\�/y�F�d���DN�b�}a3�^��:���ʳv,��'y%�������2�+C*���ōp3��N��S-�����N!�}O��<F�;�dHC�$���(�&�KuuP����l���Ǘޥ��\j�E
��Q��)l�<��	W�Ua3G������'"�>XB�$����`c���*��'��O1?߆A���Ć^���x[syo���s ��j-�流�5�A�!(A�J�Hc�+aˌW(ZA�t�S�н�)��)0�cT�K-r��~r�k��[��䦊/�"�����wTԝ��
M�(s��QؤоLR)�<�A�*��B���Pz��s�F�JУ��s`��p�|
��R�DX�&j1Զ���5Ëy��ʡ�õ$f�:K^�\Jۤ��ᄺҰ�~���ą���?>�M$
�P���x�ӭ���n�S�W�=�/ח�ݨ�y��A�b��]M��yw/���=l���/�<����w}h�yy����`1����17�W�Zq'��v�_�`-��Ȇ 5+�'��m��H̭Ͱ�C��	}���x���"	:VMI��f��k�M���Ɯ�}ku14�#��ܤ���ߒ�����xW EgX��B���-|�Ҧ\lc��C���$�/�8f�{n<�-k�b����e���*~;_��x�v���]���H
<;` �1(�	fjS�΃l�Xx�$]�[n��H	�qǘ���n���rt�}�g������<���q�A/��L ��lm�������������6\��h��֙�&m�h�)5��n,K���P|�
�K#���b�B���U��m��V�o~��s�������]��Șzk����[������Z����h|�ȭ�ܖ�`����:`u��ԽY�n��$/��d�2gD�4���.����u$i�7|H�!N�Aug;cѹT�����'�y�握����KLȡ�E#���8_>S}���3m��mWJ����ǆh�y���~橷鍹���HO�O�I���39{�8H�aY�p	ݣa� sU]:�yA�Y��aӪw��L�>�<�{��\��	��΋_���iY�@Es�em "Ef׊@U��;㼂]H�u��GN�7w��R!�H�uxzە&&tٶ�iK��T���?���ܠ�/kna���puv՘�0��i+�����
����4�ƒ}~�(�_Jѣ�X�"��H�
B�*f��G�`)6�X�"���ک&<��1f���NP
ޚ��R�$0-��k9�x ����V
���w����O�
U"��E'�1�[�	v�܀������w}KQ���??o.���.�8Z��{"z�?���s����S�ً �~��`�5�wP� ��tD��qCUx���odF��K����r팕I���g���(��\��jx����=�\m���}8$�M,�h���D�Gea��	��i�C	�׆9��a�}^�r�`W^���c��מF�A4��ĕu;mԥ�o�N#n�~u�b����O�[ʽ�]���%���mzw�A�~5���8|��,�wVi����y�oP%�6͹�Rr	�����
�oe)���&��b���<�Ai�u|����T��"�)�`�خQhps���Kt=qP�t��<A�p��(�P�+�5��3I`�uPm�M��~F9���4b9�_:�����ȵ��et#���oq�Q��D�ۚ�{IgL�9m<��E\�%�bT��`��;L���t �=.��	\	 T.e)̇��xB5Jz�-�Z-�mػ弐)�b����ȫ��cWԽ��r�t�bez-=��5�24�s�W�U;�^Rcg����Ve:߭Ȓ:���cș4i�F�)A�Z�{�#~|@��fm߹�/M�lҡ�����
�b>A$�����J$͑�9;z⵻K��"�ۅ���`q7���_�9;��H������ԏ�@-C���N*܀oug���u}��z&�pW�q+`�^A��:��>d���D��G;4n?h"&^GA�Jf1�t-���٥p�w(�sƧ��&J�l�Ve��7����yik�z0J�v[52��^��G��R��597�v1bw�����V�QQ{~bҸA��	�����cr��X��4s~��o�p�8�ΐ�DD�@R�;q�X]�휅�_�
�"��S�*��r�u��Gw�i�ig��ΐZ�8|Z^-j�j���^h@�BȤ1_xr��z�L�$��~Pd1̀D�pf\So��g�6)�rU��i@w�����I�~�:�&V�Qy��9F+;�L���qMI��b��Y�mWe��Y$N�,'j��|�p�7��"��^��Wh��wl��3c`Ft� ѰЦ��|��x��R����vl.�$TQ
jm��#�:M$�-��`��X���UbH̳����(���t��E�Ʒ�����N���~������� zn:E��mw �@4a�'[�/7�dԑs�1���餝�� ���6������(��M���ѣ�m��A�x����J1��H��A�{�C|V��,ϙ�Iq)ԉ���K���.BB=�dS�q]��y���P�+E�Ra	)�-�z�>$��Ԣ�V`8p���i�x����\�c��@J�߬�G�v����M�Qݡ�`�{�A��]�J��j�ڗ�6���N��kP�U{�Ej�,8�,]���(<CŰ�j�j���� %-ȧ���^�s�)������<�C	c�B�S�AE?=����_�����m�PGM /j�<���e��$"�++ߏ�����=#��Νj"���j�i֗���ډ*���!F���k%W�Z//�1�<P��� \�S��q׫����c|��Lx/\�1:�O��Z�a��_�7�}�`@8�n �=X��壂¥���J�Oi�L�¿�yN*A�sĞeN�,��;�jފܪ �N�[��������������Y��k�Ò��0���<߁��H{�v��S�t��H��X��f�K�Sx��Cig���S���oep�d���3�	�8;�¿d�Z�p�#�ǈ��`lpΤ-Q�?)2�5ª�E�!�z�.u|}Vj�T�t�r�P���\Vix����6�HHx���m�l��2��=������W2{ U|*��eU"�Ξ7�bf�/4��JV�d]�J;�6��/#��U�f��s�#�*;	)�QC����kg;<G6`8�]..�Q�����Z S���gk�B���a�5[{۸����i��"�=)��\�I4���O�׃��#���m|���j ��E�Β (@u�@�j�5�_1y�l�pmg']����w�X����(Ҝ<�G�c?����E;�}��&?k^ �ך�	��'�������Pgh# nt�I�d �_V4�'8|�" o��7<�Y�XŚ�I�=�CD�ch�f`Ь|��W�FO �3'r�R�*L�F�@��DK�F�Ɣ��>MˢLI&��3ê��?"�R%4̹]<0�2 2�mo�̊j�&^�E��=:혱z��(b3�0�;��+���`u���`��I�I��p��1E�l~O +&���|�-HS}�F��hn�B`)���j������]�01�$Bjr��P�_j0{�7��l�5��i[1���i��~�\�;��g�)��xŪt��S/�v������`�z�O�)���A�▂ף�/D`��l���4_[�)O{9&B���qH7?�g���iF��3 bU�n�N�G�ݰ�?�h�������+��8P.�mF�>!��`�w�?�E�� �[�u���k<	9T4�x}�p:�&t�F���U����RɃ�Ð�Nzs��l��AZ촌��5%�!�ܭ�W�ELģ�}Ei.�X6���-��-ZZ��˟L�;��<W�>��Ȝ�f����s�����*A�e����kƽ�u���G�q�Oh�H3��#ڗ�t��I
�i�cn� �y�d@���b"#C��kфZ�}�0�̾Aʇ�������~��/�<��<B���"�!E��ߕ2�F�	�K����8%�'p��ֽ���z#�"�R[�)�?�R�+�Y/1������ʧ��)t?��*A<g�}^�oU�1�=jS`���JT���QJ@��P
��+>X`kY���Ļ(T̋����S��V̓=�2�7��:w�K����5 ���!Zc�J�[؟K���o�c��W��ܫ�_ ��+��mbw˻S�xw@M�]qkMN��н�_�{&�f��7�
D�̜)-N�Fuڋ����.�e��$�1z~%>���5E����:Y�p��F`�R��\w�1��0^��t S�L����a����`���.55B�dG�QF*�ƶgԢ�'�������� 9 S��/xh�}h`��b�: #�̛�E�QU/c�ª�x��牉ҫ(,��c��RoF��BC�wQzB�f�f�������{�_]Ÿ�`�o$_��T,��/�
��o�4��~�&�K�B-�Gf���� Z�ӌ��ԥ�:��z��rEX����E2���*���k�B��[0�i&=�/UD�s����lDaYu^�k$lҨ�S�����|����2� �Tvȶ��a�����z-��J7=��#~�"S�6T+�B�l�,�l�O������q�T�"ı�.%���+[��TH��RT	'�4g��4��1;����@�[��a�5k��)�1D��W���z0��� �"�(��`��Sr7���d͚*s���ɗ�3@���	Ho�����}]*���mCpY �h���cp)<��<�����aF
����H�$�Ȟ`�6�~Hڬl�<�M�K��,��RŊ-��e���`�����j̦Ѱ�.y��X� ��������0,Rf��J��L,r[C�3o?K �V�~���(p����a�BA�-x���?��P�w�/�w�J19=e�p��� ��0��
�-���!õ�?-�Z�x7�����y,��L뢙��	�;@���Ww�oL�h�*&��~�C>ta�ԯ���KH�T�wQ��^S_c����W��"wI����M�'�z2H���n���w�U,h>���7�51M�Q=q���V۰WÝs-�Q1���W_F%��0ڸ뾌��l���h-�"@���2�!��_�a�&*+��I���Qި2p�W��G�0��VÇ��'��#h�$L��FN��I����e5�����Nx�^ډ�ۖ��V�?�S��3������=����ᅢ[\���gp��Q�q�7?]ގ}_�l����9.18�$�(��G����ms0����0�zJ�V�JC��>C�Xt����\�;	�(�L�A<�9��{�]��x�ʞ]�ߎ�MV���N��>���=�Ɲ�~7�2��3�@�暝�x���`s���jѩ���HIW#ò���c�~�۪�_�~?wo���\�S92уK��#�R�"��<����|]9��ɕ,0��\v�&v�l�Uz��0���bgc{,{���Gp�1�;W�w�H��9C��C%���C�3� =xL�tukfH��,������ugj����B?O������f�Љ(��B���:9�r�� |>K��m��U�=�T7����Z��+��t�"�޺��	HƹY~y�
{{|~���B���5����$�	����x��W��ђ��3VcS��R��F�P���m�:@�����	��]�c�>�Ff�h��ȧ�%a��6�^��^�;�H�^)������
:������UGm􁮆�,S���ڔc�|�&T(�cc�_�7����4@Թ� Ő���mG����)ki��U�}RURL�ku3ј���2Vr�`m��Ì��0z�4}�>�l�hX�KVWU�W�*©����NA;ۂwk��M�������c{�t��M�)�2����k�<�Io��	��/��$�Uc5cLh?r+�r+�*=�kzƨ>ǿ�
�/٦_ m�sվ<t��$����h��gJ��<�����ƍ0u���R����PZ5�#�D�Wt�w&Ȱ;R�ީw�~��4Z�� �(N�z�a�	{�90,��\� �t��jC���qm�=/�"Bc�拫��)�����x1��҅B��UajEd��焛�G��8{p�*���@�2��X�=i�fE��\�H.+�B�f�F��Q��(6^�CA�Y4qجڥ]���$���ˮ���]��Ƅr�Z�p,������V*ߎ��� �W��P�JZE��'����oc�6��%��Ӕ;�}�r6`���.$e�J���Ԁ����1�K:�ָ!yG��;����p��A��g���I��T�Ĝm�����o?����K:K�k�Ĥ㳳CH}1�7��lJCt�,�C��.}3�ȫ�6��u��~�j�˦|�(A�����pqDj��;���B�)��\U4��n�p�f�͉��	�7}�ojԡ�M PM��d_E�UȨ9�52��"���(Iq|��aM0��ݩڽ/��Cs�VVˎB8���i���DS�O6�N%O�40�ʰ�T鹙���\�6L��4��,���P�d�.��j����E���bD��^���V��]l�.���aG�o^��k�M��c�Bv��+���o�����mPa�����P���DPy#00I ����<���������!C���!_���3���G\g� yz;@ J[Ї�N��T��
hi�9��Q�5s�_��̜��� l�LmY��[��MY��#�E �&gM���Kc��*�o	�3U�%��;��]��S%�*��pTt&��&ґ����=�@N/�a�;�lZ�a�E�RzW3���fO�)�
�oQX��C�W�I�R�d��]`C#�*K�	���:R�U͋��SdT_Ʒ�	����̼��r&PlʾQ
�oi��~�v3���|�t�[�H	K��Ca�lãD�c�s�I���&F�!+ЪJ���h�m�E`��g�lX�dwt- �Uf6�G3�W�f�HʞV����J@�%��^,��|6�L"��R_a�?�U��2���GQ*��ںmLP�J�޹q�֯���˶�߯�x��{ݘ�jD햣�}������7���;&� �Ŀ�=N��A��%�|���ҳ��c���й1����yfH0ҨmO��?Ԏ��<Qt��"�ZJK���1 8X� 68��KfϫB�p���^YY��t4��w�,W�P!{���;b�7���K����H�'q�$#*Z(�]Kv��B=�Ex���Kd��a��0�y��;Y
��g%`�3����B.'�$J&�����ݲɓ0T�O՟�_�{+>jZ�?3�3=&��?v0�CV�G,�6颶
����8�;kj
#���*�;ݧ-�I:[�3���dt�	�<3�E���F�Y+0�b���z{�qE�1��?�7?�K����JyφD5�6�������|��T<i��,}0�uw�(�a\��q6� ��r���������dV��^^_�{ѱ����E=� ��y��AH�����w�O�s>�إ}G�����-�˰��x����v6M�Gw��'�lh�F?��~�r7���mW3����"����1�=�^���J��o8����HC7(FU8�(��?3�ls0Sl��D!�b�Q��<~Vt�$���R����S�ύ�N	�O�|l�%Cpo&����چ).7���+�!;�f�����H�w1g3�`�w��#���)G�n������u٥�tT���K��h8���+�\� ��A6N(�1��W�4�O��P���O�#�@�1?&���Bȵ%u
+fQ��v>�N6�����P�sq�%�U����C���s+�v�S�x
G�j�Л�tX�(]�W��F��H���(���J�P�D����.�¿��8�eӸ��-61�}a�
�OW&���}����n+#kՒ��p�_tQ��g�!��鎥�M~t��Y�v�����s�R��pW_u5���x&c�|L�s�KL
B�11*z�J���v��g��,�I{VG�h�<�>`�B4��c!�U���0���_T��������c����-0_���*G�傣�J*W=ܕ�����46g�B��	�J�Wl��Y�2C��
}��_�
�*H|��S8E�ݒ����,@0��d˙�U�a	x�Ru�i9zj1�N"}�HKzuc�(T<�QbEob�d�oo�����	s��Gv�YXU�3pYI��'Z#:j<{���
�.��nˢ��m�f�g�AchQoV�׍s����)$��[>j�,n���e}�,�`���N#��L� �,�?�<��/eS�O}���g,.xx1Y�`3ds�}.-�x}:�|	���vŐ�T��y6�Fws��H�b��AKz� 4_v�ft�gE�ؔ%p��$pPv�BRJ��韅!+���MM�4�v5�p�� ��OJm3u��fT>�-A7�e�,�����*Sx�����v���3�X�kc���/W�B��5[�Y��}��6���n\�� |F���h��)��qj��T���<;Ҽ�#Rc��_mG�!��O&�;�ȵV1%��E+I(՞.p�;���	�A� 2�(>�n��O}[��S)J �!�H0�TCC�xo�:U����*�Q��r��ڙݷ@Ӊ�h�;�G��S�5P-�a��d7����P�Y�bd2Ёl����XV�?��w���L���P��"�<�ے	ζѰ%b.+q{�0 ��A�=�f���ow�xε��O���4��'�u�%,�gΉ��OW#r�_�'NE�*C	�F���S$7H�D�;+L[�yldU�bu�d��i�x}���@�X��5&:=5n
d��p�����
�ڌ6�ܮ���ځ����}���%Z����1{zý̚�y�F�2,l̮%g����>=�k�/ހ��V>��~��L��e�v0Q�+�p��~خ�WVG_ ��e�ޗ!��Q�N��¶�|��.��gGÙɕvj`���6�q|��T��|�G>pa�ؠ���B�J>�oײ�PcL�,Ԫ���Yc�����6XK���)ug��؉��h�r!Pm���P�h�B�*!W�Mn����輎�y� �����{eۨv	
ߏzƎJ�nN<H4
Z���6~�f !��
�F{KC"B�8��ӻ�-�<�f���	��#e�@1�V�@���/f���2��x�D�S�7�n�VSv�cp�̚�!������1���H�c0(�L(#Z�Dڈ�]��1l )���'+ԭJʏ�k�g͞� ����\yy�ɜź�P���S+^�V\�e��R�o���s"����V�X��w6p� �
��Ì��H��؝�����������!{)��B4��XD�:I'%�l��W^j)|��7���˄�wadC} �i���/�\đ���~�Ѭ�-�D�'�~��3� ���Kp�n+�)	�5 �,P�@�վ$�-
�=�2:� ��5�������hv 5����i��Ƃ4w��k��<�6�6��
"��ӂ��bK:y:TT��Q@=g=;�+-���냙U��Ц�'*72F��5�M��2>�e�����zM�Р`�j���D���5u�w�m�Q;��L�R�:��P�	��U|���ʲt>Te�k:[��U2cOD_w� :�: �L��i�̢:�$m����E�,��zֺ3���3��5����㶃��~���7چ�P�����O'�{	ʗ�3#C�7�F^�-��^���BG�Q�w}�o�� �XR}����U���5[�^j��®>��}M7<�{!;_-��g���>�PA�p� SR"�|M�TQ޲B�r!kN�D����5�34��W,ُ,�����H�Aԡ�ے�>��h�;���}�r��r�<��5�F��\�_�f�qu��lNiz�y�r�+{]CY�s,qo�ət!���A>���	���6�J��~ͮl3���󧩢��7n�_�z	L�m��[��-0��և%j�쿲���|�j�.��|�5���Z���?��]�,�K�y�>*�1�o��b~�2}���v����=W�Z��Lˌ���F��i��Mw$@Z(_W�lbg�-�SLl�xKP���Q��,�o%���8U�O��/aצE�O��W�
�[+�~KM�<X���z�)��.U����_�t$��<�P\N%ićn/�QM�夕�L�ܐ���N����UP�D�Ub��f�U?�j��Ի������*���Qe�a1�7�s�Nj�.-�G�DN���H�u�TBgU-�4
�;����l�����73���mFw3t�㞁�<l�1�%i�>F��&]������ٲ[yJMq���7��|е�����\q������7��'z�?���I}Co����\h�b��8�f���K勨W�j�m�~����j[ ��
#���������⥻e��w��鈓�W��O��f�]Ç�C�D:^����Kv�T����0�@��:rӢ)�L���d�����Y@D�*%֍h���zf�C�����$^������ǆ���(�zD���B� ?����,������_*�骻�������
�$�r{�Ys��>�����H2%��ĥe<]�ק�$��A�J��n��>���5hV�~2���F*�b�a	"�Pא�6�7����1kP )�˳`�p�)��D;�Y��d\L�1��f��q�>V�qh�kH̓l|E�	GC��啀��wD�����T0%�#�t�� �fv�C�%ę2�����-��Yj�_�����Qd��l���f�)�X'c�Ry)})l�/���>Tg�Q�R{@�ຎ��G�Cp�&
8]�I&� i�8nnԷ��"����T�ϔ<����j�����D�⦨t�a�v�_��\�gZ>!�Qj�H�{�;�����F0�R3�������Rߋ��4F�����2~���z�6.yAr����a���L�B�*��D��]b�3<3����,i�����)�^T���Uoa��ݲ0���uQ���piN���g��I,
�c����ծ4:�]Pb������(=��;������;w�Ι 髵�{����~��j�"}��(}診��/7%m�L�_L�mj%�wF�^n
�G�	�BnFʬ��QV�G)��J�_S��.�܁�د��s:�;צ'�V����<�Uƾ�����Н����z<�����VQ�?nN�Ěi��(�H��#�mh�����
�t;����^)�?[���p'��f'�^R��u�,PQ��/z�TlF
��B�o-Y����3x��z�0�M��1��O��*X�w������
Z"�������M�b��
��!:F�c��*��a�l�)10%ppW��B��<VM��N ����sPB��v�i�˒���p�����%Ro,4���zRb>̊�`�lz��9s�U�����<~��&�W��'�U���k3��x0�y u���{W�:!�g1���}���j�^�P)$g,,�./4]�7o�y�Ǜ8#�w�ek\�K��B8C6�� #D�У0w�$�`��4�������y��@��DfؓǛ|����,A@�֓�T��j8�|qujR0�r�&�cf����{�"Ǎ�>K���@�y�OCw\|�)�F)�3/w
[BKX�bR�zt���Y��4���vG��>��P��22�H��s��������F4�G%`��>��+���0ʅ��;����Fw�x��TV�L��#��< �q��7��AM,Y�8Џ?c\kh+Y��!�rلa������@g\j����'&�Zy��g������T9�ut�*
T����yMc'�Lw �[�;���P�C'e��V;fߢ�8�X%�r���AC�@�����Qr[؊(a��Y��� �-�P�Q����>�{Ջ��ĵڣꬁh)l��:�(jD�ҠdWr���vR�4��)�R�����`�-���oSA�1DWw(��!��O/K%������F�XE#,{]vx�i�aV�:%��ޝ�����3�IR5�Mߌ#O�TAr���XTU�L_��f$�1���5�D�TB/��Q�����#s��;=�:�V�E����E�|���W���l�;O��eT#���8L�~F�RѸ"��P�:�s�'��R:�8z���r��I�.�*�����3����`NF4�3����g끱�3�J�T��FRu��۶�$�~���I$���*���[`����"��2Cre��]�/�<7�yx�|�IV��Z؂3q~��}�X	�����Y<BF�a��=���G��n���J����أ�F��k.�-�r��@��˦�Ka�8Ʒ��I%v.K����<L��<:�?�F�/#��W~ ̨�v�D#N�P�5:�4L�F�TC�@KDR.-ko�5��� ��9�8w?��o�"_��>���c��}5�!Q�0����qi��L�Sɶ����B�Ų�?�4+t���Yn�FGR�B�~��1͠�y��>��l��w��_���|�EJv����}2*
�3pZ-$�k���`w�E�c���L���!�I�3��I :I�����/���2�	��
/8V)X%Q	��K���*n�o)j̧�O���9)�Y������K��j�e�6M�w3��{�L_����;�ݳc:��5&�|b���K���Ճ��!)U�/�vP	G7��&\���:�
Se/ni���lX��#���6����i����T�GhA��5�E4�eiϖĶ7�w��a~`��8�ܧį��)6��٘��#�73Z��f��
��NY�%B�� -��u�KPAz5�`</Y\g�}!M�8��TG2���x�zb�S��ӵ�WK�<?������N�7�揑fo
(,2?E�$&�|�=���������!`Z���-��XvD�z>���\�gS��t���|���
���r�i���	�DA�\��C��"��L���{0�S�Erݓql�RH������I49���8�&�U�������N�I��k)�i�+�p�H=1{O��U�1�7`NE`3e�8�*�74l�|_E	!����w66sԦF��C.~w�S�G�d!M�������z���^^�Eb=S�r,�黈�᥅��w[)�h3	�ؚ�1�� Wd�>CR����{�Yp�dA�Ҡ�=R������X{E��oI�H�f5�~j��R7�{oԽ��:3�[[����ƫ�d�%�C�e��]�;Ƴ��yh�����7ka��17���O�*y�b�*�{e?���5��"0ʵ�I���`	�\9� S�LG�A��!|�ɃieA�U��$�ﺙ�7�[�"V���PwB`��>�"�r����	GƷH�n�i�y��F��Cj���&��{▮�Y�(=Nu����n�Ε}+�'�e�(�oo��"� ��@<(��-f�;��~�45��ܜ}D4���b��_F���;��0��S�T���Q55?�OD�R�p�p�+*9�%����ƞ��.�r�E�j���1��Hv'Į���lH�g�T d�ZbF`�)&�1��iz���3�)��,��n?h������K�۸N���ϫY�q�U2��9bQ���zq�Q���l��(tX	�6��`su<|�чN`�rƴ�ބ�3�3�7�k�[�,c�ER "U���	���V�T2����ȻS��w糌��w�����<N�acGyuE����)��-���[��C�L6|�y���(�GWD
��4�yA`%���=�nMR����o�t�"	,��:���{�����`��pd���FU7�֫ ��Ǎ���O��3��!�F�)�C.g�b3���`}�ꭇIsf�5�eGͺ�a�`���mfr�"�\�}�Ls0�[Y���P�V���bL�n9�V�9�0���;y�pf��4}A*3���}ݰ8:p�kY��>n3B S�S��+nA���f>N3�x��=B5ʃ�M�LS�\$�	#f��"9��&7�W��Bk��߾D�S�i���A�uf����:NFM��~h�)���7�+��H��c9�K�z����)�c>T���lbI��G���;���A���c��)��o�4ۺhAGV�T�����RZ����B��!ˈ(�f6#˝�_Т~͝�H�I�$l����_�]��k*OS�?���(*T?*)�*� $B�s�Q�jf�q�f�Y׉$�,�A"K��f9ֿg�]�%*&�������t��kˤ2�
Qs�D��݊ǯ������Ж�0��D4M�n��]&��?��[��#.-���1f��M�bUo�KE:-g,Py��@r� f����/�.���=��k��Z-+�(��	3����k���>	�<����l�R���K�Nw���_�T(�6]����H#q�9KI̩㞑&�s6��-����7՗��ޜe{6�Ki���95Z�'Tz��vT�>,y��Hw�~-aOk�^hʭ>���3��9��{���/��Ӂ�~$�z6R*�Ubx��WI���fh��i�m��Q1�d�S�^I� �fkp��#�L�r��,cXkR�0���s,��B�i�h.Tiޯ�������n� ����e>��p��wA�Y�[�ƸR+��b�/��t����A��ǯ��Ҹ�MZK;�9~�J:��K�����{�!ր���-��9����׷� ]��4WjN��n�t�b��b���G����@���,��4C�>��7I��4!�k�ω���Y,�y|T�.��/����U�,��/�E0�C#|[]	.-^"%�Ϟ�k��a�a!.����ig�, ��v��q�O��|	�� ��@�d,�(/�-63
�o#:hvtl�P`��S�<}͘
#j��Dp���Zu0���O}<8�W�bY�xX�I�O��f	��U�y�}?^�oG&��ޕ7����RQ��p������ȡ��6^���(oE"��Gqk�ƀ���6R�� �A�\2���0��T8{�A�VY�POF\Iҕ�)��v�E���c�[	�io�c:bA����P^�.��n�<���ʃ[Bj��,��=������m����jn�nm��jTKܴ�P���%<��(�� �d���Y��f����s�N���nȖar�z|Z��֯�����G����a�4i	[;N}\��F��4�8�X�3c�G�_���^�08�f�����:��
���7�c�b�}Sz�x�{�����'�<�Q��-���4���X|=���oP�� ab�:!�L����Q���y=l�U�9�t+����#���������)B����|)W���n��x<��)ٙ6gk�
O�D�]<1���D[V;�صt�G����1����H�ݍI߾MܶM�04�σ��/�K��}�v7�4�oN�vn�f� �[3�G���㼽M5�cۑZ�~(���L
oM�{�������[? u(@�3��c}Ma?iå��G'�T�r�cD�lգ�~�����c��e1CJ��h&(ݔ��+\1�i�)�#y�(D�Q"h���;������M��d�sT	��h�A(��ki�����eˀ6+���+FF�>��0�1ؤP�2M�%ط�8{`۔��f��]IR�ʻ��6*{�T��u@��w��sә\��MBp���6!��2�*=��FbCN�a��-
Z�Ʉ�X�7��4r5�������[
VI�C h�e���'�Fb�m������4z��ZY��5��L��e�ٺ�X���9Ů�?+��JB��oڴjt��ᙇ���5��/Xe_|��1EJ�HW��fχ������ 3T��k��I7ϯ��H�����j�]���vk��l��\�7��Ey$?O8�S}���Y�q��HfpQ�PD����V��PWŀD������'znj0��D���n��v�g ���:o@Ba�#<��Q����a�[Y�S`?܃��xJ7w�x�\U�W(�.���������9��s+Uu�fǃ�=L�S���_5�\����W�ĳ�(��}c�#�N!�s޿�j5Q8F�2���nwq}�H�]��x0��әu��pc;��gf2Bk��/�8�~�Y�%�nC%'x\W�'{w��˴��A�����%�Kr��7�kw���;�;+�����6�b'Å�>^�F܏0N+�׭B��V� �X̱	���V�jż�Zݸ�=���z5�Ap1
W�CJJ��-���2�� b����+8��������b/�T�sC����Y��B�>դM���0M�m}�QC1��	G�ZV�mH��w�|�w�6|��d�*�v� ��� ᕚ�Ɲ���*+�C� �Ȧr:v�\�S��'�M��B>Q�|�1�2�A~� (����a�R{�������!��81����6ad&�a��ϵ��,?Ɛ�\w�m.��K��]���t磟a{>xl}G�dȶ|�iq�dAm��9�J���p׳�ߨ�z�p�:Gl�0b~�o�aA��=Iz�&�|.e��m.���44�OהS���-a��o����H���L��j�&��^��/F���Z�Űpv&	�m�����Pw����x�Q��-�u-��PR�
p�<�F��qN�姿)UA��
�E ��f+Е�o�Z'����!�)�@ً4k�Y�����$[�}�Wט���LL�m��.e�Z"(OB�K	�_cx͝^P��ڿl6E�ȶ�ad�oe�x�Ӣ���&�����D��$\}�|��K�2�y]5"L񾑲�T�po�YB�*��_�"*�Ȟx�x�^6a��.�NZm&QS�.� �9����e)��J�R)}V�� ���[��<�tĖ���hC �ȭ��MY��*R�nb?N��0�*�
�mw};	�N���w�R=�@��b�N�}nIZڊ��1����}%/UL��:�S��i�����D������Oo-W��u��bD]?[��;����H�5@0�ѬJrU3�F����m<-4w�N�,w�e��A��PV�EC�h�WK�#��&Lu������������5��n~2^"��z��j�"Ihѝ�ɒF�Y$)�Z�sg�?w���d���r�FA�E5��)\��J�ێ�^�ʺ< �M�F��%�O���y����BJ@����}��F?H��,E��/)Vb���{\��ps@2���<�o���z�5��2QYYW%+%���(�\*O3�X��iҥ�$c(�J�5��rr���۟�[�yx>bv#1	|�����ɣX'�k�ؠmP����뮈��r׉����Kk
�S������[�Ե�&i�sd���,��tʩ��rI�
�\-�޻oXTi��v�4��!>�<�3L�(�Q�Sv�|"4۩Wb߲U�Q��J)p/N��aVBc��#B���
a]��R�yyҋ#ˣH�p�=�͔̜ʓ�b�vc�i+BsU��{�ڔ4{��fy�%�DXA�RZ��u�=�`��7 4�=�ڎ�$	\x��S��Y#����CiJ�A�"
��3��H������}��y��������&��c{�Ϛ(�0�U���A��:9�p�qFC�<'��KP(�ؘ{jѫa�nt�[�.����8��*�i0k�DPhX������+j��L<&���FA �Pk�rc��0V'�|����2K%
��ZG���f;�/����0��=��Vh@_V��7��x�}��	6bЕr�L��ڒ>�j1uW�똋�A6�MԻ�ɾ�Y��2�x�&��l���g�K	州X.���'Ij� ,� �
�}�I6HyI�ac�&�;�u��6�+�gZfϚ -N��1͢ޏ
sK�@����wW��.��[�.��%�轄FD�¶��X�3[�J�vO	<�w�:�F9xx:��&�b�l��K�{��?��=����������J�����' ��󳠷�=��R�#��r��7���)�bHnO�'��Tߞ�S#X���t��d��JtSZ���@v���S]�F�<?�\q��}ie � ��X�M�؛m�J�F�t��$ �Plw�~	�hՇ�oQ�`����@�Gŕ�h{^˧�xH����mH!Q�l�+U���0�(�����i��ĝ��s��a�y˄�?��"��(�R�G/H���?/W��`����D�������0@bΎ��6%?2�w4�^���R{Qo��9���Y�{��h��٩�8��J#��t�n�@u���φ*��)н�5�-�QO�!6=��C���z"ɦ������gwx1�c>�� !�?�QmP\f�f��jS�{"�j�y3ę;�9J��.܊���o�.�͘�Ł�F%�oW�Wb��H�G��0`��Q�=�Ο�º�V��q��J�3PL%�x{�\,:�����%�[<�!7��t��%�=���i�S�ܭL� ~���\�%s�{E�wM���`��MrcلL]�/˫������}���HQJ>�y"ǡ�40�տ,����T>������ ޮg��_9͹:��x��B�l�쉬�Pz���] ����j�;�M���h� ?.Gy�n�5���|��*@��#f�-p���=5M�<g&.^T�Q&|h3�����i-v�W� WNy�o���D����9��5㠰����w5͕Q2���流�t,Wz?=��6@޺�ި�&jTF���BQK5���~t^)�f��R�x�ۜ��Ē�H�&����J6Xy���U�ރ�`��1�c��1�yW��BcD�#�S� ǐn�Tr(ڏ£�X�S�0-��T*xe��H����_u�;G�y���������\A7L�hL��8�X�擃-�9K=�\�ܮ6�ßB7����.��+����✞\'��?"n�x�+�L/1 \>>4��4���/�����3
�/�K�:��F
 ^�6���a%i�C)�-@��ɼ�z����ps��?s)�0��yR:�1}�ݥ1�����Q����j����T���X� �����޳P�4�6�v{g�|bK�l6�@�_O(L�״_^N݂)k(%���s�#���