��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|ۧ[���B=PKx��{�Ƈ�����3��[��M�>���.�|"H?�E�9���iͯ�;�����UC�	g{���u��!|]���D����5�[d��0��N�n�;�C��2 �ϑ?z��`8	�a�c!E�����۵�.�R���3�X��'i�P����T�7�g#A�)���`ls`W���h�g�)�	֢ϛY@���9b�%L��/�4DPWJ�����>"��-�&�s��Fl�W���*�g���M��C�%��I��w͊!������t�����ЩKφ�ҹi�j�>�^*��<2�8��I������.S��Յ�*�Y�VVYϫ�5�A�Hpь�͊����ֱp�ɡL_���m	�V��o(�AVke�P���ɭY0chB���i��]
EDm�+�@��^���ݮ� JCiQ��Js���i�|����5�؜'���}T;>��4��  ��h{��M$!�Lp��e�;��E���s�k�025b��/���}�v����<,e>SɅeBN�a�����E���r�}W����G���idiMw�����x�0g�Ȟ�dL��~_�V+ә�-����
�@(ョ2������l�-�����ӈ��ޚ�Z�ð����P�>�TqMҲ�چ�m��c��kէ��,ע?n˂z5���!F.z8c�k�@7��܈�^G|K$?1&�:��{�8i��9���	}m=��e���]c�C!FX2<F�31>&l����LE8�x8�v^ȯ�Kt��q2p��%p��ym��l|�fӍ1Rt��Nߴ�S�ó������$E���'bʬ�B7��:cCJ�X��E�%�{\�V{���7��N�T�L��G�l^\a����9rɓ��g��18;Ko���"�{���@��\�pJ���}���55[k�<�M���WpQ�3s*nK[v��t|W�ehZ�w��#�d7��ҫ��X� @�I~ri�b��/}�ddx ǋ�>R���>.A�co�f(%����ڎ���`2p�.�3�|���Ag&��/ 4,��#�w�v��4>��x����Z7>(=��l�0?�t�Kp=I��r�<36C �M�J�ڸw Փ�kfX�]LK`аT�i�I���[a�����E�&�n)�M��t�ab"0�-�8��U��r`��P�|���r�PvFI�P��:�h[���'=���W踨�b�n*�b�40o���h(�6�5_�<�^2:��9��i�̹�/���C��Qg�@��؛I -��� _�u�C��ˮ�p��ζ�)�5g?@
� -X�S潺%3q�͹�t:�K�	�M}�zE5t7���D	��]����-Z��-�jA�� k�')d�q�}
<I^z���ֹgpP�B2��R�W��7�۲ܗ�C>W׷R7ר��޽!Z�g=�f���@hn4?+��bUgFG����1���I�I�M4�+b\M�bY�U�K���4b��/O���
�y69�p�or��5D��T��-hYB�$vr?�so �~G��W(��4��!a�g ~��X��+��ž�xE;r,��l��!U�]r�S&��Lc�sp�v�Y�w�����z�i�{ }���7V��Ч� �W�3L���V��hY����b��;���V����ǩDt!�2���荖�,�$9g���/s�y52д2"I�멧&�V��2�MW�pu��`����u����4���,��4�<���'A'�U[.B�̏��C3�` ���r���$���!�&ojb����7� mz/�v>CZ7'�����I}V�%B�B3eR�a�x�{a�=<��"s�qVF��Pd]��BCat��"Է�I�u���g��^�`��A����h�������2��U�6i]��[,s�/��ֶW��!��{�9ۭP�n,I|�d>u@��hKc_[<A�������Mhն(��@���X�0��/t(R=���z�/dg��]ȝ��+��;�-�@�b4��l	s|/\�%��l��T9{W�����7]��dF C?y�Y�;͈����	�����O�	�B{�SQ�Y����]��:�IV�;�1jLJreʁ�F/��M����zD�����#�ά�M��m����J��+�W�h�;YJ̵��"��K�)�>ל#�� �U=����s�m�gE����]���t<�E)jG-�N�Ks�9A��EJ`���F(�q��W������X{u��<l�i��JQ?�0�kcJ	Ni�jbRJ,�J������I&|k>zl����Üa�.ik�1Ȫ�6�Gq2-��ļ���5��Z�>��+|j��bP����ǅ�����˸�?�Nj�VFtXG�j�=�F'�G	�r?��,:,��M��G���P2���r�ާ�S���������p�+ź���c�T;�0�fQ��<A�X�iX�x�!��r	����|;P��i�59>��q&D_z)�pdl�n�m�Ә-��2?��LC(�	�~�Q�N���v7�������0	<�ZzęF�4�e���t��������@�F�w��$W:Ѳ�uU�ѓuP��)e��0�����سQ�)c�X=�Y:���	5I�A9����0M����8En7@|��|��v�6P�r���m#�m�Ȑ�^=�-ۨ/�f�oԬwh��oӥAPM8�Q��s�f��k�H�&"5I^�+���E��q��-�+��+��i*�.V'2���W�c3_��3Q�R��q��Lk���*74����y�s��R&����dGm�s]^P~�de�-�#ɹF���*�D�jA�y&���$������k����)�+�!Z5oϰ�kYD��vh���(�o�O<�_%���2���5;h�d��ܕ�7�����~^֌��;n��Ǣ���׶�ߺ�"b��.ji�Қ}��v��\�c�a,�_;����~�����lZ"�=�<T���$�9�*k`�T��������4;��_=Ӵ��G��.Q � m͈��+$]�⼔(���J՞��]��k/����j��sJ]��t7q�2M1�������sPd�ö	zRF�4m��[�&_�%�s;� �@�V�/�y�e&ld̵�`�r��N��G8���r���c�b�&�[���WA����u��c�C�f��J�ob���9�"�,��Q���!�^��%��WO��I��X@'b�pܥN�r��ᙣ��c#�Ty��2*uvQ�R��3�0��$L��m�x��;�RKQs�X������
����%j<�w=��������<��������ng%y���e^[h:*�BO��j���.wu՛��1�Cu����l�34K�����+O莂�o4ܵdTr�� �%�66���Sif*_�z��w�[�S v��¾јۤyh�;kf��L@4"�q�����/�҄�s?,������NQ��	����
�(FS%z�ě��e&�#`�!)!k�sKI˞��j�[�*���������߇�T�kQGbqQ%3��Ÿ2b��b|��vw��e&һ1̒��rx���C���-W����|�	�|�B�&�#"�y��YW��Σ�����zp��)x��^}!$j�+MA"]�g����3C��Թ��'$4ڌ%�X��B���B���֬u.[$�;�!��M�Q��ᅍ��QG�O���]��C���	@���`�}�A�L��P�8�|��]�O�hNN�P�������E��d������ë��.y��h�{�j��=�@T�S���3�2'x�]7	s[ȹi�⑀9E��cq���{.�߰C�2�N(�f0�s��mw�7�"�
�rv�.����g�ݫ�<2󼘉�Ύ<��V�ב�P<2I�˸MX/���ٴN�א�(f�U�w�#�K3�%o�4�9Wx/+��������nH�	=��h�ccD�x�����2� )A=/�M^�Ij(���E��Y�/�����Cy�LE����ȑ��p]����\:���@�<o����&O����=�*�u^�=h������N��(	�<��i�Y;zz��t$�|��b���A�5o�K�n^
�H��q�{�X��J�\ =�m:�$)}�BG����	R8�7���Ɓ���oK��<������?�=��y?)��E�&�ѝ���Z@����x��=�����K�Qt���1�,-�� ! 05�E�ǈ@�_��Q�tX���Xi������!�q(�G�پ�.�����v�X�zMy���l�e�HmŇZ�@0�*́�b�%l�G�8x��s��P�*�䬇Av;t٢��O��3����d4rL�.�$F�K �"�Q�sZ�9vG!]�GX��v�$^�ɝ'���s�:����zr���n�Tb��i�HzX�-#�d��߇�F\�&C�M�/a�w�=Cf�b�<�X�K� ��a�JA�}�����"���:�Z�4���+�[����4�ͪ:��P�p����ſ���2
����l r��ûs���o�"������G����q�:|�����ksł9�h���F�Du�衾l�/Ǩ��0��l	������:T�&�X�!g��j5W^e8�ѭU`�!�<�fg��K7��J�%�Յ'���`\����E����w�7$I���?0A	��sIֲ��U��\��8�®E�����WLl� ��} ,���J�{Vb�����x*T�m�}Dxen*FޝE��~�{�8<o9+�ɠ��/w�mD�k/=G+�V�v=Z����0t�JX���ӕ�W��������2v�Tڽ.�4�
�\��?��mG�>m�P,P�
�F��^G�(\g����=s!��0Ӏʇ/P�"��@O��G����'�:�:�OQ:�8�@>a�'�l���$�ð�<�E��d�/�,/�DcL-�1Z2)R�M,}~�r��	�Up3z������<��]M����H�Z����􎙕�O��Sg;K[��vA�l��Е�U����!yr�7J�>���lv�y�m��ML.��U��j:a�W��Z���Kh�r��&��ǈ϶h�e�^�����>��Fw��ڹE#�]�Z&���q��#�Uk��mڬ���\�(nI.P��2�L��C35�|��O�
QC����ݢ.4���l����S.Ɵ`I�Օjii� =#��N�H�%W�l�D@�hl�Qp����G�,�Cn��� ���ϥR ���(���Z�P����E`D�E�O�L��P��j"iQ��@?l�r�i�Us�%��u��mNGF�pޙbBr�ӯ�S�U���.|��ם��<H�b5N��[ޔ�q������^�jY��a�u<v���\�A�h>�[�@{�"���	��]�~J��Mж`�������#�Km�+Q�������(���z��)�" � /�����W�f������C�qp�V"f�`t�q;2�߿���㇤��m,����E~'�x�0���J������>�*F��ӦX￲��CF�_��b15?�7nV����~U2�@���ۃ����y�	�4@=u8%�j!5W��j���.[0`h�3+���3�TO� �@�u5N��˧�XK�J��}�uS��Q��Avp�b��HG�S�_�;�����D}���s��-�	ºê�H�i���l�&m�G�#�FA56��S�[��Z���w
���¿����ho��w8�*n<
v��*j�����Y���7a��*��nD���������b%�R/D���s��klQ����T�ct�D:&�	�h�������:���b�6	i��o���T)��$\oz���\�U�yܰ��/a��3��>{bfeD��#�4��c�C��ǄG+�X��*��9���e����n�mww{��le��E��������<��������\�ǃk�`E<��d=TNޖ����&ⵗ(P�� �@���5BJ���`]�k�1�`'j�]X7�3�n�۞ ��?��@����xh�ڴBS��]�1��0�K��֐}���)v�we�ӟ{a����;�c���c���V9���DiW�/�q������,�D�wp�2����{��,�{]��uw���7eS�㚯�]~s�-�bZBE�v�َ�?�����}!A+z��u=L�ci�p�M��/����(�6�k���a��*�SWj;�о�c�����{\�u���6��w�W�W�� ��d�ۻؿJ�A������7���-���C�'%���r#|S'��P���Z�"/���.��Q��H��M>޿�`�($���-::7R��SD�t�&\�����@r����*�7�i�&_�K�[�4;�-wQS�s����P��`�ZL��܊��nfJ�Ӿ01�ɋt��N��"|l��=n���|�*�IW���ՠ"�����ԍ���s��Y�nsȌ�A���=3Ю���q9�bV%�\�#0Y�V�C��pP!�@�]����7��r\���UTt������]��_��b����!~�&<3���ӎ�EVm��<g'B�r;^����K��2����	�f��j�Z�LȆV]� ��z�7QH2q��KȬ[�7���4�&C�̾i��g9~\�]LݓJ�;��);z _ò)�jkw��|4�씼h3\P���˜a�ԸȊv|U*�S�~��2�/P|�V�)��e��I����wsVcY�
[dM��T�mf-�U#�e:3D�6!��)O,�Ww;ZY����j#S���4�7��n�e�3��f��U�?��:j���;���\��E���z�.�f�#cVs����B��v�u8��-�	��Ʈ[z�4��M��.}���]k�RskogS�WEC��L�v�}��L�:%Vlus�ߗ���׷��Ȃ��GS7w�TS��0�&R*���6!3��(��y����6�h�J�6[҂�1F�a/�g�9��8�qLo�j�]���7<�`�|�qV%qE���~ZI/N&�P�-I����_����vIT�g�ɯ�A�k���>�2ը��a�S$2\���y�h\uY�AdRI=	Y����d�Kzl��.�u��j�r1t�6���$�ii��7+��w*�������JP?�s�ݴB�m������3�f�AR�ξ��y^�ʣ%�0�K���釜����tw+�W}�="x~&\+��?%��N�"�";���D�UOVO�P�p0���(.R��e�q�g3=�w�����`�l��րR����W��PE�X>گa?�o�z�2Ϡ�s�R\��M:]��5^J�����S`�.���{"���0�Z���eUnqc�$YX��zF#����w�%)m�'ڕ'�`FH�o����U�G0��7�3�����m������󔹀�Fh�T�
�gQ"a��<Q���c�p�PG���xT��t������-�AC)W1i����w�[��<@�;}~��}��$�L8����W���ӏ���qcP��N��X�s�$HPI�vb�9��NA
�bA(������Ls4�a���J����>�}� ٪׷#�]=����6�:����_�k&��8�?\�ƇKEn�}#�d٥�����3Sl��m�BV㊞2lHd�.p�|�η��_��V(�/&E�����l�ӆ�wU�l [k�#b�#�$����N b�÷n1��6g��J	\r�����:����J	h��Ȉ$��z݌9A�D�3>���u�'��E�n��Ҩ���;�b�
����5��D,6�L������1*E�@��n�y�A�p �$е.�0N�wBî�-��v���T�Jg9XΙ>&�r�0c�� i;e}Lu�`ɳ��I�z)� %�gozD�Ɂ�@T��<JMs�8��Ͽ��2�Sr#��ۦ��e�)aC����.�M�.p���}\����%rkR ���<��0���U�\'֙�����!Ǒ�*�lwDѹ� ���\��z�i/��e�Kj%��櫤���/�e��r^�Nv\�Y�z�%$kz��qi.��S�_6/8Rh��T���l���Æ��K�μn��kT�'��`�&M91��z$AD���b3���-�>j�.Wr]��`�`�I���ҹ+6-�zf��M��*u�וT7���85|}�&��G��L�����UN��
9�+'_��g����3O�&�b�l=
��K.,�<a7�;��>���X�^�,�j� 5r�P����'��զ���+x_�Axp?���*|&)�W�v�%z-���7%���Xx�7®�����-u�MT��Y��BZz�2j�|n�x3
%mn��Ӳq�h]!�<���:n\�����ɠ�G�2��W���R��Ci�.���ͪ���#O��[֎HuYU;S�Js�b�,�z���n�G�ص��gq?�v�N&�sHk��԰�KS�ޅ�ڳ���%�t��p;���T��g�Nܸ1��G�9�%�,v�F�:|/��۾����@��fq0����j��DtZ<j���@�\�L��$���:�T?h�3vY��eE�y0N}Y�n<��4Ej���	 �S�2����0U�g�k�*�gY�5��8Ӭ�Mڍ!0*��P�jN�M�8���Ƶ���)4<5C�ʰ�1��%�P��M\,ο�N�U�`T��O�Q��O0�V�gO�����6�Y�+C���ᇏU�#�L���U�e�pӶB�A1Pg�[�w�f�#eF�5�oXp�ρO�{_/���N*q��@���b!ڵ����ec;��T'�ҤC���{=���[�Yq#:���� ��Wo���ZS[O7 �m�[֚9��Ī���EZļ2�g�[)���f����mi��65_F�&�z0�k�tWSv�ljjCnn�*�H_y�~�âز�=_8����K|�FF�V��oN|HNj��A�%��P�G�5H��D3
���"\�7�$���P�xU-�7^b���[,��E� �S7��o���CS�N�:��浃*�b�G���!.�&mķ�^Eњތ���Hg3蝲5c�E%u6]��1���5w���o��A�&0J*]@�eʹ�kB��Y'1ⳝ|��H��5+;���f쌄�C��Z�v����6�6]��ȿP��ym�M���32��l�-����M��X�����N"C��i���n��ॶ���GF;D���l�%z�������앗�$����Dc�CB����X(Υ9������)I����P���Hׄ�T�&��flv5=�k�a_43+[�۝�[bAu|��B�VH�0U�q/�1��=5������uw070�" ��$��������[y�Ҫf�M�������7���f:i�vL\�6�u@��*B��X�飬%��{�z�<GJS_��/��rn���U�S<�5<}�X��a\DK� wpmP �:ev0m�Qd�4/rh��ݾ@��A����S�bԺ�E���S��*��3_u?g*���H UJL�"#��k��1�$����6H amE�P�A.{�I�'9SC-�)�=��2SX.��%����_O�]�Y��߼c�A�Xi�ڿ��J��M�<���#�Y��j��sT0kܞ�4�������:ؤ�0x)��Ĝ�ڹr�zXl� Tr�=�!�҈=��6+fg�])�K`$	*�R�\�1\y��3U�+<X�?��R�n���Z��|�ꄸ�(�\8�es����»���1G !lD��*#͚DS�֚��������=�l; =1����Է�}�Ќ��5���D�*�d�?���ጷ��2����N��S:��<t1��?I|Ҫ�,��\�e7=�*,�Ç�y�-������֝E����'�c�[+�(�y���n}���)g��V����l6W��&v����S�;�vʻM�F
���0��GS��,��
��C�_zg{�g����/���c���Fu�1Vi2���А����ҕo�"Ӕ<|��j��\9��[9�	(�͎čɱ迖�}��O����� %=]����Iz���[b����k�*�>�2;�um�ƴ��asR�����������������5���'N���5���y�&�ªf������\k>{Ts���tjc��9"[��&+|��'u���d��f
E�c{m@PO7Ī���;�@�
�jQګE��z�g�����J�~rH"�L� �b�0�g�9�*\z�V{�A�n=�k�u����O�*���
?{���=�� l�R[�~���M��/|n�A>㧇05J��u�I�^�R���'�n�HD�ߛk�PnF�_z�Ñ,�F� �CE�U��^1!'DKF4+�Z>��d�l��\%���N�M6e�Z�Z#�s�����0X�_��~^a,�ˎK·#OW�ʳ�K��Ft��Q�鞯,��fn������#�]��&1�{7� 8ܧ�+��H�4'�@&�cJ�78
�M�/k��a~����.}v-;��D{��E����R�<����3*����֜T��铟:��|c�����B@�X�4n(�j3@��:`�����"ӕ}���B��fļ�>�J���شy�9E�!m8D'��e��T^π i���dpB�_F���=����9�֛A�]�ta0A����,�a�fi�y�@�-�.#����]���
	�W��}Jv�}7��8a�K3K��F��FX�mG����Z�B��qRO�����2O���K�L�]à򷡊v��f�`v�	�K.����\��X�� �j�	�����}��$7�y�>
m�9$��ݧ�2b|�##���cSI��'!��n�jNA�t��cPr���Tt�	����?vS�ʣ���	�� ����
)Z1yV�B7-���mX0�'M�c3?�&TB{�[�ן�D�c�B��S����h���w���N@�(�t�}�ju�&�4f��A���a\,�CiU9|�ʤ��}��i��
z9 Ԛ�L�;���`B,���E�� =�"�z\8��9� ���]�j��BqՀ��B�����1-�w��Q��'���ٚ�$`N��X2�<�I�c�@��~�2�/�3�!Ӭ1�I��@>Q��$Q#&�}D���a�`!V#U�#�����+�c�Iz�/f+\��G�2-���<��i�>딐��@�Hƫ���QT�uX3@X.{
��Rߚ�G�z=��0��7�|��D���*c%2K�ِV/��C�;=F�_�xOz��h��o��9U��|0.��H�RL�%j��q���
��f�U�̈́�^ׯ� ���e�b��bc�@faCOX����ˑ�;��^���;������˄���\۠�k���LW�@	2E�t]���D��Y��bM�DA���Nx�a�j t,���R)lV�b����' 50�(�
�ꬃ����͵+���K���!0�GCq�;ϵmY���L��D�g�J��jھU����]`�⿀��lm}��q,�R:,x;VgI�PI�]���
��9tu�oV��0AQ?)|�Z}�F�_[;�TsG��4��n�J·��ُ[#{M3��臭?��qW��eO�[�8�$z1٦^�Q�/�F�wE��:���.I��&)����^ѷ�_t��(e �&���è騳�ٶƧ�BlW�ʊ���s��=ҕq)3tG�k@�߹꒟�Z���b)��#3P' ��>u���۹�1͒J�����A~~[IO4 ����as���y�;��}����������S��N�M�r"���YۡtN���&����x��뎅��3ɋ^�cXi�g��X�Ѭ�D�n>l5����������k2���U���%�p+��u��O��u>%��+[�vdo�|�q�{Q���]!�FP��Y�'�H���՛R=AK���vJ1lu��Vl�5�o�z[՝���"�	����EM|b��f�-=W�?^����f�l�`��:�� �}5>���Z��@Q��]�<�0���7�@h)�]��m:��b�f)OGI0��N���H.6R�0ʈ9�!��@F�ZL�#>��F#�gyK�7̬���/͈Q+��RUb��|�H�Y�D}c�_R�g���%���z�|�B8��5�3���&�`�E\�5<b<�G&�0��2}��ej1�&8��~�%8�4���@�G�G�W��Cir�����g����˔%2x���^�=i����#+g
�I�o���Mm{e-���,M�2V��^�;�D�[���É�k޾L0C�\����O���ix������ ����<��~L1��4rҺ�I�f,y��N����>y=�J��=Р�@��m��r��Y���X�]p�~�x�|Z9�9�U�������̻�>�65򿯭���M��'Ӊ����}���}r�t���	h.cn�&Ǘ�����n�]��Ǽ�t��bS��F�H��<�Cu�&�i�@��������P�޼|<I4�O�|��W�µFҋy"	;��pa���n��w�'&\ H�{H�)η�*�/[��#ϖ=9���V�Q���C!P�$�Һ����|c�$���ϧb�r�I�$��9�[��igս�j|�xh�T����)-f�=:҅1|���TV��$�;����ȶ�W��{�fU�\o�BgT���ݭ�*`�������L��41 s��z��,bx������c *���
#���17���- 
��(�oVf��潾9w6���wb�wB��6�3�sJ{�����ױ��j��_q�y��K��ZͿ�`Ub5�1��0�Nz?��qȧ��}x�a�����>�3����ʵ,��~��6�����9���6�/%R��'*u��Ze��`g.�jT4CJ�-Ǧ�5����������d���Q��H=1@̵'�����9b�6<�7�7}Y��𘿒h䦌kqH;43��֛���� 3��@1\�P`p����r�LQz\f�o.���8~��z
m�D���^�5�0cҫ.�=괐2���G�M��2Ȋ�����u���m�v0��S�3���VCn�Ryj�!茄�{��aܒ��Lk�8�nٵ�i��b�}W8y�:���;�/� y^q��vJA0e۪A�H�M��01$�#}٧�����l#���U�p�?'L�J���K�{I@���b#���s����<�iFܪ.�7���޶m$+qؚ��z�Hf{�� �Aq�cJ_U�#�k��&X�E<gG���`��T_?����v����d�S]�r(��}f�t�k���lT�N��ǿ֥ g[���k��ֳh���������C>�6j��9[vV�N�����0�۠vU���z�=�%$�<�vpõ�7�l���5���`�4�O�ƻ�~U�O��OX�"G��nOOz��:�V9�G�	>���Iی��8�`$���y*ߔ�Q ��=��_�X����u�SZ�6{�3�f�s1]X6��y�$�~<^$V�p|P��¡�}���G�+�3�R�C�,ݺ�}�ڨ�����o�7��!i1��>Z!���&�Q��Nӄ���"�!aǪ����##��k0i]��,��<���K�t8zW� [��P������AI��F�%���o!J�i���<wQ�nl��fQ�N�m38�M �gO��_u�ʍ�H�6�A��)'��u�W�⚹�g�H���C���{�^�-5�V9GZ�b����n�\=eݽ��ž��n�JwgЫ�8O�-N�&��S�dwD�o�4���cn�5��ZzE�`��\^�򢯈�C|j��LZuѽP�ο��C��F��3��G�9�R�dp]>��3��ӧ
��<�b��K	-�q��K���Zb�a������Ƽ�_F��W|��e���'6�A4��ގ��g�*�����$��.T+�m^���Ӳ��pv�0qDMQV��M����x]kزQ�(�T�^��rKְ���m�̏�"���=�f@��J����p�v����=����H� �nU�٣��3�3�D�|��V��d���x(� �r���8딂�ϰ���ʄ����NP���Oy� �9�稗=Un�?ME�
�'�Ґ Z��Oj�MR3�3�M�2���ߔ�f��2J`~,����ӕ����N�]�Q�ݐG֭}���ZC��v��M��}��A �c�����6 �M���Jhj�)⽁�W�>Sġ��C�u۠k��0�y�֒]d_���?�<I���cq���/9��e�A`�KQ�\L,0j��@֥��(R�(�Z��d�����u��mq���Cx/�Zf�����dZ������tkA��>���9f����\er2�%v�'��{++{�����5���M?x��_f8���1}�&���!n¨�(~8�v>%3��cI�Ž��� ��V��|%�O���nJk`��=�7�|����A*칎� h22��f��q���b���I�}����)�����<���	��5���JFh)�pj9V}<S��%l��6�&D��..�w6L�ݝ����q�S�Jn*c�{I�i�����5�@$I���@8��@���y\S���+gU���I�����m��y!.��w��h���)Ɵv���%?���͇�>1e��7�z'(1YOA�:ǉ|?騸#7���[U� p���u��ɧ��p���jG�ɵ�v�l�j��^��M�)��S��E�~@0�p�o��<� ��ҿ[�T�S�4̿	��҈�6r�<�ѳ\A�8g��=(��[�jx�a,N�^QIQ���K����5��Nfr5��u�E��w6y5����$E�>y�e�,�W�~��[9��	�@8���i�Q�9������A�^q(� �nx�B���U*�#���4)�2��$��2>����*E��־o]�ֈ�R��PӐ�y8I F�m<;Z"4ڂS���8���{���{|�E�����䑠�y������wed�_q�м�w�%���{f3�X�ߟ�݁5q�r�]<�X\�E�e�6M������+���.x���x/�E�s}N�K.�z'��Oѭ/�=]+��1%�S�v�.i��+|C,�^|?,���yB�$k`��c�9R��M39���W��<�T�����4�MwO0X���B��L����wɣ5�* D!�|E8)�r7�����(��	i������|Q��X^ �C6�|C�g����&���#U���hk%�.�����8�����7�N'�ӿ3��B��pȴ�n�������h���t�D����f�9�L�w��b��_�Ƌ[���S��"�fp-I���U%	*��B+��
� �2X��yS���,��ӻ��3�Da})f�~�fj�k#��5޿�E%��%��Ԃ�[[`(E2��(�B*��%�=>����!����4oUڶ����un��Ig�H�+F�����Ey��A�
1~4�&G&66�o�I��㪭Ir��)��W��4�&+��h�&�u�4ŗD_��oM���h��t
��zq����1
�u�Sbג`{a5�I�����r�y��˱�n&Ζ��=%�y~�d��&ꘝ����w�x%:�彊;�b껯KoH$������|���l[w����h�5Pv�6!iZ[�\Bn�m���7�?���xnc��=5c�ђ%{Ӽ?�����qj�L�� 3��j�
#S%u+�o�6��QN�ܥ �XM>Bd�)m{וu������8/�lNNV,�ۜ��&��L����PK������}���(�! -Þ����d�)���n�
&�v�dJ����NT�����Xb�<��ar|P��:`ֆa�/8֪g���/6;~�\��2��O�a~��y�^��Dj7a�6����XN���6�Wo�F��ю�J�e���c�߾2��LK$���Vg�+����4%�8|�p?iN�]�?ʃ�,��ҕ⍿�ӟ����>\���é�+���Q� V��t
��#�E�X"�C
�J���P����љ]㟽#U�˒�����y.ZX���a(�Ze�=�f����s(�Y�}zD�yi1a�#^�'����iod��ݱd7�.�.�5j�3�=_�~���ϟ�z4Ǆjۋ=q�N[�/��j�V?�!�#Lb�N���zB��3��K�g�d�U�l ���"�j)��	.�_�o%?e}�b3Z>Vs�����o���hurzaci�Ԝ������0&��8����lR�Ks�'��*�}~뱯���l�8��p�c����!�#^P&�0c�f�/�Тjr|9U}���,u�d���+z�kk�I6���y�zp��"ak0�H-p���q�.��n}�yu5gB��a4�����Q	Y)�V�6����"���n�c�z�A~�k�m|�"�T�Fv)�պܦ����<����6yiT���\����2��v��"��yM�t�Z±�w��5����ЮD������"��=�,�'�;�ɐ8�,�a�x�z���|)�v�ꏯ݋�Ͻ	��AeއN�~M�O��/������YAi�l�#0��-�ؼ��YD����!���O/z ��K3����K
 l���#�6K|��[��8�9/B�9��<j�gS�{&%�Z[^T�
�2�헰��ik�uf�eI�';��Xv�����CЂ��ռ���)-z��j���Uz�4��CzY?{&��9��J���,�`��F�|�ד�m�w�-�8Z�e��S�m�)����lnƄ�.�mI%���<�T����G���rw���H$C�ND_o��y 	I��2���D���[U;�3 �=�*��̓�xk�'�$/}ނZ��;�Lf_��I�B����p�ÒiZu����U1�*켐6�d�pg�.V�,�9(߰�U-֟�6�	ם�>c�c[-:'�k�[�D`f�߱�`�u�h�ي5����W�z,��a����jA(f[�.�T@�A�,��ζ���-�Cjl�!� ��ZrF:�Ѽ��n�?Ux�.㴗�A�e@vd��q2� &aƉ�B5־.[V�?�C���nYa���J�U/�-W��YT��Ky����I��jA�/1�p��<��Ѭ9͎����ʪ�0�m��@��R��1u��8��P�
�Lkg>����|��Az�.�;��J�����S��0��{:���/DRݳ�m�M�yF&�Ӫ���� M%JE����@Ңh�l� y;H�Y���$z��]6��-z��O��ޏٛIt.;�;d�M���m5�F����R�����4�2� 7.vs����OCM���f���ӳ����YRpS�	�����4�}�[�ofuԼU��>�4�q��YR9d�+�3'�4�/j?�#���2������n��G�ZT�!�}TK�Ӈ�1��w�et��':�=��}f\|�ʑ=��-i'4(�7��@���4I]�%�/ΏKHU���MGz��V�*���"����y~�L�5� ��Ue%_͹LU���X[�MT�����5C����Qgo҈��N��e���[;��� Q����i� �9?W���
�8j~!5��ʪ���	�z�`��#�AتTF�H`!]Ik��u/��B��C<�켼�n	���EݍFnV�����Y��ȋo�<I��^��pv,5���Y�?Uh��E�	[�1�>�{��?O�D=c����|,����K�(�ɖ���@og�`�`���qX$��&���8�V�E"�ʕuX�����0�/� ��NV�e��`r�`�.�w�I"멲�,�]v����9:T�����+�UO����B.�Q" !�\&�>�Ch�r��9�z������^d�ڃ��Q���r|�U$A��}�q��I�$5B����e�1?�M����%h�D
3 a<�� p��o����'|hn�sc���G�����V~
f��JO`�1`�y�І9�S�$�J�N������V��oʯ����	snya���~ʿ?}/� OPAXy�����HL����a�xc��v���/� �v�.)�ģ��A�A�wo�8��Th!c]��6/wŻDx�]���!=�쾶g�;�a=���U����묮�fr
�d���o�s�:Bo���B>�������k>.�ьX�<`e�OF��xg�e��o���e	��_����=��@��Ȇ�M.��yS���F�]��<p;��{�}N�rK��������N�~q*��'�JW�d��	z_�颁���9�b���@��&�`��^!N!l�h^=ݘ����1L�w��޲~�b{齅�_Aā'>�E�O��嚊!iF�JW��P��WPSc����*�z��^3�G���6\�O4��ȦGiSE.�	Af�į��ق4���3$f�����$q��ѧ/�].��;��0H-A`��G_�:�i`&�ۓ��E�jA������M����V��n��&��8��=FD������*����֜4P��R�^J0���prp�Rc]q���ਸF6l���+J�3>co&DiF���H��~��_�p�k@h��Гu\��/k&M�.�*�T*�O~w��):\�(e^j�}cs��+��P��)�-�쿃a��6��!��c��/�
�����
�!��f�E��
�U��}Y.IK�L�_�ѭ�g�'� �����_<���2���$#xP�
���S�����U�i�����U�0�W � ��X.B=���V��l�|Z=��֙�]ȨUG{��;������=EN���:�z۝�u���"���8��cz���J�z�e�7�D�y,#��>]M#5�U�
2#[¡R�ѯ�%:�>�y�G�:~g��)�Gy��'r>Wr�R�W��� _������G>���R�h�yߙӤ�~{��O���u��u�DA`� {Wħ5�=�LO-�{N�6p�uZ�dC=U�k,�5QT �:�������x�X�<l��E�){7����UE0�؋O��0�9<R4�;�ʏd!~ӹP'9U��Q��W�8��8�"")�����%���&0�,�R�.$H������ �� ��/�0|9���A%��T�j��� ��R+*N���[y"E�7��O�6��9�k'nӬ*̬�r���z��F��Q��.p�\n�;��d�7̶�i�WI�i�� �`�ͩ���YoDj������O-��c����F�qza��`�1B\z+;���WֲE��[�D��B����lA�H�`�o,��p�,�]���ѝ�.˾����\:�S7�	^��,��M:YY龆�UΫgޭ �/W�L���}Eޛ=%*1�z�n�G}{>*bd�t�)(���L�:Z��L ���Л�`e�[�T-�G/It#�*5J�2g������-ᶟ��i�2R���5��V��R�M��>&i��Eb2��1,��;�:f�K��J_����'>�� �}BQ�0&N��cw��~�p[�Lp'���-s3�PhXR�$�o�����;k�e��w�Cw���:�8�k��={f����&�XJ��B"�r�F�`+6p����Ѻ����"�x�{�'YJ���N� �j�7:f���ݯT�.�D����aG��Qy7ٴ#��s���b7*���u�Y�P�6L�Q9�*l%��	]갬�\�%wD[6��J�e��|���皂ԳBw�d�w�vj��p�
�Cz��FƸX����;��	x�s�B�ǀw��;��:����)A��K�]��@��E[U6$�HP ��{S퇳�R�NP�c̝��{�ǀz�O�t`��{��6\.�oa�
�kuQ�:��v%j�A����LO��2�r;	C��>��X��x�[7��W����r����eHղ|���ea�*�_�`r��撎 ��))q8�׵ղhZi���*�@�n��!�Fa��:�~��1�&Y�k���;٠w �\���M�9	h�0������|{A�����)�Fpe�=v[|�dR��`�Pڀb:[ld\uѽ���[�J)�d�w�����$�
d�w#2�z3!b���:���[}�0Nl�vR[����s%�Hz��Q�-$�'�b���=�^�������R�O�;ԥO�́6C�TH�Ψ4b+^��zό!���I(.B���G4i�g8�m���QZ�CJâ�3n��2��v��! �$2�hۤK�̾�H1QFv����f��Z�
�:�^��<oQ-���v�R����x�%���GJ�sR	t*4w�h^�Y������F�sJ��ā�����~ޅ�<"���奴����Q��m�j�-Ǻq�Orhj���obȊ�I2o����%�,����Z��"�c7�ќʒc����X��<�[Hr�z�ß�f?��}�qU�IRZad�m"I�!��ze�1	�����9D@�ˈWu���ǚ������F�Z���B�u���潞�m�������+��J(Z���znb�� /���,B��p�O�������C�H��$����f��BR>�[�D	.4��]�"��.d���Z��:��� ��!R�M�k��x��8!l)s�!=#��d��-2o[�����$A�d�0�+���WR�	j�.�{�)�Z�=Z(7"�܉�[#b�夜�fd!��k��I��������X7�c��6O���9bH�B;k�խ>�<��~�����bz�9u� s���E0�m9[��jA�#K��v������2�T-[�rЈ8�աp�Y�&L�$��鸚D�7��U �^F�U��;^��4q߇A��8~B�&��?��N�$_e��m���1��¬IB���z��q��׍&��h�:r�.��|�`��
�C�G��4���t�O+_4�Nҥ_ń���dɓ}��9?v�j��)Ν1��7�W+���0~���}W�=@�3xVF��E�4�'��Fk���FZ���[���3��8ߊ ��TTl����m��fJe�ᙍ�pF�5��d^�ϲ/��y��lhw�L�}P� �Y]��ҝ�2֧�6��R0�ѩ$��G�ٓ����P]�)���#�0�트G�c��ɭ.�ؘo����29m@��,�0����#U����b}ir��ho�Rh��^^:@��BΥ�����<t��Ml �b�}O�ԭ~�g�2��[i��u��m�n��]c�C�,��Y�^4q��
�v��5~TG*b�M��D����l�'��cx�>���vH}j���B�N|&�1k�lEl��<�����:��MiEE1�<=�ˀƟb~�q��L��l<�P��:��O��*�g�K��3ix�e\�~�t�zf�ۍo�E�23��h��n�a�.��3 N��B�t��!�KI.(q��i���W`��"��mn���[@���"]Ke��Vn)��#i+������}��NXCP��@�u�f��VUav��&�m1FK���_<�9������Lp~' ��*J�{p�AhX13�	��G�}���"����>�×����#QK�o�����)a��D�����(�@вƮg6�9� �̱`S�w .E�Z]���*^�s8z����N�w�b�Ak�|�=hMr=9	��d�t0a_,��>�{�>���.�s�Π���rp76 ��U�qj�or���G����| ��C�D���4b
_��͉��e��9ė������ ��Ka�yzDE._��5�b��U�*��#o/�y�j���	�6�s��+���S�=��i� �W�Rv�>����h��f�D�@U �i��rpZ��cfNP��x�h�L`o�����P[9�OY�tI��8���-}�'D/�Ep�V<6�C���$�M��X"\�X+��r�T ��W��k�_�r {��c0O#��Ǡ��JU�-Bo�v�a���{���C��K� q�;��c��U��\�(�Ԇ�0��� #��?j:���G�P���ӿd��B&[OE.ZX�����,rs=a@�E%,W(��� ?�P髇U� sL���ݪ����C�M�$��̀���&d�-�"r�W���y��>U�7[8�����YƼ�Av=$\�G��!j�etjK�aMA^M�Ŧ�Ӂ�6�.�8�p~q�Ђ���1L݁��%Ю�*poj�
I���á��-L��5�VE>��һ�ݾ�[~��B�?|)�E��1�vc�pD���8��d��L��o�fr=)`���@�B�m�h�</�I�O����3�y��I�1���r�����}^�~���z���k��%��ҵ����{5,�� ٫XF's�����ua��%x��a�0�ѿ�5������vr�9�C�{b����DDFq��u/�w��ӻ#�w�а*�E�K��1�_����P{x�Y���4rP��!�eqF$�#�Z�n��m��%MY� d�\L���)@PU^"��[�H}h�jF���B���U1�_�%�!ηt	
�W\���Wͦ� �'"T�EZr�î�U	�;���^*=�fe����H������@�`r��J�ǃ���R�MH;��L�۪PcͩŢ�xި�D1Q��o��!�,d�u�n���xgD�w�r�H��ڏTJ o�W�^i�^�HD~����_75�=���{P�(��N1>/�z����3#��0�wz��gkJ(�%�8����̲ܲ���m;�N�o���X-l�
��\f����v}��,����(L �B�&4q�ʗ����Э�%��l��hA#./�|�����1n(b��&$^؊D8����^@�jbJk�vD6�&���Gj�9X���AH`:�̏��Hqo���&4h��e�����3��{.�8^���-���㔸�?���A��pa�� ����3���Ӵ���1uRu~�c���H�Kk@��`)G5Ŕ?�I(%��6 `L�	�ރ���M)�/��9l�H�s�����F�D�-��R�=s�vb`����$W��Y��Š�P�7%�%�%62S�z6��	�x=0���^ ����:�=��W��!b}`��5:���*]�`�+�����10,����-��CTmj� [�dcorQ��]F�$�^�W'/ 7q?k�>j�I\��#��kX����JP����v|�)�UJN�6�����ܜΣ���"�e�T�X��{lR�ʶ��e��/vX�ޗx��ż�8
gu9X2I�j���/,���z��>�u*�WT�v�I������r�#8�S��E����V2T�L�FĨ�p5��m}�Y."��}�V�ҿ�t9:�g�x��C��7)ɍ[7�tA�c+z.���!ax��l�ͫ��͜	�����cCv��v�5(,�A�(���j�����⤀�#����r���N^ ��k�РM<�H$���e����+J��2�ʻ@��Y��,��� jt=&I_� g�.�&�EN��ݗ�X��KO�:D9��ӴjQ��w	�.{a8䃭�R-'6
>�l�v�Z��Z�L4I��1n%�	J�aF"��_J�����~^�j���V����A��*U��wd�C#�N|7�.k�,�XO��M�R��{���mԗ��m]����[�)f�����*
��щ��NCw���� ���T��GB�rq������~&�M:�x�WS�(�J|~
�:���-�Ib����H@��w��w��{�j������t�\4<����P�4��1��ͫ�R�i�s���� J2K��I�/�l-I�-}�2�tG�wBX� ��ͤ\�-F�'��%`�K!�_��B�j8աƇT��Ԩ�	�{��1P�X��+�T��'��Xs/���%^-Ӧ6�`�~���
-��*PEޚ8���ȣ�Q��>S��d����Qؽu�[ �|O�#�J��=[R $|N�EJ<��~�Uy��o����v�F�g����ƍ˴���I��5�큡��WS����Rg��m^H�����k�^�=UlU?O)
��r!:vhe8'�䮩�d�	�Q���F�zN�������_��`|��
���f���(����x6@����=%��!���4�gg55`�[2|�u������9���7�[ 80$u�9eÀ������@�!�ۇ�8���k"�>�#���>����[���4�����XÊ��JA '.�9g��gj�
�}��;ʨ*C����BW��$�w���u�Rk�'�o���A�ʄl%�+��ʍ��׋��c�RZ��Lc3*u�7��q1xB��hڞN�8���JG�s���b_[���p!wB�o���}� ��`
�V�����(
�h���Q�%�[ӓ_��{�b����G��i�A��<�Fp���xK�Oұ��x:���Ί��@�|u�`�"&��`W�+�&��l�h��i3�y�5��g�>w�E)o/��e��H�&�;�Q#�c��fʂX��Q^��L�&Fs��@+"�?�dv�����֕�uu|tO��a�2�ΘUC��*�?��G}l�5�0��U�@��i\ߍ���-�%���~���"�G���ۯVD5�y�}����|��bBUf�Tu����~2�`����/������0,J��H��w��0ۉ]��Oo�=W��o��#�v�rZoH2D7�&||"_W{�I��	O��Ou���1��HćA3���}5�E��l!��/��Ì��bW�{��-��-?����Bё��i�o�	"��_@9��JI�Eø�Z��j}��(y�.�ru�����"љ;YD-��d��`��K6R���kCY6ă{��n��cQ�#��M'�+��G���7�K]y9s�y��ƿȍf�Z��-�1o��_z����Q��T/ծ�戥;}������$n��@���F�P�p\�/G��$�9�b�lfƑ���v%��-�H[^���xq'd؄�l�*,ë}���(5Ғ�J<eD�ֿ�,�4��hB��ږ�F��MJ�|���9�~=c?_�6��E��������`M���`��m���s,(��[�Kk���^I�&��*»��ؽ�H��0��s��d��꫹}�S��q^K��S�D��n�&��fsqt0#��s��XB�'�S���=��y{�W	�t��_@����R8:j67?fl���^5Pn"�G"SL+ޞ�B\��L��l��R�ϱ�h���`	* �%�^�o���@�?���d�xj,CǬP��2d|�I2]i�������nU�:�U�9�H
��v���5�<�X��)6�B��*av14��"nW���f��Ҵ��kLp ��,�|�}��{�ێ�@%���g�v�KS`r��v���i"����ؤ<�H��Z��'H���>����
/�Ӛ�y�y��Y���Fغ! X��YnZ-�	=c�FX���)�**'VIb�u�0�P���̈Z��`j ��k�m�����~W�987��m�c�O	v�M���߻�'ԋD���\�BK�,<���<�z�ow���ls4�\�9d�x��CfΫ�'#�k��r�Z��FY�&������8��)�!�j�Q���������-����0�֘���״�w�ϡ������+��Te+A)�k��u���4O
�?��G/��(O�B�����>� fQ��FQx�=�<�R�$������m�A�k�d�s����MN[������:P�9=[\��_�|Q�+�eY��
]�]�v��z�CYA�z!rLp�J���ot:̜��\:���VU�0S����)���q���,���r���?������%���[���/q5.�Ғ�/��� �Ǹ�v�i>��e���g� �G��EX=�Ie T(�������
b�=��N \����f�e�XU�0s�Or#|����s=��2o�؊J�	%Ɋ�V�4��|q���m�Q��d*ߠ�9~5�4g�u�E�"֗UYܰ�=*�yǽhu�w�Rv�3�Ȗ��+�w��A3Z���ܵ3��d�T5���	�v]T5�lӛN�)@y}h(��ݸ!#��`c߈'ùY>q���ߵ՘ؾ���h�;����g_]���?�&�%��������9���� 
�~�.r=���'<8���+|ea��"q�M�7	b����ǦOL�߄[\2k�>ꕪ���Z|�*����Vn��j�)y���c"���( �t���ɭ�"3���+��f+���@;DT�Qj�@)8�͚�̀�o臆,����F%�Ăx��7�p1��}�9�θ�O��ҩ�t)��ʵ��PQ�BtO��M��e�o�{zb���.R)`�"�tr�ݿ�B�L�v� �sX����2\RN��YZG:-�����$�,����k�o���=��i��|����j3�X�kEM;�g�dKz4��i gn~�]���RdY_�����L�q���z�5�-V��U+p�jf@l`�X/6.i#X`ME��-|����C�DI��G:3��T��]�����jT�{ë�i���ц5��BA���"�ݜ_��`kmj4+(b�z��X���vT\�;!ja�C/�@�p���#�����q�kaW_wq��*����I�HVݓ�w�`UP��M��oUKP�h���~оY�f�W�~$}Ml����k;·��%� 4ށ�
+���D�?���>�_�Yl9*_Nŗ#:��ZBx��&����k+�R�L������ݥ]k.a�niŻ��aS�候N�'+5�-�{�­\��E�I�T.m ������P|��|�Qu�VX����tD�Q���l�|�k6��8{(%m����+��?���Nt�^.�{먞Q�9ND�Tz��.سC�+�P�է�U+��5D��#��ɘ�rXp�Pf-KLڬ���v A ��7.UWK�����'U�%bV9�[����F�h��`�P�u����%l�ރ,aJ�x̨��)�7��,Ұ�>k^
y�c/|�C�/<H�6����)�$�8OP<�i"uA!j!�x��j�r��
6�z�Q��o>Q��x�:���N�C�= ���)��vC���o��A�I�s8��v"ȡ�u�ͼ�9!N;�k0��)��i}�xƽ���Z<96�Fy������g{�l���D��z��J=b�g�%�5�K"l��ލ��9�K�s�+�a��d�b!�9Y�����`@���Y�9�x�c�>E��?]H�!ٽQ� ��nVv�ma�z7�g0��v�mL�G�,�MlP��`DC����JnTR�b��N�S�z4�!�	�,��+�k�I�-�ێ��1�V���MX��dQ�겆N�GO��x��-�RɈz���>��|�!�����Ge�c�V��#��Q_g
Ş�rB'�)2:����d��X���o�m�ϡ'@���XCe.�D�nPŘ����:n3��������V^>���i,��ݝF"�Z��-��(�J�����G���[��) o�XO���ϒi$m��Oe/�O
��I,��V�h�|��طt�j��b�� r퐿̗�a���=�\�E�)��P�X��Y�fY_�Re�Y%�C�*T�,&V��K^Q�a��W�5��8�-�3�0�I�:�Q����G��4���?�vY�+�.�����8\���7��QA�Yցѧ�0��Zrؼ�t�:�(b$�W��B�__i�^f�OI�o��<3���b�\a�B^X��#vꔖ��Z{�n)�}@����} �E��a�����G_���)��ǡN�c��U��[Z����$�9t>�>�`�kuڵI�+� �va�w���2���%�z?(u25T���]�9m6`�JfM�.ta�N��[�	�J$\��y+�8#0���o�A�z6�E#��iO F��^`8F�o���P5۹���O�h=u%@c~Np���Z��4$���/����;{�\��j�����+A�W�Q���}0�pe��) 5��o�������R`�^Cnh�,3�N�hć{���w:J��۫c��<*|�m�P��~'w�@s6���ު x^�JB�wk2�r�	_�����)�tXQ�=^���!^����nk�E�҆U��Q�?M��pa�]u-�b�`�Y�̕(���y�/M�������{�s9u�j�i���l@����E��֘�V�X�I�8E��;�#��1�v%�釘O�S�(xE�f�C�N2/G��,��2��=������>�,ƴ*��2L9�i�[%a��B��<�GEO���3=��Wa;���f�G�o�Zm��_P�:T!0�f�,�O�Ɯoj���U�I�S���V��4�6@� e��B����Q@Qs�'6FC�V�Ik�d
�z�p���˅�ᗾD��'��^3k���iWϤŉ�M^ϩ���!�/���!����0������6�}�a���V�V~�l�o_s�A^F$萀X0S�N�x��t�Nu�`�#4��i$��=CǟP��� �M�/\�x�W�;��510p �����:١4���~��I�.�2\MK�?h��5�`��{����|��<�C�d&�³�۫����i���B@)!|b-���Z�դ:Jbtvi��1�ޠ�o��7�M�eǾ�x�ybC�D�Ż�q�F(WJVAl��8��4��Y|�PE�8Q� =����5Eේ7���u:W����/c����W������q-���f���3����q���G��������o�����51!3~��:���lL����1��E��ET�atQ6�6�� ���s1#O<o��54!�!��At=I�(��T�
4{4�#+3x�gh�p�~ ƺ!���j� �8��SL��L���&xг�^�3aӼ���d�Xȼ�$"�.}& �-��껜8ﻟХB�ID�;�s5-��5�M?Q(�� b{�Q櫔f�ARr*�E�r��b�����h:3�&���;�ii��<��ɨ��b������"��pM8D_��I���J��+#}h�q�*o?t�6E�ZȎ+���I�*��I"w�o����m����[��gb=	��� .�"� �	�a��Xߴ�!�GDy�nL��Ħ/��]��!�Q��	@<�����W��lگq��V״�U$l9v=:�O{�X�>F����e�X�y�K�W	<D3�,�e�Wb܁�B�;���F�Ч*3��b>�GC�N�m����S��_�O�~�E�<z�Ϙ6��3p5ʹ���S�*�G�\�*0�+�Ę67I���j[h��3�hNG��l:S��e&���7��0Ɔ�h�@B��W'Ҟ�7b3��φ�I��M����%P�ײ�������!:��,$u���0EB&�G �@����k���'ѷ����?��A%��f&Fk�BeG<�jO	�YwS��s��m�K�Fs"��\���uz%�4!��(:7o*FAQj�J�kd�����d:[k��Z���K��+��_Dg9�6���8�ʢ3��zzsLw ��}_�U/���x�k�Ȥa�eu��́bcMj��KZ�vWv���A �[W�r��#)W�/nWХ+�ax�U�\Yʒ�#�/oF�C �2�D�*���Y���s�1^�U+K���G,����/�n���a�.��'����Gh�|�(��4IZ���6�k���O���Nƥ�ڳcH9���{�]B�bx��.x��w&nBx���|k��U�w��X��u��;���1�Z:)A�� �{���;T����K{2�]��3��L���O���C���i-�Q�X��,J���6@�HoLm_p��/��$>��1ʌ�>�c�ݛt9^�3�|X,�^<�W,��&�� NK�;78��;���OIo�ܯ�8�X�cv�:oA۽8Ƙ%v�F̧�XPb��_�䪉��{R�Ŭ�R��y��V����f�m��ł|���{��g�t�C�|��@<�j��8�Sh��2/`��	�/�����>_w�?���@`ѱ�gXY�H���u�7���r�f�y��30�.NT�{��)��q[��)���J�S�ǓE�o����� �hR�+6���]��y�Ŕ�QR�Ʊ�*�TYŤ�P^lht(n��v�lu�uQ�2���3u����|��Þ��"c�w�yj�d<�Юû�a��X�$�R)�ڠك�Y얍��r���_�2r��4�'�#��[���� 5�Wvh6��P�W$X�}wa/�-���1�
��u��}��r�1�x3�
�e�;��ΥvD|O�Lr�K��9u���c�s�=�ݹW�qk�v3o��vľ7��Ƣ}&%���;p~�RI��䙖OTX\C�,���� �L9-�`��M:y�Z��^�]Zږ��H7�q^SGQ�j���A�D�  ��\0��LC�궷Ǫ�)>/N�;3�S7����O`,���=C{qKS�V �|���_����������dk�����Ђ�a?x�i1��Đ%�Py0�1���#!ޅ���h�6�z�������z6��$�}|���+Ł6���j��1r���[";�&2�3���x�8f�Q��;Q�Sq A�1�8	��RvNo]@�A���L�%$���:�\�����""�����ȿa�����WԒ�d2��A�x�ޜL�6��y�i�'!i��KW|(���}�?���q����LPEͫLw>�"��A�h�M�[�&���?y36�ӗ����Ǐ�M���~�)w�Z��� DM�r�$�8��;����	o��K������I�g�2A:'�Dձ�8q�� ���.8/���=�U�B#�`��ؾ�B�s$�A4H;N�����n�}mh�����^I��ұT�~�f�2
Jm��a�Z̤t���i�%|ʓ;B�����W�{�[�KA%x�(��{�a��l�PX�5�rO��g�pu��锱!N�F���t�F��MO }b�~�XJ���*۠�}O5e���r������(d�������s�U�@E!5�R�4˞'��(!^c�Գ&�/�0YQ:5��댟���Ļ����?��'	l�L��7kdԁ��ccCNT=6]�j�J��I6P�L&++G�U��^s�i��ơR��7�t�v����p���ՠi �vi��F	4���2�Ff2@����z������/�אM9;�yy�E,��BN��/�8J�P�����VXU�QT�hSz�h��9�����D�_yF���:�<#Dv:�-e͇?��Z�|�\18��~�4�[9�� �c�J�o�b2�������H�V\��u�(+;��*Rn6���g
7sm��s�!���	�-"�5��!��0�Ie��!�Z���)p�ZTY�ř2��7(Iʠ^�w$�4�Cx
���3��5i6wƪ��j`b��d79Є�	: @��q����V���\g��ڶ�$�bG��2J�$ّ-��BY#�nJ�w ��\�?�`�6�K�R�^^�B	m�QJ�e���t�'US�u
����gj6|Ũ>�w:�/n�-e�n�R��!�;;�?���mf�Rgk���c�ʬmG\	DV*m�3q����S���b%\�z��Ѫ�w��M�UE��rW��%:�ۯRN<z�M�$��;Qf�Iu����S��A�A/uq�$VV�� �q`ދ6;�N؍z
�i��s��ϩ�E�~�'��40^�0�ƅ��c�`����n���a*%uo?��b
����B����d�M�w�Y�����}�'4�6���CZ*Ў�g��w�ƬgE��2�^���%�pL��(��]��lO�07XNA�'`��}=ԀS��Ì+�{��j��Vj����R3�#%[5P���4��޶�}Uhyu�uq�N٘G�Eȋ�{o��e��\�M#g�C.Ȉ{�,�[!g�p#
Hk��ֵ�*m
�0����v-��ϡ�����0��S�����$�����@�;5ꝷ�c>�Ϋ�	WaL唡�H���(�PZ�u�"�l�}c�0j��|[�⭔���i#�����"�����V���V����Ж�G��Q���5�Zs� 
g(q�'d���rj�ʶݗ(�_� @f>�`*7�� I���o��׍�����GG�&�^T�7Ne��=���>"� q�O����~cI�HL�Xo���% d�#Ҳ�m 0�k��v�q���R1��P�4f0x��.����SQ�I)0���(�6k�݊�,���-�s��6&��Ѧ�J�~�C���:�F
`�����Q�4�-���nxZ�ޢ�N �@��v%��[����h��Ix�;P��.��0.0�w������sc���gMEG�M&�A�QӅ��gY�gƗ���9�\��g��8J�,%�k��;�er+q�X����F�
kƱ�lr#	��O�؎�g�����@�a?���R2�i�ȳ�G1)c��J{l�����5,y��{`CF7�6GL���6��C��]Ť��i�5韛�P���d��6��!���;� �m�̱8g{9އ���`�Nȣ�2��[���}�-ˊ��T.v�q3�1�.[ ^<��6  �N�/��&��i�pș�u���Z�K�Y��	�5��@"�m�+�)�e���Q�j'��W�6�N��hu\Qy��r.��͍<"^����������Q̬w�l�|��@�p�{�ѻ��j���V���4Ӏ��)���ָk6)�R�k�@k��ޤ���դ'C�Y�cE�P3̔r�M�����Su��6�A8!Hu�^e�l?�\bC��ʼ�<���i�镽��i�����P�l�' (^^�k"�OY0Ln�/=N�{�~��j�BU_�"��dAX��9h��m5��ɝ�+/t�i���c�c�B�ê4sQ'�V	=QD.�&��/�dtA2ׁ��n ���y��9��į�,��>�D���1;z�uZ|��nko��呹��U5Z�{)^+�$2��dA�)�f�Ą����v:/u�����#W����nYuhv25W��ײ�c&����}���-S��QI_lT	���*r���#ȉ`��]lI�?^�=D�cV�U�avy�ڒ��=�oRiy0��C;X'GC1<��,g�Q��m7X�/�Dh����1�<Sn�H�[�Xu��yw`�����n��6�� Q�b�Ys��a��,c]f��g|�ܩ�+h���,�-}-� �o4w� <�5���|4fW�r=���U�Ύ���Y���O����Q��1�db����ft�A� ���$l���j�[��N�{g�5f:) @\#��9�=]�(�V&��u|a! �AW���}�����&L��f;I�r��!��n��C&?�J>
�Ip�Nj�"3@޽<��^�g�����9�H�9heg��G|'�.U�[Q�d:���Ӥz�O>Z�Rɕ������9�Q�칮�</�������"X�jeh�:�+=L�>=��Y���\6S�WWV4�����fP�Dxx=����<�w��rQ*�\֠!�~ D=�?����;����e,���ެ��t��P�N�<i���gGֿ�<u��mi�έZFHI$m�����|��㻛 ��R&0G��9����߻���J4� ���no�yb��n4ߩ���@�3R,�4��gw��ģ˥�A�Es�h1	۴�haH4o�0�1�Jˆㆺ;�5\�#��J�sy)D�IF*H{���>�?�#�m�Jr�'������T`�-�;@;|rЍ.�P��=�'��-V�5f̪v��Ǟ��Jz���'#B��Y�>ش����É�h/
�vZM���q�.x���
�N'&NZ!��+U���)��X����e֬z7��I�!�ȱ�<[�gc��r�{f�������u���V���#{���g3�B:w�ݧ��6w-^1�jg�W�[��64���M��������{�ޑ;b�eEh��'v�f���U��U�^M��1�J�a��X������?�F41�Z,��|U:`�w���ӵx�����5q�Ҡm���À��j�+ƨ���_B^re�(�9^
�����nL1�]���N��s��%�8
���)�?P�d� &3! �~���|"}��#��ԛ��D$�XSJ�Թ�$�i��!�;�x�F��z�\�@9�MF���L�;�-�jx�y���I{�whG?�-�5�e��կ"��M��-x����t7J�J�P�_U�j��j�,����
t��:	a�|Ih(ƞ3hY������xhK���Y㜅�A��%W4~zFN�`QH�� ��D�T���b	�e+�6w��w�o�� JNz�9Eڰ㨆�����V�;Q䆁��&��H.�=���m9�{�#Tq�$��H�Z�zM��6K�Y�^��@/�������<ydm�& �����o�3;���ĥ$�6ĤT>v�EL�2!C){���p��('�=�-֙@)4ȵ���	��\���*X�,��9`#���&�oe�Ak]a\ My�|JRu�6�ˎ���7%TƆ4�l�zn^b՝>TT�WW!��{�}邁�BgI��僖����9(��t��\k�x�
)n�uJ��H��rd��b���~ ����n�������k��3�[2?Q�"��F�1P?���+_L�U�ֳ��G�����*\��_h�r'��xO�e���Ing�`�Q]��W��b���w�*U��e��L�����{O�C����?���w��EZ�4��N�3�ŕv qr�<ґhJW晤�[���䄴�������<ftH�i��	Wa�0L$��=�E���,��m�@y�ٝ��:��a�a['��)y��l�Gec�%� c�֬9m]� �ˋӪ/ש'��h�]g��~>���0�9"�`���{CS����
1Ñ�&�S˽6��X�S	�'
z��A8��؝k����ps��~��6��c��m�0:�I�u�!
I]�>eb ����Q
��4�AK�d۝�o}
��6�C��� �����W-�Z	���˚�S�t���f�w!4�u����wA�;�ą��x�auz��>�DT2�ߩ��@w��A�3�l�%̒�4�3�|<�n?�[@��1ԱI�������9�&3�ؗԇ[1�U�M �Aj����Y��;���Lk%)�'-��:�	�@�O���ܸ�FP�D.8ۊ��:��>Z��4'�5ѹpZ��`��[F M�ȓ<gA�0��B�:AEM�e3�Ȝ �h��~-�C������w���ϩi�����,!mTWĲ#;0��U;�\��`͙�})��剥y��Q��c��98��#�m.<_��u�@�����ç#��9h{��
���&}%6ִ��Ƒ�d �(qai	MU��~�(y>��\_
����(� 6>��yZ̃�X�i=c�fQ��~Z	��]�9m;o%^��;dԏ�P����J��דp��F�y�:���Æ�L!���3�_ ����N��o�6�V��BhqM|L�\^��53��Qv�y�c�K�p�߉��$"5�E�'�A��ϛKi��-�a�k�k�Mq"\ŝg�fDj���B��x88��=�����	n���uk����-��G���	*�[�0�����gJ����by} �/�~��,�N�+�]/�Q�zT�d*x�~���G�B�'/��gUJ�k�pSo��w�D��8�f�FF��3w��O	���ˮ_��8 �)�e�w_�V��������d�SOF�&��!��H\N'�����eL2�G�O�g=X§�/��i+��{#�v�P�c���,�A��s�r����H�BB+;�k>;/�X>��=H"��~�����^Y�?��}�J�{w5��E��n������];��!����%���]4.h0�-7��j�,���I|�x��	!���������n����(��}� N*�F`���7�1��� A�nɬ�ᇲ�cG�����09��@L�S3��D}x�Q��Nt��Sf*��@x��5��B��]s�^�5T�Rd�r:�<���&67'Y� *��d2��4:Ok�~�M�yBE����Id��9D���ܗ�;�'͒wB�nO��Zv]V*��=J�`�7�t�9��T��5\'�iN����#��Ի-�2�G��m}�	D��Ԉ����)�&P�F^���@�VE��g�Я��@�(7��} ��`�t	,�!�(�I����(���Oz��Rc~W��t��oaj�gՠ�\b�����Rc�j��`�B6�����x��^Ƃ�6�-�Wwy�Pvg(p���O����G�	����4�XW���8��b=4̏�3�����A\���(��DH��,0��b�赗#���@<���ܳ��d�Wܿy5�z+����+pM�
���	��!�|B�F�p��E�EK3ဆQ�cΔ�g��tI.��� ���2A}���,q5��{�$p:u`�M���N2y��às�p�<���?��g�8kyH]8�`:Ӫ)�����V�9����=Z5$���O5[����5(�j�Z���t����HF�t�P���Y�$�Y.�jgܫ�
�8�I�(����Y!��	J����T;纛y8����t����TF��E'P�5i5�DQ+ҟŽT�S�Oau�؋B��a�M�����f/o�a����SJ��|�SX��W�,���5y��7j��P�s� B��$ �c��C�����f�4��mCY29.x�'�i���C#����H���C/��krC��޴�N��������?:j�tZ�qQf�i�U�R���0VG���?�9=tR{]����?z�@�ӧ�y��~�(<I[��֐?�� {����톄rU��sM �9*lS*�xP��������"���҃�a��M�Y')��~=^{���/�Gi22��5+�
�\P�\m�fP�R9��FZ;���3�[ �6��m����\��8_�@ҙ6�#b{����W�t ����PFe~촎�x���y��'&��u,���lb��P~�jS��)ݾmY��$z���	���Zl��M)�Fd=`���k��q�-�>L�.~B����K7����������T&�CkD��]���Ɓx#z�hU{�NJ2��7ǵR�lr������|0���?��#�2?���ݝ���dý��.��`h��\���k��%�ib4����7��AB�[`��������)�-	��I��;�9�u%wH R�9E����)D��=����E'�9��ި�}��Y�8�r��^d=��2m�ؖ�>���d���"'��4�(��
�A�D���O�g��O��Y��' ?��h�4��F��
�?�t� Jx���6�v��(��U:rCO��X�Ҽ;�%�����'̰� �d������Wv�xWd	�}��B�  ?,�f툩�L��Mq���V��^��$���v��:�9�v	$�j2,�C,z��ME~�G �T�����st��������j`r�5ܙ�a�,y�.�DVk���p����j���	}����@0+3uM/���r@��8�[�7� �� ]�����(T��j�Gd��1n�9��8�ط|����)�g�D
�M��0�-h�ա"�IPN
Rj�_L�W%,~}���O�=iTʲ>.
�5ŵj_���Og'*E��
�+?oe����hC��ȼ���>��O�M1�D����:���5��g�ՓC�5σDq��X�٬B#\zn���46�bd��<�|�?C�0��SR�e������g)-�`QB����{1&��n��b�"�ig�O�Z'��2~O���f:3e���F~�0?ŊY�="�A�����$6���_j��A��W/���2�6.���^�C	��O+f�q����l����r�)GE�[������00�!�>�٣wJ��u�'���?cP���A��*<M�f&;E��H��;'�U�N}cpH�l��&px(>]�0�� ��6`�b�}\#բuC�ה].,��C{D�<��Y���&�uKr�^��[�b���3�{��.�U�5+r��iN��(��e�yhpW��r�1]&�9��������e�bN�EP�Mfl=�d	pſ�:٢ؘ]?�i�z���k	�d[���z��wR� �`����x]g9����j���h�e��@��4?UsrΣ��|=B
�������:��\��>�G1/d�h�������ON�[>M���Z^n�R(D�I�?�fg�n���?���M�Z�
L/7�a�r�H�+��[���S�u�ge�r�{'T���rԏΏ���Mx
W{*��qoNU~�uY�9�I��]�^��r@�seu�i�:;?��)���^;���[kf�F���8�rh+��x��A7�x��3y�����]+��l�M���l�p|QlMx:G�nh2M����n�7�.\%But�Wѝ'V�H|%�}��ibi�-�UA*A�x�ۜ���Ċc��"Jř�|e
s�RB��L>I~�~Q%�����O�Bf୽$(�����"Q`����ً�^�I�!�	��}.� �j]t�\���]'�� ���k��(0-�|^�,���A�:R������q-����W��.κ/�;(GA�9WL�Y��} �~{Ѫ�o��%�����,�Q���zF�#���"	>�HC�5�~�hhsd�HxdՑ�}j�NZ�Kwbx�+��׆�m-�G0
UN5J!������a而݉���l"AjvӐ�|�OW�*T���/��e�[gh\(�݃��y�=�-¡�2P�bK4GyҩҚ,N��'�ً�7�5\p+�ɧ����@���H���ʞ/�<l����٤��� KY�� ��M�^e�<���;b�Y��Vdz��7��_����|zl/L��E�s|�AGѴ׷�Ύ2/P��^��Q��is���i�r)U໔Qx +:J��Uq�ׂ�7B�fYq��;ҁ�$�*�@��* >��B����%l�o��2!+
F ۺ���j�aR���}b�fM�κ��B���R ���*J���s$���r|��o'���~l�!?nN�`>�rB�됄:'#b/��֣Nc�1��C3� v��n�K%&$n�[� �˴�� N�~B�5����A����S�:���d�=�#<Q������ɚS���@���C�}`��$���S�"��0�h�<��@wT�����nxQ,���1kj�\���AKm9�A�j�+�[�8~�v�_��8�"�EuT��+-Dt#�X����w��
��H�9���VZSL�_)U��zV�/EL���9�y�Md�l��bvD6���q�K��E~��W��-r�����~�:�pGi-y�|/_ïx�����1�2۲�_\���[��h�%�J�5���Ud��t-��G����L�Ьn{"��y�zn�r�M3��`{�<��=�a)����Z���[�F�:a}C?`5���7|���UX�A6�c���h�t�j�N�vN��_Y�È�'wK ,���^�����m0��ۙ�]�|q�fX� �n�DRx3B8)��ך&P�kXx/��Z����R�~����zB��'�))1l���O�D�kb��`�%[�]|�B�20��ĵ�&Wyu���&*�J?�~ڠ��������f]��r]>"�צ���d��)����uD[h��K�u�9��_�}���mDY��R x�l��	�[��Ya��b3�H~���|3��]��aE���N�n�ח�9%��&����7@_Xk�a�"�-l�OK��|��Eg���}�a�'���Gd�]!���P�~4�y&&�߮HĐR>�Kn�fJ�8 �Oh.��yh�i�+�{L�I�����-<����fҺ�YPT�>A0h5�A	q{�HE��_� �8R̨��?��>,�XE�WϺX2_|�"|�z1o^N���Ԭ��pDIP&v������{CJi�V�<���ox�OS�=��D�+�Ԉ�D��#�RO��L�䓩�Ʃ?m`1�Q��5���,\L.M1˝�B�����ɑ�b���Z�Q�֗������_�����pn��o�&6!�lwoT���X�5���m�@��WF�r�^:	�8kC���5�)��t�/�ޢh�@���?��e�����$�1t��Go��rx�������� Ta�pG-c�����ױ̽67��:ݼ��-�H�T���HK�#��+߰�2gE u���\����;T�fߔ�.ga�u?BY����B�jvh/g�}�E���m�M.S�bPQZ���[�&�Za� ��n/>`ɴ��#��1�J���\����aA+,��S% �$&��w�\ 8��y���;j<�� ����o?��&�!�V�reG�+(ab	��=�M�8���oD��z�U:
��t�4�ܝn�}��
P<���HEnteY��cI-��'M��;~{�k'�*}H$=��OaS��G��?�:f��Q.ȟ�P�{*:tu�(5@￐qD�ޞ��q���r�m�tg�G� �p�7�[��U��C�_����]o5��s.SKIsU�UWˏ�8m��T��q��S!O�T��sF�ڄ}���Io��7e��!d#j��9�7�|ŀV�R�� >	�
�H(�Vi����F�r�4��B�/!svR܃�����$W5�Y��~Ҕ���\�K���$e9Jm�>ļ̠���D���l�QD]|�%��Z�8�R��{�H����D��y-�Z�&0kI�����	{� �Ɖ�0G;Ĝ���3D�[E���SZgb����X�k�����#��QF*w� �P��XL*���Y�t'I���7��Hl���f�y5��)�?�׫[Py9�s�\;&��c(�%���R�CC���	MJi�*�M����h(X�<��G�t�Ph��� �Y�{���Ù�[�Y��G���)�f�0�p�ݣ�-�R�Y4�v1���ŀ�nĎǙKـ�1m�� jǹD3�a�\�wx�i���͗$�sIY����L�֥$E�ʴ�\+3W����,����ۣw�@6��Z���b�FQ&.�F��6�M��㷪l����}&\-�sM6ޫ!oM
��Gk�1o���h�ǁFG d�wn?��*�H�.q�R�{
��՞�ԒH� ��	c�-�7�m�_���+����\��tE���f��:i^�(�ң? <O���Ӽ�(�NÐ���j"��l���e��a�껨ۄhLI}�ף�,�/������u�ɬ�{��ޯ�q�Z�Pv(��vj�=���y�PI�H ��vW3,O���׹x�NG\�f������9���tg��c	K�*�4Z�֓��MuR�d�	��lF�d�V~���St�c��E���p���G�'=g�͉ ����}�~���L�ւ��Q����$�����!|�4�vo	�ˑgq==%g4Q���#>�(T�$�!Z��t=W%f!���[����?����Hl��>���ѩ2�g�t�tU�6�$�֛M(
�xQVB9��ig.[�}w2��^&�� ߬�0wvv�+�G�=���q<'�
�:�{�E�~-[0RN6�X6�cM��I:Y���y9��f��P����y�N�W�F�}�vj�8ȫ�W��Ċ����і<[��ZO����,~;P����¢'[uf{�L�anђ��V�]�p�^�����Mws>0���w("oӯ��/��H�C΍������J�9�N�a�`�s�
r���;��|9ʷ�����|_�Ư+t�}�ϧS��5l.���/[�<�x�f[K�I��d��ߘ�h�(j�<[����r�5B�	*��������D], �������/&�N�����=��c��B`c�-m09�Mzo!�w�����s��cZJ1�׻�:�W_g!��������r�ɝ�����v�E�/2 �L��"{����m�܁ά\��:[t�;��7#5!@
l��bAÐ1�P�uI���:�w3�F�Z
����E^�='3�W�������wmH4�-b&���#v���zYi�p�'�<-�;B<9���A`w�ӵY ���ƕ餗3\�S�AԌ��Č��bqd������v���qp� @��u�(�Q��aWEM�C�'6��VK�ZU�m��%ҕZ%�Q�¶ix�X&,i��h��ֵ"�3�/�şy�q�B�A-$��{d	AA�=�O��?�5�9-�q��ϖZBj%���(Lz�\�kS�ߝ��vոG�7MY�H%���[�	��f��(���3=3n,&����p�K~e��ƭw]������%��,$Qf�R�F����議#���8�c�n]����6g ���Tg������.��p�)�&�'�0�5K=l9Z����Ga@���XX�GNw|��	<�vKA�os�V��ʢ���X��m���]��R�o�hbp5�q�'��P1Q,�M�=[�,���F;���R`�	��Ŀ<�4�\����ʥN��~)IX��ŷ:�;�r� K]&�S��X���������.�X��M�U�oSUH���6��+�2��r���V��Z�c�_|s��-��ʣd.f��	O� � ��k5��ս`��ufh���3+�>����Z��Rnq�ϻG�
��UxU��ZԱ�ϱ�E������_@ɗ`1&�f�j����\��K_�5�q뗟X19IN�ء�d6�A�d� �/uw��5�ʧ�f֥��bT�B��#`�k~jȟ�=�*���gI�AG�Ir,�˝�`�E��*������*�+=�����b�A��A�E5E
 �8)�g�VI���c�%�uzw�Ƨ��y3�8/�	9C�0�c\�PO��ZgSW�Z����u) 	�ujn�։�f��{\���@��;*Z�x�t��D<vG��;V����@o�VmQ��ËD�$��NEa+�ȹ9���Z�K��L���Ӌʑ�$G+���΅4��l�nA�.��>Fˍ�w��xƌw�à�3<�Ve%R�^�Չ�=7��'*|��^d��UןP'�;۱�eؔ~��M!2�]��䚱<��>n�)�I_��O��+Q�>þW�x��y��>�_��؏4�L�<�b;����Q��T1M]��p��3���'�	�~c(>d�jhV�z��`�,���Ͽ�i-���+�1jʺV]�y��]����@�p���q�P	�V��հw3���!9NeHw�Ŕ��U0��Q�cMZ�c.̸Ue�҃9�i�q����v���6��ת2��H�~��jM��y)ﭙ��$�L�	]����S�?Un�����)������m�\�Z�������J>�����&UԳ�P�&(�hŃWb�T������G�o<����X���.�
����V���)F��L���B2���nq%'|���Y��|M��Џ����2���15��Q7ό�pu�9�Ð �d�<���Qr��&���QR(H�z�[2��r�5��k
��Hˈ����0s>�n��u昹Kn*���l��ød�GaLP���΋����y��\*b�ͦ7����>��a�k�T[���[����i�������S�Q����N�X��W���.&P�O�3����2�H�����s��>�h�qm����'�����N��
��Id����T`I�S�����E�c���!���� ��A6+�M�
3�ٓQg��ۭ�(���m.�<E+:a�n �ӉR{X@uy�]�/�<5�+UQZ����pR�6�_7��p`[��GfG�#u1��u���԰�wd�G ,�s	J⤠�ܪ���T���2!1�AP4íc�M�ͬk���� x�{aq����AxFޑTlvF������J�� ��,�EB��Xj��گl3���=S�ʜȻ�g/Ι�M}��]L�[��"�%�G���m�����H8���z�3��8C��1%�%W#�v�o�8�/��������`Џ�5�a ����]�-��~�\��Q�9jg��A�'�zɑ����������\��AC�u�e)�F�ʬ�]��lhGz�A�If[Y��OK�k��	]� ����P܀	G*�SȮ�o�<<��ւB,�g�toF���׹H
��u ��;�O��(��#o�̃��M��ĕӊ#f|�k���K{�1?V,^Gw�ݸ����_��c뭉���U�Fb�6 �M-�U����D�G躲NU`Q�����=��Ӌ6%���
��{f��0��$"���y�b��\^P9ɪe������\AȈMt�dL,��5�X(��%![e�OC��\9c��p/�_�Vś�(sA��)7s�K� �P�DY����OD�y���k��O��t��]�+�����k��8G�t�vQJ��c�H�zP��T1���M!bTv�8��,��J5up�)d���d���h&4�{�'�u5��srI�FYmǺ��s�p)M	�3��v��Ƣ�Vq#
UE�,wb�i��xk��/1�"���^�&`�ʀ��N����fsME������u� �N6��1�B
ؚ�°��`�*��� �K}�Թ,�u̯Nw�0�ϛ��+�7	�}R{#�KT��g�js���s����Q���d�F��`�H��:��gM`�����ib���2��v� �����ox�\eS���cQ�5�+DCd%G��8��g���J��Dxc~<u�|������$9{=b��D%/}���M�f+����U�^�5��!�:{!L�zxԻp�=%WaX���4�ҽ66��=zvR
u�ə�܉O���gC�[$�ҩ���xZI��_������=Cd�MC:V-�#f��� �Z��;��I ���9�T���͞!��H�bm�M�������)~���0�Q5V��1@�h,%�B�n��%� �T���߅�
�q��&�L~�xZ��8Ƨp��yQE�Xo3��'Ⱥ�Қ�<�:%�[�gù�A�^%J:>���l�%�:�7+�5�b�v8���5�����7{��k�
�8BD�����{�Y����*�o���2z��}g�˼�$�Ib�$I<�+>gy�A�;��_�.Lp��_���!4�Lo2���:P���	�n���-����J�j*�H`�B��e+���6� g�������C7;^��sL,>	8Y�%�����G#&OXA�c<�S�I�L����c{���u�������V�kR7Q*�hDа�]����k^�U�E�-��ܫ<=�����T!#�-��A	>���W��|P�'�@p�O+�,W�"���Z��u	4��L�ǝ�5�c��?�U�a���F~�GYKt������$�ZB�E��2Q��8}�_	���>Z��(#5�K��6�D�c�&x<b��2���*�B:5�wc�7e���.�����-�2�8h�(�Q�=7j��'����^jby��� �sp��iιCwm�-�h�7ĽTJ2���7��ts\��N{��[���ί�))^�z��ǀ��)�TtN�+M^>P��[K���bj£�������F���G9xXڋ�=��ݻ�ߤ��q[{�q}���*&J��1�YI�a�O�T��K���Nx\���Hg����\��q��3�z����"���!#,�S�~��E�e��*�Ϻ�[!��G؆�R� ||��oٓKI�-�FN��'En*VK�r�s6U��%�pn#���{t����%��fs�%��q�	v�d�_��O@cQ+����?�o�����5�����bK��]2�����5ewS�ǒ��hfe���1��3����lI���PGy������/����F�3��?��P���8�����䥵�L���$��?�K�33:"��+�#�,{�ˎʓ�����H��#����U�iA���pm���d��K�Qk���������cT@�d��4��)�`竣?��\P�C�RPC��������!�������ݚX�����9��1�O����Y�L�=�FH�N��Q�ܦo�0l�	~2⹥)\�X�i�!�|�C�v�-.r����!^;���/y�����M��?�vBrCf	.�A<Q�b2�J��$��~�����/���/��4�� ����ؕ�ql��A�+s���C���o$Ӄ�T� @�dv��:a�d�N�kp�g����������1Ё�������cɱ��㾃�A��-�����aL�c���V�&���T�lX��N�,*3��fa��L��[%v�{��@���|��ո;S)�6>�U&x/ �a�Y�K�`x\�r+�+���^az����5�>b�j�egU�݂%��r.�{0�b�[{�@%���j��6\�<���.	="��԰Q?#��Y�H��6�[f���?��qu�6Cx̶.�,)npA^�@�YW�(_��.]T�p8Z2���>KCrM��l$<������KQ�M�0�w���q.@��k�Ab/7�9W�&���Q��o�m�g�vL%~K��Z���ίc�����S�S]@�y��)�wǓ{kTX���~���m+U��bm�)���].I�d��
�h����O�9�fv]5��O�]�����$�P�+׀�.K*;�iC��Uy�"��=J���L4n+����l6[Z������b
�, �|7�9ǝVw�_ڀ��J�ݤ��p���0����ŋSb"�*S�#�$��񙶞|���q��������G;�`��$9�іZ��WsS���"�zI9f�k ��Ĺ����36�U<hD�(k����̗�Y�Ş�	.����A`g��54� ���W6i�pڋ�t�T�4�R~�t�����t3�t�`'ߗ3��UK���n��}u䶩�ݰ[.�b���}1��([�4��4d�qE�6>a�(��2��oa����#D>��q��kb�CKB�O̷(��ž��=�7^4=۞�y�c�x��V�k
E-^��
K�v=k�x}G*2:X��R�G�m�Eb+?�U33?�%E�r�&_4m��囹�j�"����+v��Jv��Y��*>��ROMZvje���]^=����E�42�:��E�y�r���Z�q���j?a��%�4SZW�ur�����"���E�p�������a�ƻ%0�%M�_�z�*��o��IP�u���f2E0�fh�J���H��{����+^EX0���7�D��i��⨠.��<E~&hP� �Q"V�5��2�����nXi�)|�L;�驨��h�ӎl.(7�>4�D6�IL�����N����1?7]��B�-t�8:"WC�hڋ���o��}������oyq���W�j����T���H㞏�M���������b}!v���ZŐ`�!���h[l�؏�7 �"?)���b> :�U��G+ة3����r����r�/*�b5��cU���]���f3�$=W����q���	ݟ ��=��,� ��#8�����_��0 p�6�1�ޣ�nttj?+\���«�_S��z���K�G�V���&�ɔR�y�O��o�\F,��������,#���]'.kcD��i�Q��ҸK�@/���P8�v�]���ɲ}}?��<K;	Ā�o5=�3����*�$���R*�Ӛ�Rܜ#�%]����D�+*K���=��N����4�l��l�_�N��M���y�
����J������cRg�Y]`+��S,L�~�V`Eʇ�jL��~��1it�R�g��R�*�/�Y���;�/G�!��x��2Σ���F��^���͵�M�iZ�"�I&�З}����t��d(2uh��G�:�"�%U{>*?I���Eg��4Qo��w������)0�J��e��L20G[V�Ԙ�r�XQ�b*����I����vx*2��r�	��#L�֬�ڿ	�>.}kd�1{�Vu�
ɨ��m���3b��ږ��+�
�-��:U����-����C���u�c�R�S]q��8e�Q,����]1f}�ϋ��U��%ϴ�%��q�[#>������j��wK���0\�Iڮ�U�z ��t4T�Pl�H��eU}�]\�4tC|�u�G)aY����f��q����["q}a�s��?a>J������(��T������-0�êF�\RYXa�R��i,��z�������Jë�p��)�P.�2r�!�v`�Y	N5<���k����p���4�ny�U�X��H�??�B��E�@$�!X��_��Zu?�k�9q�k��iq%�}�aS|ؠ�����,�Q��ԱS�v��Zm�w�V
���ʃ�E�r�{u��͓�oh7@�X~��I1/k��Tj�ا�@�CsP��Ɨ/% �S�,z��*�F�տ;&�c�t:�NҦ� f~
A1A�,��*�;:���}�K��ѱ ]߻TY�����%h�|�s��]}R�;�]�
���s3�x�&���sc�=��0ۜ�e��M�&�	g,�[S���u^ n��`��ۼ����O���F'B�Xu��0�R\��Zoa g#�]�R&��,��b�l��)�W��[��-`Y�"�	�J0z����Zȵ�;���
N	���bH���ӋSEw8@] �+�v5ը�X�vǈN�.RN��6ɚ���S��A�U�;�`��C�I�MF"�LJ�u�"e%�ث�A�mzE�D��M���P��ߺ�j�nK��j�E�[Ê,��K�g�a����ܕ��څ��s��\�]P��(�'���