��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P��v�"<ߞ��&'��k%P碶�R�ӣ�sĞ������FY&c�W��f
d�:��s�WS�_ӄ$����(m��r?1���as��l9�����ݫ��˹��/���:SP�mj�\�@Ǯ=��
���������ʺ�F�G��o��p�f����E;t�df�� ïKK��Jla!�Z5k�M&�I�N6(���;�aJ"��܄�ܸ��G'>J9�╀]��krJN2��$kزז���ӭNV����4�H�:ͬ�!�9�#Xkz"qVL-M0vj��Q�!݀>�ҤK�,��wynZ_⺷����V����}`�{p������S��Og}/4 �)-��͟b���H���	�X¦T��B=Ό����/ئa�Ŝ;����O/��t��%6���~)q��j� y�GQ.O��}����=�H~O�^'�,��LmI<���QbA.������1�
Z��2����<�5~ac�b��dz�j5#�R֭���v|>�=�O���Ľz�?kR�X�+��`ZV�V�%�Cw����A� �:K+�i��=kqcZ"���FrP�� �7�6P��37��L�JԜ٢�ǥ}k,7�0��7�u��'��F%n�!�Zҷ�F�H���-	���D��'s�b�}�1QO卶��2����.�#����ɉ%U�z(�7`�-2����A��"ӻ8A8���Rs��ei����m�g�H�M��P�j=�J�#���*�ZɅ�k��:���ŇV�B�ª㉐��e�O���f'�>��H����_�y�+!n�#]�8tB�z�tn���,��	Pƨ��jyKt�����tS�=�0^��KJ3p�������S�3;�ߏ-A�9C��-�7g�EotTH�,S[
y7�� 5�K9�g�MӝÖ�y���#9(f�Q�-c ��K��K�W�����Я[�^y�?%<��8��x_x�u�_�W�Gl[.����-+��M&�	x�O5+A@04Oc橿����Dʻ�(�s_Hq���j�U�����$�����c��-��M)&/9Ю�pt�y�D�D#8��a+]���8��`݌G�E����u���Τ��?B9�Ib0m�����
O����>O"�5�Wf���[�"������{��уO�a���y~������{��Ũ�B��T%�����7�:��N�\,��_rj�d�C�kQ}� 5��S~���L��
�z��~�E2_�؆<� t3=[���حG���+#����gէ�r���Hyvi
�>ҴɦE��6"4A4-����Xw�+_R��ơ�OG�=��������!�� ���r��7��b8յZ�]�����Kר��
Iy���'8�_�c:�@h��ĂnKQ�@��7�s�'$x�mlYk�dp��b�C�֜F}ӐoB���#�佔���J=��q��GQ�P Ř��4�!��ʻ0"x�M�/0�NV���m}�,Go9���{&b�����8Ϥ��/�9�l��
-3��R��uh�z�̓U��k�S��{0�7d�RTm�ك��~�����r����0f���X���*\�3�I����l���ߍA���� m����H�<)�!@���u�Y<E��Z�{p�g���&��g``�V~��iPەɱ�K��J�J#kC�2 ��[4]+I+�e��[�s�ʖ	; mor�%e���yQ�ɅR�:?�K�l��dl�y�iV,�LH�QW4��c쥹3�W�WUN[2 :���e���P����v�F�p�7�X��CڪNo�KP̄�qmi�|���%�/�轍���ڬ�(8 E%�W���|U�M�U�t.�xUbI׆����Lg���,���t�?A���	�揿0
�9�:(	��ב�c���۩��q�.	�aY��H>����vZ�M<�~�d��A�EF��YV�C]:&8%�zb,���[@S����ًU�Q볻D%��y��bd��,�J˙|>�a�p�ރ��K��r�� Rk��C准��P�Qʡғ����O����~t�"�3��+�b��������G��M�c�p͸E�q  j�p����#|��W�*��덟�!�����<��ᷜ'�H�7��[u��hp�*����$V��߇9�����dЏH���~�%%�4+�'#A]�!P���ʔ���.���E%_�6�p1G⾹������2�|GW����Z��|�~�ZGe0j���"��h=*���x��ɓy>�D��CF�g��8�طc?	t���#8;)��7��j�y��Z@�����f�p�bIcGUn`$`6��No���>�ldO�[q00���PB��c�[A��x��1���B���ľ/x�-/�@J!���X�8H��ȡ��V*���9í��Д�\�xM$�~/�<�!!��w�0=����<��^rَ��N_��#b���uY0��4�]\3�(}���X��.�
(9GK�� >IƠ]�Z�p|,)���m������D�W{fb��1��k���2ֹH�חh��H�3��[��y��0~[��pt��6�0��Uo��Y�l��9�(��.e-�pwאw�^"��89���OiGf��X,&�>6�ܺ�_���ʞZ��N��a�m{�/���WEy�ncz�t#F<&)����8f3&xc�Hnl�F�;��+A9��� X�3�--_�Ӱ��R�-@$�FN3�3z�M��%Sc�{�mq	��Y%��9�5����$�5��A��[E��/ע���H��v�!̿����R���K�ň�7���SH��W�hbXɋ����	V�	^"��S�㧗p2@��H����5s�cW��u��s�L�'�6e�JN�yIBp&���#�Q��|3y������$�j�������Z+w믛E-0�l%��}$aJ��5cJ�>��ljQ��WΪ��Lc�?W�h��*�v����p�����@�0cf�� ��л#f�;�p�ߤ���0&�H�'�5��[��RR�X�`8���cn���J�*�!�m�N���Z��EO�=M��AX6�je����{���@h�R"o��Ȼ��(�;ZPL3J���;�Ou��dXV��{��@H8���ҝL��D�J2�d72�� �՜;����]��36��:枷��M�UWH~�d�,��1е��%&���<&>�Ɛp��uL��P��ۓ�_1��s���אN޽�|؈pͬ���'0��ο�VRE���D�99�zZ�M�l��L��ޝ����4�ňp��	 �S�������V��yC�O#��ciW���ڂe` ����;B��D�	�ޟ��y��q����羿̏2IBix�����Ľ�b�f˸�`�6�\Z�HDc�G�W��QG��LV��!3��E�G����hF�f7gE���uF5��rsTou��%B
{��ޚ-�ϴR���ko��tc����Uns���q����T�-ic	��sE��}�l-o������Z�����4�j���|/VayP���gڬ�!���({��eu�$���F�&d�_{:��ķ��-�Zi���ݘ��7�tM�z������C��tT�"���]X�5�:h�M�[�ܻ��+�W|WM]��\�!Y⭚��qK/���L���$�v���8%�x�x�aPZ����6���[w�~��G6-6ҧ)fl�&�����F����ti2��g1�������ߢ�6���fiSj�M��|#б��s�v����єr���_�*4y,��RO@.��֍�kV�;Tֳ.i;��)k���̞sd��(�1܇�$�#X�����)4ԅOv���RP��)	ܸ��E�@��V��qosE���-7&U(�X������^�@���q����/^�BΛ�ɝ��xOC��n���iԖ5`I�NQ6�;��)~Ԡ�sK$&�_��-3�W*�R�Q�
ŝ>�]����܎0-	#�K�QHm���Z�>=[8,�%��~j���g*flg�+��/BҢ�0"��?����:ħۮ,�d*���<�H���xn�GR������g�Ω�y�m��E�ì+�*�~�>o.��\� �U"��i�GN�))'�68G��R �����}�_s�
��f�H�k"D.ul(���>��(���	�����vN�1������q��\ �x�K�������r�����1܊�2�ADõ��T�%Y��/R��r����!��_�}#�s�s���w[��-���4�����f1Dڷg�2�;9����v�\������fJ�ҪyR�~l�Y�#��&�����ȣ�ŴC��Nle�T��l��B������`�������z����uhV`]��;�
�m��}�P�r���:*�b��\�(���9��y��ö��R� IY���������{$F���9(��2quZs*@#�C#g�x��f	�4>������0�!,��̨ș.	���zZ:�_=�ͳY�i��e����&͠m�\w��I+jHDx�����RD��b��}g��G�`�%�"K��1�����ߵV�t�$$��I���O�¸_�PWW���)�>��YfJ���C��p
�|��ֲ��#բܯym'_�%�[��lE^R�V��L=��P4�֧�)[��OW���q��<��!�ë������l��-�}ŷmU�S�9o��Z��"so.��Ň3��Wjy�Q9?|��N�PQY
vLz��(#�����׮�	��:�r�-�k0�ܙt��'�K@��N��r�[�
�h�AVӸN���؍��r���� �R�ѨPi�r��(���T�ZT�!�̤]�i���Y`��0"��)͍�2�:���w����J�UhJ�ex�$>l�?��bnSe/��I�l�Hb(i��� �Do�&�˔���K��8Y�x��N^�;y9l��<֏3�I�}���9K�Y�3���1ژu-M8��t��kj������f��y�[;��:���k=(��װc�Ѹ�9��H�f_N��a��[��p���`�7+����=�{�Cs�Ѻn�&�Wd�Kt�n[Kth��b��Y�9|
 o��/P(��)������-�P�I�y��p�%EV�۔���p�m�����8�V.徰&k¹�{��E��)aSV��Ml[	�tnMWq��-�6F�"�	;̂NvZ5u��(��ϔ��9�ȕt�����@�A4�*�s�[R Dڢ񸔛����?5����PZ�z	�D�A�*d�z�[�U�^:�a��&0�]8=�b"�a�Qʻ39""<A��B^52��v'.,�.�����ZΡ~I���v�:3v�?%쌆��%H�����x����u�6v�ܷw~x~�N'���X4;`�T�cP���<�Ƹ�ФG�RJ	���m�v�L�zm<�>���d��[��U���^������}�y�T;u�hX�i	#uN(�Xn�4ık�ϙ��֣�*���.�����U�]X�?�3[N�����H�Ou��j�x��J�l�!�`�'e]��Z˵�r�Cş'�� r7-H8REKL�^^0Qn��QT'�i�h���[�Sɀr��i�7��k���r3 �X�n��#�jX��nջ7{d �vפ��n�~��k�]&Y+8���X��'��� =��|�G�^8�T�����/�{�2�0���K�~V2��]�b�ڴ�BUTI>�1�?le��m���B����aY��l�Ͻ#;F�޾���v$1�1��9\���!�}쬃�YE��#s��[��:!˦���4��צ����p��p��}�L4��8`����� ��;:���������g��L��w��Mwf�z�-��g��A��\m��>K��}��M�A�(���� ��%9x\Sx�����NO�=�b#�OCHd����2���?��h<)���OѶ�/�� ��=�/<�Gm�ԱԆH4UmJ3��'����� �l�)I�&�̺�&���Ҁ���l��ۆ'�ww�a\\ݬ���ը+�ܲ�Ǔ����=����,��3�׬�7�M&�b�nS;��W�ē�3V��U�m$p���,)+�]e��ē��7?�!�U#n)��7�{%B����2`��mTC�}�����VUm̄�]��,-0�# C���E�Ż��cts��o������*�-L�ru�tR�Β�c�:WGsXOn6�
��5j>��q���^8�	�������߱��W�6,xp$���P*���_�4Q{/)�l�MH�X\�X}��X��E��j���YKv�}W�^�����Jp��\�{O<���0j2÷�2n^Y�4�n���a[�2����%����Q4���*gZ=֟ ��9���b�}q��Y�׎�u���it����/PG�C��?G:Q��<�e{� _�U�-y���3�~�6�F�&U�~�K�ir���1_�Zۍ(�c��"���S&3^�ɫ<q�r�Zx�y��H����Vѕ�����S礍��UZ�����zZ������/�|7���:�ڴ��:QaC:A�f-��-��L��(̮�%����¦N��K����Ei%��&��o�(%����h2ds�[;�g/�6rܾ�����% �oN��}�a�]A�C�RkLIo\���b
(�JQ(��'��FB�k���0�J�p� ètZ�z6�=/&oV`�q�<��`3�	�S����M�T�*3L�O�d[�@�}�#pA����Q]':���$���g8�`� �k{���k�&Q�Ht��e,�H�Б��(�a�(!��U2t"Yq�
�_�`]��0G����=%�0���������9�n���]w��$�d�W	3������%[�e������;���LA
K$�Ƈ X3_�̕�wm!�6W�ET��. ���.�t~iˤ>��f�q���I-�؟���9��~�3O�A���wH/	�%�(�n��U�w�?G�
|�"YmOKN��S��nԲ�j����3B��w^;N���@7����f�M
Sڌ.���9�]�M\�*>g�d��q+����*�mq-7��(��5ݟ����A
!�霛��mj����1�r�Zr��ۋQ���5�4�)�T��$I�.MP�ݞ>��?����@扌�������%�ʤ�O�e������mR �ˁ6�@�94�~pTeb�s�Ȳ��6�к+���r4�cX���|j��@Ż�C�R=hA�����7��
�{�#��^��p1�:�^(Fe��ʕ/D,�M��b�o�<��Ril/2@�=g��J0�g�ɜ[�/Y 5��1)�N�-|������oT�i�j�k6�����X�4��(�$��H�����9u ��2KT6��9s�ͥz��Ɖ��Y�Tkl�y{�Qt�x��0@5󨔷��e�K����vA�����=�#M͋4 ��6m�fT��)8�7������ͬEh9q6�VI�$�}���
�)`k��X�ݭ[�>j��+K
��>�]���	�J��fg�V�������(�z�Ks2� B��/:s.�I�o�ʏ/��C�K�̳P}<w�w���9$	!����GK�q-��D�P���g$.Ґ�׸mE��6H��i��~p�h��S}��x�e���2����[�=+��c�_i�5�Ү�(.��|��*��c~
��/��w`��}z{"-.@K���o�U.��N�`���J1(u�ӷ�~\!#��Id��}T���ds>f�:�	;�,Z����,	���A�Ⱘ��[PR~iC�c�)^1R
WR�·�L����[W�#�y;��= ח��t�������~{�g��#8���������� eE���^���*!���D�T�f��'���%1�9[����LM��8���]NV��I�at\�)_�4y���X����e��N��-���d�|2�K�4�?7����ԯTiY8�I�n}4=����͒��xy���[/���	sdK���Y�bA�*	K
��쁞#9xS��n�{;�X���1���.sF�͑[��s|��e�ѿ���kL���+\��PQ���
�"�(��3�R�˯�5��"��[J��!���	�	��s�kg��+�M�V/�W	���*��t�{hA|���j�p�^Q�0d�L �,j#&��v�{�W**��_�G��Ϣ=P��9Z_D��)�c��H]i� q�6�*��(K�����^�&�l�t��鲃��k�Q#$�E�"�j�{�
���1�U�+��h_L毮�c��;p���>�o|�\�Ȭ<1M����,����x���<!������[��V�8�-� `����_�Jp&í$��뇡VH�L�ҕ��5U}����];%iIC,�"0��u��'��$�2���p֣�5�*��y�X�^�S��Қn�
&fdK=����\���BX8�B�
8O�l�Dpa��~�|@q���G�.�4��ȓ������