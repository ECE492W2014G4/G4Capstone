��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P��v�"<ߞ��&'��k%P碶�R�ӣ�sĞ������FY&�zH����/Vu�T��+9&$��2mN��5AQޥ�J���Fs�$tI�"[�:aCL{5�"�W+��Bco� �%�DL=��R��ԥlEb^�g??bsd�{2�hL/���ot��u�N<���%���V���ͧptRAib[ueӎ��#�ғV�w/�F�D�a��xc����>�|�3]����m�k��!iUG���a��t	d�l�>��)�����li���y���t<��-��K�I  U���_L���SޒyJ�����?��,$#���\!)('ʿ)���Cwn�g�D?(�~�&���Q��X��^k�3�����ַ͝,�86;�g"l>�b����+=���N�,�b��</++K?��{���� �:Q񮗇\0���~Eǝ�Ⱦ���J'�3��\�+��<���e��P&�󞂌�U@��M?��<��P"��憅�s���Q��˲���	q��/�}���������K��*�uZk�|�ljUA-�/L�=�]tj�9�k��]i(��Ҏ3k��xƞƀ�l�![ <_4�KS2�k�J��go��
�]1$b�'S�z��"���N�C�o�����}���/�}/���� j�[Bg�q�>����Ԕǿ<Y�{�U<���k�c`�<�}�^����`��1^�M�e�z�)�4)B+�dQ�2`Dv��	
��tº0as�hw�?�3�����l��6�š�ss3a߳�1�إ�ΏCY)��'-T����wE�+�����Upq�{E]F�s���Rn����U��z����>j�	�z�р�<��ذj���D����O&��U��O�5yhfW�D�H9HNt��U׵O95��88��PR�����Q��7�>,�u;2�! &3�Z̼�%���!�*��ś��u w���i�����V޶������������NA��wd�>�6�v^��q�*"lw�i�$��t>�Ā�6�tS",Y�w�څS�dR�0(	�D���~J��[#2q�g�RR�:�s�)�Gي����fÈ��EumSgAUK�Z�3��Q�b�KtE��OU]R�OA���0�_]�,����Ep�S;Ki���>8�Q^`�ɸAA;�����ҸXd���g���.1��0��X��/���7�x��Z�	�O����B���t>��@�:�ç�#B_r	��wI���!�i�W��?����3Lnv��v�!�%)��1��e�;Mځ^8�᷆�#mw>7=#��;f�?I�³�h�!+//�+�)S�>&���cBe/Ze����n ���Ժ���V/�+/)����G�i?���o�x#�-7)c�b��+l�Y�Z杻�n�G�.C�>��|���X��<��'ޢ,/��a��~q���͌�H��K��������㺋ӑ�t�DE��:X�-�9����G��W<�?��%�-�O���N�a]�-sh�/2�7ӆR���n�&D�D�t�J�p�`�&#/u�t���(�G삭$�d6Y���U��j��Ѯ�D}{<��/l��������I�h��Xg�Yu�v�r��&*��z�ߕ,�{B�}��e�I�DV��R�bP���:m(�I.�}|���]�t�o�̧9��wQQ��^O"�dtŖj��	��o��|�̡v��X1"����9��%��^?֍[@�񼳼$���\����U:�7���v��o������-��1�߹=G�~�rCu+��$�
�Gz 8���]�6|:�.N�4�}-���Jx͒� ��2�+:1��j�`R6��~e�֧9��T���|5��
�֥�$�9��n��OZ+M�����?�ķ%mR����;���_ǿ{�2}�{��v�1�e��#��0��q�%��YoW��_�c�5M�J~�漶���3�4[��)Ҍ��Q�[V-W�7���3&^��-�y���d�Кz�UL��ꚡe�{K�5_i䉜H����6�5�F�8M.����h��v�/,�FoF�vpJ%a�P��]-���e�Ks[����S,cgS�A��P�<.p�i@������#u�_ŧ TH�V�z�խer��E������E�3O�?�6Ѡ�~���K���-Z��3G��,��\���)�j[C�im*�ւ��V �G�H���K���	��lp�e��0�@���q�n���	������:_�Ӫ�梓�j0��Y_�0i3Ģ����7� ��zk�JV3�������si�CԈ����iם���5�.ӨG�=b�`aդM�!�8M,��J��x'�f~�x�t�MK��xj��Y�/�{��T\<\s�Z�=h�������6
�l���l6k�]4��\��&X���K�Yop��]wbQ���� i�/�u�o�Q+��$��ܺ�@K�����4�d|xk��;2#��'�௦R��4�
�D����O5�i�m9n�%h����%��aSu/��M��I@��x���V��^�ɿ�����d��w�3] �m�������JV�T��EV�S<�_:��;�+0�۶pH� ��m�p-�sY�^nmYD¾�F��"��X�q���V�����~��L���B��V�����a�[����"���;�P%�l��=��#`�
ԟĽWf�;lS��٥$[��#��!���%F}E?�jҘ|�ɸ_|C��`&Mݭ��ٮ"���m$�u�0q;��Լ�����dG��ն>F�?��1g��p���n�ZS:o3�Ǎp�f�g�n�V5p�G�2Z��#��.9���foePĿ����O��l�e�N��Y��L�<r.��1��)�h9�	%Z\�ł,
�E@��H�2�&�,>�F+�����uS<Ғ��,�ڵ�|f�tb;PB^�ITxD6��	e3em���5#�ۙ��P��;Df�O�(`�h:鬅�T�*o��N�&�]ެ������ �)@ۿ�H�2�4��}$&�
Zz� �1��cuu�9b�<h51
��N}��3���t��J�|?,���Nd^s������H#�x[)�H�d�(�X�[yh��{���&���F;��f^P:�R�R(�^~��YV/ܽ���.�xt�᰹3
tZ��:��L��c~�b�;�^l�� �+w4�Q�v����JÇc��$n�Ci��@���V�^���z�ˊ�v�#�7�^r���oTԐ�~���\���h�f��J� ��u�V�9�F�����d}Yn�YD/\*��\Y~�D�{�$������]�Q����I}~uԱe���/��X��l��0�=g� ^��î;��m�S �a�t�+q�k�\d�u�����.���i�uCIT��XĔ��dO#Н�U՚_$sn��E����a�2�<YŮa���k�`���[1^+2�I(�ʗ�09V"��(��:#�
<W�-X^�ލ���>�#܏��M|b�2������/ؔR�+��`S������Tjs���ڳ$�)����ϖ��3g+h���-y����r�=�rԔS �,��Г	�[DC�Bb
��\%��	���4$n���62�y9�v���-�T	�ЍY��<M	���>�.l2��|�G�x��6R�u�$� ��@�`K�� <�:o�''��*�PN��xS����/i�v�+�\�G^9miN�0X��@S9vo5'/���Ʉ��<4�U?�@$�$�?��.UҌ ��ή�86��-ɧ�^-;�_7��
��@!�S������NAak��4����uN��`,��;Qe�%�F�'i��o7�bq�{ZMJ��<�
"ʬJ��e����ύ�߽�%,#3kBj2N��4���H��>�T�,x�<���_�`�}��˸l TY�:lamE�@�'lGc1��A��@@ϋe���'���9��<���A�a�w���c��K��QЎ+����Rc=6�pc�;(Y'�I]�@L��tO`�!0����K�&�X��i�@�r�=X�aC|\�g(���U1��G��;D��o�����<.�gȔ@̝^Rܯ�Vn�$� �| �9��s�@t;ht�KpU��$,	bp`E�m�d u�"
����^MG���. O�H.���N<\Sdn���ǫ$#�I�M��^��9xw��.O�m{K�80���a��nq.z�޸�&���K��^�Y̑������(���>#5i�>��w�㜨�ږ �k!E��C��:�(���2����jz>�}"|7�D+V!����4i���Ag�_���\�|bu����-^u�"^QZ�?#21z�>�?���]���G�D&��m"�ż~�z�<\I��z������?����N{��@�-����a�,�ﬦ��b����Ih�����%�/|'L0Z6E= ����
�=sC���.)@��K�>�K�&d�A�܆Y@�Th�j�?�z� �x]x��<=9>�Jw�'E$�%��T��7ū���i���ج�)�9��:P:�A�bA�8TꙄԦR�������t�=�T��.e7�P����}�9��F�&]��,cҬ���%=S�h��L3郆���~����~�0�I?�n;c�P\i��#�[�O�����'�.�c�p?o����k��[�Xb��&�1��l�8E��>U��[�f4ӗc+�������-�݆ʝ�����Ū�	���l�OĠ�c�#��0����$/׋��J�;��M~,Kh����#*,�e�ZCM*W;��4 4Z��3@�JH�1��^ջ�|5��zۺ�j��)�7�_M;�?��Z�%b�/���C��Z���x{vx'*@��y8?���]�^��T� ��YƗTa,�Fv9En���EC�p<��MLk�gdqɫ��C�g;:�){��	��U��B�߯��?���R3�޳M�J��kz��l_%���HH����#����:���:�馟�h<X���$Y��qp"�np���#�Z�b�ϰ��J. ��"�R����8VtUa��`�A�I��O�6.��f\��Go���8��P{s�,�'t��]2L��l��4_��Õ;��(���a�3�[oI8W)��>M�X�!8s;�#)b#��H�|���)�`���q^���c�'?��ϩ��>�y��e=5��T���V�G�	�D!�t�S�K�sp���դ�+hg�p:R��/�#��å+��:�}��G��w��N��^~<����m�\��SHs:^��z���&��� j��h1g������Ղ���L�ݿ���ݥJP��P�X�SK���YJ\282C�f�Ω��gKaܓ��	b�L
j
�L�����M|o�<���>�aDґ����9���u�V�V��B�g��E�9	���
������t�~��20����j,�]K��I���B]��~�̮ߵ��e��~6X}�<�@���mH6j|�J���1*Z��8��X��Cp���be:�8�Ѣ?�)�$���WA��D���x��H���{N���I0��!S�J����j"Z�i�{��-`�dl?�V~���[@{�T�$7J�pn�k������� 3�+~$Y(��{�����|���l�a�>�
��E\\���PfW8�Z�'s=}�/A�i��y-����M��߯`�TD���J'�9%���|��&�q�������g.���$_��)�����J�yU
�WiG���n����)X������9�J1�l$7]h������5�?�I>��#�m$�֔�Qb��+��l�B�����jky��l7)�A���b�ll���+��-ji�hH�¬���0��Abm�\���ve�}@�� ��`2����mk�p�X��bY�l:W���<�ƙD>#��	�G圞f( s�c�V\��>��,��k%m?���!u���j��$z�������b����p�
@Wȱ�e�x��%���1
p&@u.���8�L���_*]!���������鏁��f�Ȟ�F�WﭮX���o<�R#ׅz#�S�W<�3��\=�r�릋5Mȑ�?��BI�O�7K0/5'v�h�9�O�X]���������(�b	bX�D=h���	���w��9ɿ��+!�=��<�|�aβ���졯�A�p]���l~���g7ph��) �4Q�F�G�ڦmS`:;�Z�L�ɢ&	��J޺��h,��G2�j�s�9���#J�	f���Z���ք��7���$�/o��q��11e9H�<E�+���6K?l5���� �BrJԽ������G�k,b�z0��<�^Ұ�H�Ro�|�z�ʩ\ˀ�:�cj���o�\�U��n�Vî�=�NI$�A���8Y��	H�M���0����'������E����	l1��q�(9gG{�O �
N@c��Y̽y�h��g��uF6���0���ߐ��6i7��MJ���ދ9y�}�{�hXA:-k�F���[ZP���Hi��NV��v�q�������MpH���g��nh�:씹A������L�l�k%�	�Q��,L:�huV�Ό�*g�0�~5M��~�6-<�SD;۱���;s���p����|�Q���&2���j�BF���=�lw����h���~�� �cb��&Z]^e�r/���0�fC��������Ӽr�]w��GK�~&�{ �Ƈ�Ҡ�������&�
�~̰�Rtf<mZ��2���E��nD=ߝ
-Ǒ(��└��,׈?��W�K~4��12�&)�Li�cG��Qb�6u/�
���G㑚��stHO�o6w��q�]�����������^�\E���Gր����ˀt����:o�Q�h��5�ۉ;��7 ����[D�;�����u	@Y_���M��<� ���W�E�j	��*�Q�C�Nc�I_h�f�U0���@;��cE���vC{pO��я"�J�I(�v��������4	���zL�Z^Xf�l�_�?9G��Ѹ]^�Z�HL�����K69�HX�2R_as<�B��*�� 5%{|&����kb+U8��w��=�X�m�L�KP?}}��%�Mv��!�e��j������PKB���e�j��~&�����j��B�Rp�����/f��?پH䇱__Ɨ���-�xʿ�7,
�+��4�g��*>���O2�RQT$�Q�d�q���yc�驛 �7'wߴ��.|�@���	�&Aj+n��5��r��#?��d�u҃�w��Os�&�Cְ�CJG&������~�Ճ�"@%oh���+e���4��l��K��l����M�$�hx�F�pa���C����\+��D�z;C{ء ���8 .H�T������ʃ	p�})��p):�g�*���	\���0ǜ�<����`�l3��eHx@k�ݨy@��^����l>�WF��2 �`���p<B^E��v�ă�a�mՙ*���m�/�3^/�1ق��',�������ZvGYnA=�ܤ2w��_<�����z���]�ib"uG�#���D��t���h��~�Y�A�����@!�k��KT?5X�>g���� Q��k�"dt)�n�%�����Ӓ,�M��8������D�}�^��k�M�p�3�r f��)�6|�5�P���z>����qu��Z��W���j�
eݥ; ryqif:��2Xߜ�[�nvpȨ���0.?t�68��d {�=U�ņ���w�;���;���A�\&pm�r���m{W;�$�w~�,|�1r�@��m���}�M���<��y(�*�RF��VT�d��{��h˴K�֦�8*�m4f^��S؈P�A�e�ЬZ�D��$ v�
��$�cA��3:d�@��Y3��!j�t3�:O�t��r�T���������>HtWN�Y���_��9����xn:;�y���K.*��z�ts�j�t�h�%\���r`�������d+`
������ 8�m�	t�� 7�AČ&�VKQѓmjJK��ۂ���,��+�����8�����XB��4C��q*�d�FU��!o�5�%��ߜ��%E�VT��>W�_��Tz�;!�%U��yy���(\T�˩q�&!�����~��h�c��-z��e�$x�n���c�أǮ)�`�]���s��"":�|_-7�0�gk�Y.
ˉ�w�NV�9�	K�p���NO�
�E��͒��X�V��6--mI���%"�iHk�k�4�c=� L�3�������<I,�����3q��7~��Ь1�!���s ,�����B|�ߒ��V�lu�A}���
�3X��.��-�1��*���g��V�Z����F����%������.�o��w�=b˗�Թ1fS!���8�)���C]8˩�z��@�u(�)s/���K��p;�)��b/ԿCT�j���?2w�1��(��՞b[#R�`��xr[��s<�۸�D���wmx�X�|zcCX�8���y�$�d
��I��o�Oʍ��3�$�|�ӄv|w����	��/4\F� 7揷� �F1��גm�����8��:����$6�=��f�@�D�/"ՓP�d��0�Z^����
9[�z�J�V5�����IqU�:=�N�����0/l��L��r��+�W��,�E�8��:���U�Q�������>)mi��[v������آ��,�,��6�̓�7dS �H��hb���=��K���A�$�*�׈����$��]X|����Xik���^�5�ˆ�$�vGҢ�щ79P�U֧��c�I�a���~��珑���n`$
ߜR�\��KS�w�7"V�E�x�be��f]���6�A���������|���r�]��� }���7݇��bJk�?�s,W+���o����[�ޚ�a:�]�+��b��y:!n`��~o#2 ���r��v��=��i��������C���^8:] Goŷ5f��mě2�ٝIE�(���f���u��[f�dG�LW�K�$�gHy�K:��a�����i���O��������l�I��%��49�L{@�`��>����1����[C�J��H{�8��Mɑ��D0���Ď�8ŏ?�8$��)���O��:�MK���h�'vo�L�S���NT��2j	�hn�O���{,`��/����+�z�qf6�	����ti�Z�\��!�E�_�>�8®����v��[s���d�͐��I����Q�{K	&�+)T��PPZ�y>[�����ٻ�A����ձ����f2A�֕�f5�q�U:����+t�{��7~F�������$��z&?cj�Xk�Jw�v�0}�X�|j�#�>�R"�Z%�Q��e�-�����}�c���~zfb�hug�uȱ��Fj|\�\t#	<��͌}F!���T�x-�Z�X�d��m���yHryS��P٘��V,ɛ��Z���+�{@�A�<I��Wr�t�H�O(-���>#�̡��T{�]����݅��c	 Z{<&(�����N����L��=�Z��G��¥?�>i�sf݆9��fH�tF`�6���y����3~�r�C�L���'�|D�^�["Q{��Q*���C��$�#���+�R�1c�+�[�2~H�F:'�*=�^�
E�'� �6�CY���T[�R�7���L(ȿF*�F�֊
+3w$����e�r5��M���[8bp<I�Dة�B�nO:�[*(�T0�߼���X�r���\��gM��x�������>�:# }"�27�K�����kk�lVOh����(p��N�;�� ~-K�5?�����dA ����)5EڒU�;U[�`l:��ז�H�=�
�3!�*s�s�pGq�ի�Z�+1�
+~�#��᫝�%���� ��'J��n�䎣/"p�u�*�%]|el)�Q-�d;��?;>��d9{c���ޗ^k�4>C,�L�|��3���l���Y��>[(����X*����|(�2�a���\�Z�?�Q��ٚ��8��]W�C<뗎�vXcH3,F�Q��m�+���d�,�,��ơ]�0ZXg�~�ڸ�K\āC��!�\+4��]�w�s��s�V:���6�\F2������3vz�!���CW�����}0���$
z~�@l	 �ėQj3i	���r���S������quq��&�
n'�����/YG��Z���9jp �]������m��+ζa�a�#%J9~y^[�t���$Τ�P�a���K��+�V_,b��HF+��@$�84��33��FC���-(ױl|=�Z?U����Y�*<�&��,6�L���]�B#7�t�I`2&鷇�@�gsA�x����o�S�Kt��;�&e��h�HQ.�A�\�%kj�"�\�!��c��'��+m7g�U����8 ��R����IՏ�J�6ᰕH��4I-�U��9�K`�����fyb�H����&vi�!.-�&ts�ENp6��PJjm���D�����U+��/Hv�~���m���ꛓ����g��, [#2��s�':]��L�I����a��=�or4�\��`Z�C��Q��x�?p�&j�镨�hKA���Gc���b��>��!k�������!�ƥ�)��͈���U96`�̘���{D��a%|�z�敾Sǟ�p7n�'�ש��Jz2�y���E������C�y�)�+�۵�JXk�*N(Ɔ��.[	'R�s��oSn���rz��92�C=�KM��E��-�#���K�@��j���%S��V��¼U��ǋ�lJ{q2Z�p��TI5'�u�f��Yr8���7F'P;2 ���v�$�0m���>7p��xe���n���������Z�{m�D�Iq���)�i��K�z�T����d���D3WW�yxi���Q�쌛���m)7��r�T��e��Y���Pˈ�Ql�|!�e���Cw�b�m�[�hi�Hj;��	�H�|��=�`����}^D#N ���p�ۭ�8�[v���GX�s���u-9כ.W��@��-(45v��Ֆ�R�<�綺E�w���L}ӏ�Q�u#o%��{�z?A��� ���Sքr�t������	���� D�rg}�L�P�6�O��n����I�z�Ig��D�[�����d��r�G� cV�'�E޴�+�
Ɖ`��53M��\9!oI�N�(c_W����G�:V0u��*~����S�D{P~:&-F����~F�^�v�]�T����,��̈́sS�Cq��O.�΋�;e��"���CgV��̓5�F`񟆤�u��6]r-�����-X�f���gfV�����cq�Η��:�0�)�!�S��Z��r	+�;�8;���Z��oHLsj@�)q�i"�tqf�q�������p$
at;�@��m/�Q��>�^�U�gm��T��#PU��XxH�=��Ǘ���=�m�(�L�7Ce�9B����<�h$�5\�ʡ{��R�� �/dwSd��X�K�cU�����=QJ�d��B�q�⻩/�9O%b}a�1���d�9�׵�����]?�e	V1{��^���"�K�˒�y%�^��x����Эi/�m���!y���`�S����Q����N�1? �+K�d}��S��{��XQo���6��HY�Oc�'m�T��Oҭ.���"����0�n�fϑr%d�v5[~�1�)�t�]�;�[3��*���s �q�1��9A�b�����=�O��� ��n�pK�Pc�D��UP��JL�{ʮLIҞ�u� ec'�$�U�;�'Zp��REv�J[;�_/j�>h;�Ν��?��B�_b��̥E .N	=��t!Od�����H޻)_&v�I�%�ҷ��H[�k��gZOP��Nbn� FJ���zz��b���.d�9{?�`�!�7�q���&\�<�t��$ӷ|n�\9��.���L���rk���E6@��?�`у��-A�"�>+�<B�k^�W����oE�Y�~��j���

#�j�D��g��0R�����3��r{X���H�����~u�"���! ⏢����bq�b�:��oE�x{�ҹ���n�[&�d�u�Kn{I��i7�Rv}���^����\Y&��	FFv���o4���Ҫ�7��󖀩�\M��V<�]E����}�؎��Te�$��d����	f�D��w f%f�Kv�A����yZ�B	dKȭ�{�K6�ۃ�=N|��U��9���p �HU˺r��WSE*c����R"=4.}F���K���s��ѵV��Sk5�4�͗t�.U��Rn�A�ÿ��X���h-�������s����7`��b��1��2oΡL�*Q���|������+ѻ��UH	�ؗ�XU�k��p9����T�%�yy��V�%�~)�r+^x����q��|�������J���*��x�Ra�
)|��uE�W���#hO1��K׍�Kk���2�A�p��u�
���r���@۬���E��kvX��0߼�n#�}��#���G�nx���2C��'D^Rtt�`����'^�~�-�R��-/�M9i]��|���n��W�Y����C��(G6�%/�$h/����M��'�Y/VE=BGb���@��w���ǆ�\����
q����o��,�B5�K���>]a���X�^�^���;nV'��1MF�0L�(;�j��b���Œx���_�Ԃ�����P}�!��e�z1�eɘ�I� R0�ɘ�NPl���MOh�ߣ8D��^�Z>�/6�[�Ud�3�Ge���R%�"�Ea ���c&��M��INz�.ti<8��7��
,0`n0}*SA�Ӟ��9�+�]�rP��� �B�D���������/׷rL����B�=Ρ�Q�t��!�aEͼKKm4����1�J�*ܴ�*j��vUm��N}�v�ϴ�����si�neC��Wl~��2�������]��Vh�ܦ�́�֍�
���8�5�w��$|�p�`9���L3"��N�E6��9���̀P�����~�A{{b��?�8��f���Q����n�֗���.��'n�r\?�vl+f�|�u��y�G$�{+�Qv�o�8�w���H/��&�����kY� �J�ˌ��'Fn�Jn���f@�СwxJ=�o��뇦}�|�K~AJ/X;ݰ;L�W]U7�;����������t�+jsƣ���";is�-�@Uv1y��x&¤Vp�C�e6Fad�ac/`��g�q�j)m�m��[qrI�	��yWJ��qg[�O��7��,�m��_Zݤ;ܼcp�8�*R�T��-_�F�5�(�{l�|'�~�}�p�.��o�%6w;���zk��/꛳:ۦ�z�І4�E���|r:�A0�qp��܌S�Q��9�Н�::t޼[ل�J��X�m���A��ہI?rCB"з���� }�SQ���7й>a�Q���7����ݜ<5k��W����9GPQp�n�:�j
�c�LtPl�wx�P�T@C��������f���.I��{GŞ�����W���)��т+w��	�@��Sa�`�Ŗ�6��hݙ�&se�,�c����h�5p_8]�aA�)�� ��4c#ˡ�η0�J�{F*[�\��V�ؐ�$Β���.���������!���Ŷ����5����(U�t�'U&aQ�P��q�%/�jc鼾0��DU������P��")���S'_{a��m$�`qWt/�#̊n�.*�����D�Ɂx|��-A�7� ��_0�k nf3�B@,o8b׋0֋d�W�l���C��S7�%��E�ʛD���M����v�����`&9ED A�E��-����m?C��\�Q��c0So�gAt��g( ��>vU4F��%�dg�)/:u���opO��6�̩�t�?0Y����	;��s����J���et(���P�-�`��d�ǁ�a�Eǩ����/��2���?Ú���ioՏ-k�8�{��ٜ��½�4E�,��JA�����e�'�Z��ȹ����H�^5߽vʸP4�rQ���k��?p?0�)#M]c}v�8���8?��o���&�66����?:�w�4�2�f�r�b���e�V�p�n��Am��� i�01e(`ι%L�]]lD�5�;0��ql^���u���Q��j��+b)���vZ�.��`�H�]G2��P���%�3�-�k'H�x�'B[1�+�;J�f�KS��>~vL�BK�9��řhK�Q>"d�ƅ�?���D�`�	����I��ض���5jv��
�����B~Z��e����"t��Eٷ���6N�����M���I�o��C��i%��;���(�DH��t�l���ܭ:�E��f���@]N�0��'59����p���͂��р�9����/�)A/�]�fj� ܵ�#y��Jމ�i�5�^睠�(k��1�"�FJ:@�a"�N\L"���+��Io4���P0�qĐ�R� ��\~9�|T:#ۮ���L� r��H~�D����7^!v ;�����J|;Vk��MQ�ڌc}s*,�o
�'urD����.m/�t0^��9�g�6����2öf��O&y��Qa	IQ����%W��|�P����N�7{ZjP�dV����|�"��r�(����>=h5Q@�گ�{S�D?`Q��Ҳ7�o?|x�E�����1����7���)Hre��,,��r��&q���e��E;����<@#�_pC=��4+���N�i�1X��7���R�h�F�- 3=�pB�&�Poi�↍�G��M�(W�Ջ�d�P/�\�eBԄ����ϓtz�ͧ��3x�D���G���&�X�L8�ĜP�J�3Q�	���*�S�"폾��k�R���~9�c�}@��Wp��k�O�e��	YwC)5�l?w�_�qJut��^�H4�_�?v@�8 ��i1�;���N�-�6�wV��4%��E��2�r��v�8�E��؃�|o���U�.�}CR.E�X�*�B؋B��^ <b�P��`Ѧ��������~J�ҁ��d1�r���/Y���k"!N�5�V���]4w]N�´�D�5r��,8�Yu0ϿP�x�����+���a�fo㺿��	g�o�#E^�9�Ul��~/�Y����k�����	��や���DJNh��J� �q�M�=�հ Gb�&��)��r=�QP8�9�U�\Q��RwQz��蹚�\�%���Y���c�nԤ�7�͂P�Q��G2���`Y�������w�{�E�I������I���Űs�C��;P�>��/�̉���L���6VȘ9o��J!�I��p39-��}��ߛ�%�I^�V_��
�(��+�����\Ѽ(|��7J}ˀ�p��K|cd"��n)���	{w$�������j.n$�q�9�^3V�a�2T�R~kk����9Ex���N�I7�JA�K�Ό�\^��h>�[��=��Z
�#I�Ψ���7��v�a�;T�30nS-<2;�Y8w�b3������!����#������-�^�!����p3���ym��RS_f��͊:N�y5xL'�E�)��JY)��=��LF�K2L�̓�ԈŃ�t�fv���-�9��b�2\����h4	Ř�}|�z ��3Y(�1�d��`������(|�/N����k�NF����c��_�vW]4�76���%A��N� ����jEc����(��ׅMZ��^�_E۲���{���ӫ}0\L�W�>g��y�;ze�J9np��k������P���>�~
h�<w��b�o�����B�i�`�]L���m��D��o��3��rTZش��2����ξ�0�3��gZ	�����1�\,rL���d�dQ�cgÉ�od*��=L����ѓ��'1(����c�<V=V�-�vb�n�J
��ؖ]Z!�g�[ci(��[o~HI����ֲ�'��Г��4�#��O��e�,U&��ٰ�u�%塇'}�;��9�[���Dq�*�����^d�c˖ά ���2"߭LT�*6E�ԭt��
� ��w%֞�8���������]{�
W��z;ʟz�-���ੳ�ɫ$�d��P����CYO/P�X���#��3�jT�k�GGo7�7<�).ń�=��T�,�~0��;�cU��*/F���Ej
�\Bw%1��L5��C ��FéoY2`B��l��{�W��V�І*���ܧ�6=!)d���$כ�_J���)v1�$h�o�;WV�w���e9�T�q:6L���z��v��D��e:9��b�H���ۡ�&���\gVY]�/����k�\2a��Z�Ѿ���0�iW�=A|=�5C6G����ZutW�پ��A��0G�
5�QB������Aa��J�f�m�ދ�ɍ�����/?�6���dVG�{�f}��uJ.�" �Iz�m��w�5�My �۔�`�l��/����N�dk�RB���1Ur{�*�$~ǟ����-������v��$k��2�Xp�S�D+z��;���P��w�Lo�mw�]�X�g�B����y�W�9[yr���z�G<�7=e���(H�� '�B9��=+�7��9��#ߖ� ƕm�?`(��!�'_��^.��Zxb����G�S����o8y+/R��q��w�=��-�R��CC1���򳭊��,�����F�*�jZ���</	x;U�7���W�>M����e,;���^�5Ug%ꊩ���%d*o�2�a+(��lU�2�iFvc���g�^�E��Y����Lfi�P�Z\��DY��������pہ�k�nȿ�#ը;yP'Å���ıGq�(� �h8Y&�(�G��i+=#�Éf�ϙ=�i�����P���6�\���Y�����yALQݵ��Ћ��WӔ��w��)D4�������!fM�8�On��]Ln$�.{DL�c�'��J�Ŷ��'X�AA-Nv˞#,,�>F��ժ�R�k(5j�7�w��$�p���p=��XV�s�i�
��d8������۪�a��>��eHU����&�.��{�u,W�g�R��P9���xJ�8��-�88���D+^�gF��%�ĭ˕���"���z�R>�(.��n�jg;�h�J����Bj�4���.:�b!҃`��w�i�K\T�a��m��G��},�����u����=N*��9�JT㋍:W4+�0SS-�KǑDx�����&R�涳�{S*a2��*n�*l�@��i�H�����SXӆ�8��.,���3�nm7��:����8㘫Mx�S�Es2:{�z�3�|�`
��j�;ZVق�Gv�ad�X$���m��osl�}�swߐ;�|3�Ԕ7L��b�ǀe>8�����9���c���;������DD����ה߆~Ml\?���&h��mC���hсH�;�+e3_ji,�2]W\�0 gnQBPT��(���:P�[bk�F�!T����вA'.X!��ݹJj�''~0e*-���,K�uFm�Q�]Z_�R�'h���+��8R�ֆ!�\ǘ��nA�u�`���%���I������_�E����8?�=w*B���v�g(a������9T���C�uo�	i����XU�r���] ����T���y.�2�yF3uo�������4�V��h��+�zt��{�0�z��������c����Ք��mX�9ړ(�NU�fF:��ͭ�U,Q���uT����������#�"�t����U�G�����"~b�CSdE��7��	�nn���J��~�m!OIO֞�Ȭ�Tu�}\�;\�?UǄ�����^%��O\3�c@Ȟt�C̪L4��Qs�|-/�%�0v�8��{q7��WzRn��a1\���DE_t��xՠ:�\_��:��4��C9���뉯��8gz�5�.��x�[��걥��1U���!e鍹p5�gײE����r�/�|���;Q9��*bL`-���@�l�.}�����C�-�Y�$e�uΉ^�y9��(�J����e�o��êJ.lYA^�_r钃����UN�k9ي:��Q��ޱliw?1�l�sN�jgt�޿ ��^Y>�����j�^ޔ�[��x�87�����aN��~\r�WbL(�&v{��Z�)H�h� �T<���Y�A����/0��){�(j1�	��(�����j`9�|_l�P�X0���P�*�S\Q*ҵ���3�i�C��Z��`�˒�dק����m��NE��aŎ��o���ȣC�K�G���}���pvq Q������?��si�v?�dI��4��ף�?�
5� �S�g������rmF^,.��b�h�s�0��~�,������� %���D�%=e:�M���qbv`���+����z�����٤�qP>3 �ޭx�uu��t )w��7q@�y�\�ZW4m�2��6�, �������o��� ���ibOh����H�x�3=�;\(ȳ�$y�9�坭<���ܻ���m�����ᰘ%/�����"�������kL�7�z�J*L�A�v�F���<=m<*���Ӡ<�ӏ���\��Ml-��y�J��$�*���8t�KL�j�Y����Qh6m�j��>g�F�\:p����_�4�b� �2]M�[�?=p�ad��Z�A���kc���	s��ⷧ>��4+|��{-:K.%Yn݄��Ƈ��S2{�x�r��8Uz&����?d����۰@�f�6��a�Y|�Κo��,���V! ���+F\ /��jD%��o����keӝ-��u=�>���ӖK�WK�ݞ��3���Tj',{!7hƆ7�a�Q�������~�m�3�����s���o^#콷 b\�(��1Ԣ�i��f(ƾS����l�j�S8�(Ԣ�����z��m���H)IL��;3���v�<(%�V�j���%n���9V��N�X&.�b���&)?����pE��p��4���5t�YI4By��q��՛C��4����Yf� 
���̮y�0�z���^4���P�vAg�Sk}�*'��3���J���ݧu��|��I�J�R �%v��nk��B����[�(�(J�����H��I�;��$8�����e��u\�]̇������ђ�%�˅���*G
sqޮ���!��*���~����2,�����a����^���.��
kF��u�&>I�B`��|��Q����f%U���(�B��J������ʟ=�� ���0����k���E�(�j�s�<���Hv&�,�kT�"����Q��#�{�.uȶ��Y�z���0�5�)�ɧ��.6�d NB��yE�@���:�=��OS�ob������Ġ���!��wf7���w�֋8�ߑ�e��q�^+�� 1z0��`6���w�N��W�g�0��IL���/�!X�5h�4MR"uT��`�La��?� (o�J�/r���1h
p5��N7��M����Ԑ����|���V�Z$��2K��UԪ��s�ᚶ=��Qؓ�w~4+Y!Q3�d��'��5)�L�$t6&̾t/)��{��S����<D9��M='�x��aQ0������p����a:�"����������/&��|�~���&K`<�_�5r�yj���}�CP�2-�j(��8�Ηuf�q4�1����H�ad�~HÝ���#(��.[��~rm�I�9��W_�����)���5;��6��p\�r`L�͍5�ѹc��x��5"X`6t����ྚ�
���`���-q���G;3�LJ�}�\I?�J�m4q���V�djb�G�Ǩ�N��3�%��ȓ]���IfH��R��0��`��:��|;�f��3ߋ7=l�e��raeW�����i t�iåWз�t�z�� m��%� f�ʉN�d�l��Q�8�e��g�EN���z(�.�1= u��&D2w~M��@���mf�^낺�:Ng���j�S��@�1����:=����ؽ��eW`\8�1�O���̢b�w��~�16]��{ �C�lڲ�"�!��_Dg�ƅ��p��^U�s*f�՗%��&��sg��Z&�zf1��2�E��
�ܴ�"_���j�]���=�L���
���pl���pH3�2�:�>򌠭-G�RX����p]	LËT��b�H
w��v{�7��B��u۪�wtRq7�6d�X��_*��t����òuf�z*���Drg��+����#��PƜ�7����R*��J�$S��!�c�zny��ȣ4h�j�Ц�r�d5���T����6.>��p���ʏ��r�/$M_��YD�$�a�|$�t�8������-x�o��M��xTz�0�g�bb�O�a(���!�^ϋ!���/�4�͎v����D���m��<�#��톦�R���@(6C7�y>���^$�E-A�A%��h C�<&�e�����]|�S�:*ܳ��V��(��iƠ���g��뙣qdᬌ;Op@�Ʒ��S���Ҩ��y3�؋_�~�x�4Iع'$l�ؖ^�����c	f߬���\�V�L����������g�F|���P�ލ�r'��Ud? ��A?���,�S�D82�
͞�  ؟�/("T��|ᖞ!��c��4P�y}�X~���]���	0��'�'QJ�5Y��Ms��Bm@���|^+����@2G�����U
!X���#�8R݋a����>������[�� z�-|��Ϣ�	�����9�����X�PI���<�>g���Q$��^���!&u��(�{��f���c/L���ȅ3Wp�ͯ{�)��~���Knya�V����nu(e��K������ۢy��R�^RH�L�9�%O�Qs�E�3����_��eE+Yhy6GK�3�)��y�jȎ0��G���$Ǟa�`"����@%�B�T�a��wDr�\�(j� �Z���}��\v��N�o�a�_<&�|H�����Ρ��k�� �gҘ�L���c�-]����:Ρ��C7���
�/b�J��W8t�W�(��F�Ū 2�P�i��˜�13�Ƶ�8�2�ٯk�Ttgw��Z(��-ujBݶ5b:���]A�X3$ )�����N�=[}��l%P|�zq`�>{�����F�O)l̛�C"�޻j�ݺQWc�2P�}�N7Fd�|EUg"ԯ�������}U0�Q>�����q�q,���4��`	�p/D�0e.i�
=.��`���j��M՗�\lA,�O�' MGz�J����[!�N�F����d�o���@s�������<��)-����Iq���_ {B�D?E��5Ub���v�G��Hzh���עb���p��]�,���-"�'���A9�I%Z�<����bȌ�R\�A��a
� ��*m��"�z�u�Q>�j[I�%������l�� �D=o���2x<A8����9�����j����y����&=u�{Qn>�`q%|����.����n�`|0�1X�m1��n�2n,Es?K(q���j���!yqԅb���vZ�M�V.�Z=��ص�c��G��Wq�LW�;�=ԃN�[�k�? �ߖ���%� o2#|s�����:��Ֆfr�G��GR��>� �P:�g*�G��{v���D��~	Ë�G�����c�ѵ���v�D5�qO��%MJ`�X��UW��n�z~Eާ���x��w-l�k�V��g?���%7���[�x�\�j���Zu��?ȇ$�Ga�,X�;ɓo��^�g~s��$����o�z&T8jR� �QJ� �⇎Bugg�&�-r�Lme�ψ}����e�tɵ�$�c���ty0AkHs9���H5ӹLA9ʝV�ܿ8�p�����1���7ш����>�dt7T��1��|�3���=:���eR+�&�Y*%�N����5�m���ڧ�����u���<<���ZR������2RdW]<�ׂ�Isb��E�&Qp]����ɵrM�'2][#��O�L*�\�j��b�90(,2�H�3=��Xǎ��\�ET4��.زk�FJT��AR8�ō#�V8!*��c��&O��]ՠ���`-��U��އ���@�� $�HGZ��A4-I�WE*�� ka��2x��"�Hg7��.|��e��lى�;��uJ��:.5 C��\u�A�	��|.r} J�!�@�Z��.PCIYKO�%��Fl�~�R_"c��4$xN�Iˇ�d�xk��x�E$�;4e���%�������s�L���pj�\�1���"�_BBW�������穰Ȏv����@��Vpq-4s�,�t��@����VL�y��qB�*���(&�4�'�/=ی�;P���3�Obے�iʦe|���o2سc�x�����(#7�m� VN��O.V�/L#4��bNכ�I7t��Q�r�{�j�ww��=1�6��� �v�^�X�6:D���R5���H�����,��l��Y�͓�h<��6��5�s�R�66�B�Õ?���-�h?����T���ۅ���c����n3�̠�i4�d"%�V&r������of������mLi������R ���$��~�'�|ي�r�f�X�������#4@$��+���ޢ�X�w;껷��*�\_��T%��%�1�J�;��n2Z�ǲ �V�,����,�D�����8b���l%����2[J-)��o} x�b�Y�5��{�G �3�]�Q�&�k���V��w_�7���J��JK1j�&B-��Iaw�H��5N6�'$��%MU�i�VG`\��?N��[�K*O�>J��ůۍ��ˇEyqyù�@3�I�El��ۤV�����?�4J�ފ4�X]��}�g�Ŋ>S�Z���`��U'�Q�/ۢ��k�qV�H���#�%�J�A1��t��5^@��n�x����������=����� �K�����ł�Wz�j�݅����vj���O���-.+��v�ސ}X��#Թ�7p|�nr��x�(�-KfG�de�x(_�Wt)��R ��D)����?F�s3>Z0ZR��5�=P^�ˈ��-��=&lpS�,�{�tp4f�j�Q8�o�.�cS��/`�yѯR^!�	Z �Z�%J�������H���ujk����C^��>�WC0��a�x⧵���cɵVl���7�ç��8�r5�Q�Y$qx�����u�!���������6?v��XBIH�K(7�l��u��aࢗ�6hD%��x�($Ho�SX��$�u%��V�,v�o��3�WI�p;T*��ؘ9��}Ǐ�Pl��^�I}���}��s�M�&�!U� V���O�U2�8��H��KЀ�i�Lz%>����-l�,cP�M�o��H+O��޿�͑���Dp�6NF�%Io<��^�/wr��}�m��m}U�?����7�4Bq壺��� _oc��oHA�lQ�ګ��/ ��� ��������>�����=��'��wn�}qBwۼ���:�s���]rR�n���'���(�*^t]�3JȦ�zֱ~�q F`��_3o��,�K6���*X��m�6ȟF�RCt�K!�s�I��Yt����Q�O:� 5O�ҏq�~Z`�~���>=iU�)Z^���y4A��"A��.��;�!�Sϒ����7��-]]*�t�ȜN>�0W�GJ�^RJ��G��k5�����IV��T�����x��g���`����'~T��v�{ġ9|MEgg?U�����78=��D�br[���/h\��c�x����3/p�&��a��}ak��L�x��x�DF��߀�S2c������ĵGF��Vv2��5����'��,өx5Y�ij9I�����|��F���{d��-k���i�R��ғ]���?�!�co���\���ds�0���f+����ٺ���O+)��|�p�<�?�ݿڸڼ�s�/��1g�<��\�<��t�F�>@�ѩ�8��K�b7��T2�Ÿ��(��C1�]�_����Ŕw���O3m��T9^V�N�I�ݽ��t��*�Hpx�`/K��1���:n�W�9�6`��÷5�ѩ������D�^>��m�τ$�h��,���� @��3$3��}��+�(!����fn�7E�,Jt �`���(�ل1��t����C�c�E֐V��Iw��g�IW::3��M���� ��H1�l��s,8wfp��]0��V]����n�|�/� �c� ����~^��LWb��{�<����9�d?�� |U�S�*K.�(��PZ7��܄;�vR*��Ҩ�J�}ڮ��O��s��������v`9� F���S�����H�/`_��R�G�D�"7�Xi~��Y�}�Zs��ǥ��q'`]4I"�T�v�p}Fi�'r���C ��Ad�8��/K�l O���!�r�l����������9&>�1e��=TP�D�Q���eH�������dL'��8���I��K��vEn���:��ظ����h���b:��.��1���
�"�<��H��������\F�b5z�ٖ�\�!t4m�*�&����p��\�hh�c�|%p��Ua�?�P:��gD1�X�l͐
/n���?6�ę���]^LU�',r|�K�XA)=0�`��S�2����
!d/��	p��A+�Lc�B�U�$��i��G��T-B���mK���'�t��S~C�'�CG�Ă��L�"���@R1��R�}xCesQ�h�~�Iju��(��O���%N���2$�K��Y������jP�jW�W4��t����_�_��٬	voc���"\D]��9k^�gm�\F�����f�$����`�Ҹ#(��'�>�/fQ✯�_ļ�a���6=���@P��LAK<�׬%
a��}q�Q�g�ź�~/�\.����ϯB�/�-a`gZ��;KtӋ���&f���d�yb��D��^�#���d�Z��X@��E�C�O����=$�mG��W���bHL��$�O��VTN\�̓�81�
���C�`~ا?
�L�3�4ة�G҅<8'<O����CH �U��R|��,��I�`�����·ǔSz[���ю���Aʯ���w�!O��#�����I)ݧ�3p}`Y��h�B��hzW���T!.>q��?ީ�⊧S�����1k��!��1�� �dn���&�+�/��44R�A��$����S5,�V.���_=� d!'d�괼�՞�� #����VJ�WKi4��h��Q�W�X��U��`�����]C���D��ץy�U4yv=���2L�t�����",,G?�������RR
WB׊+|k��Ϫ*dG��2I�h�QN�?Enh�9#���\b{�R�/
o�i�a�Ja��{��O}�]F���Sdq��D�f3�v�7��+�}�7t�WCǊ��ю�:��|�a����L�=��D�z��a��͛�N$��m#�|��t�rmeph~D��L�������\�FbN ��^r���_�tEGro��0O[�e2���4��}�߹�z �1 ,�J���\�X��Z�{Vy��W���Q�����
=���׏�����a+�_P��u�:�xe��TS9c���	$xQ�}�R`^+Q�GM���=c����E��z�я�Є���c��|+�q�UƘ��9���W��`P���*��U�����G�TA��t��&�	O�k�r/WZ���`��:f^7�L�2���]�My�x�cj��<��U��u4�tf�|��1���(=��?�����?KO]�,8��yù⛶���B(���0q���"fv�?ڼ��ZH�B\����]��Z���������=ЂY������J	Zl����
3���y��	N<W���:�ʟ�4Vo�YZ�;��b��Y��0�]�+Xm5���2�G�e%��0d�|��(6�>w����m�N�rmdq�҅9�m�[�H[jT��I��Ĭ���Ar��L��+i\FQ+
j~>c�_(����l�G���	ܴƞ���1��~o��m�/�=����b���}���=l��'m�+lVEC��)�Re2l��=�m�۱��"��ύzm�!����ܐ��"�E�ӯđ���⭹��D���Y��5e!�b���b���OQB\ʿS��;2�Y�G��`���2��G6٬���қ�\�����0ړ������u�5��Wy:�j��:Bs����>�<�N{� �B�/8\�}{�*f7T�?�p7ױ�e���m�&��o�@@��^�
l�v��UP�p�C�
�#��c�Ln^�_Mg����1|����K��5!D9���o�{��Gd�LGM$��ٰ�z��)0�op!��b^:���m�}FDs�����t�B�{�)�[	��)֟Ջ�w�K(I�x��4�-4�6q���:�����(0��xdM.� OG�4`&��T���p^���Pڨ���������#�F`��A`�G{�C��/_u-a>����V���#P�04X�O��i�L��c�~�kД#7�3}]侫I����|)`N����l�&Fʫ$�����ٜ_�\�֬����Kΰ��t@m� А���\GK1�Sp�c�%�[�,#�T^���;(?)�d������4��e9��N ������� .kn=����uLxo�=��눴Ў��>rD�"LE��G���㠷*��Zj0�\jQOJ�|��;5h�m��7�"����v�����)DY�ŋ!��Rlhm|{����W`��2|���XV>���=r4�}�:�$�L��;5@�ȵ��&���,}�	�P�(���bV�2)}���w[���L�5
 O��e�����}�c�Ղ|���y��Y�s�:_N��,vg�S�4��l�ȭ�=4�{qf��1�&�"��SE8�ci!�!�J�V�C~�Pv6�y���G~c#8#5O�a�j	�]�R��Vj�::mZ��N����QO�G���n�8\_�*�v�#r��ܩ+mA���7�� �r��>SO��z%aд�Cq#�* Z#�Ֆ�>�8�u5F׊�S 8���z�?�A��0b�����`q�ݎ�Q�	�.��~�ٺ�(ѭ�z}!�B��<+����������ц5�a��������g�0�ɩ���u��B�H3㙾��������&���%pUԍ@4O	)?���A�@҆ն������QCI�_&�%��2� �9�v �و�`_�I�Pxr�D��{ι��re�~rn�TBM��m��҉п.:Bl�$�3�87�~g�����)0���f7*�c�4'� �ӿ��L�<�f���m�x޿��Q¼�CS2��./>����vT��C��[����/�ތ}�_QG�`�
��\���<���)�;N��Xd/������2|�� �5QNNT�k�� s��Q�[�ԃ���)}�F!����浞�ݝ^�\��52U�g�yE�"<�P=+h������ky}7�T*�_��\�Un�Ȣ���U1߸� �� B���6Y�����T����7#������?&/-2f)�c�%�m��h}��i����/^t�0Ҵ3B])��G�Z�i��m�cʡ��D���;�lq����E#��{E�>|�Kԋb&��a�IP��n	x�F-�Xݏ�BS��x0 ���]� �(e����[�z#��S_���|�̢g��������Ʉ��ۮ� ��N��wCű'�b3�Q� �O�>��ݳ�|q��ڨ��`��O�-H���2n����}�DJ����N�8��G��G>�>��\C�9�����&��v��꧋�W{���K"a�(#�[{H��+@h�/H�a�b�#�:�d�׹z��]i���?����b�̦���R��1�$�����I�srB'��$�g��<��Ѯ�r�Wbx%'�F/�[���}|H~��ȍ�)ǀ?�,٨�'4zB�՗{��Y��rѹ}0N�҆dL8�Xy�XEd\�u�P}F�d:FP=��ʧ%^�0��u�O$w!bW�ƀ��T�V��SBX�uQ@\����ф��-Ea!�d�ȇ؞m�t�"͂�0s���0���H���D�s�pWֆy�M��w䳈	�߱��^,����M@�p&O��������_���1�@��7�i���oL�����6�l��^zg���kB��H�;��wJ��&s�N�>P�b5�S�ʞe�o`�<BC����ߘ�?s�.��	R���T�����ljY�(@pu��D�e[-�.*����z9E��F��2ω�#=�����$�>���Z��0@𬿚-&�t��]U�^-b��9�e�17��J�F�k��l���C�;�٫���*��	��%��J�@POsU�n\��^�ya���)�^���A΢-�Ebm��6}�e���a�i�A�D^������8���|E�´(�q��	M�b�g;���"�뷶W ���"�b�xjN !��1��q���\�e��1t�q�zq{� ��((�P���<0l�+��Q���A~��ŢB�,0"���Z�����𿆉�4�f�3����Q@�0�`l*���.�4�Tn
|�?�˕Aj,w�12�i%63�J?�/��(�^�q��%�����a�
 ����`cq^�C* �ߘ&ʫ�vo�O�7�����$!fߢ�� ��h0��`���kZ��6������5���n�	h��t�t�B������_��V���P0�rGh�J�+8��e�����0�_6�e/ � Mi����|l�U�����o~�L}���`k���;�1p苕�1\+Z��~��.�u�F�<�U��{�B��")��#��8?WIG�����x4�JM	���� ��^����x-�E瓀x*n6����|�^Po8��N3�ǀ����F@h�VS�1��¥���jy�����w5"r��z��&�ưM�8v�_��\�Y���R���G0�D5JFh+���1�b����fT�^�\��٠����+�D|6c�ho�����^yB0���	�۱��)�&�b�g��#�x�a�>ک7eq����j{byE���9�O'�3 ��w��A��A�5�1Xm��<V�9m��^�f�����V��y������� ��X��o�A�c��͏#l@T��^�����u� �y�I� ��8�6H�gKYՉ[p���|�e�w�6�Q���)�����[�XlR��L$%���s���8������8�ܯM���U��o���kOw�"�u��&�1#���X$���\O������`L�,C^���0�
��ҳ�y\`
<�u��:MKD!tԸ%�	 %�=ˋS^�=䗧�~nd�܀n�R���?��?ɳ����\Y�I���<��{�m�8��$�>��$$J4����Q��8�,�Ȣ��C �(�_��8�����(��8�s�ϲ�-
*��ܧ�%�z�$a�o_���#���������qt�&�G���!dC�ӚZXmb�H��7	�ӛ1�>�^��0�m�J��j��3ŞY��,f5̷�|�e��.��MJ��6m
E��Պ?��A�-�&9#�Z��s���%��.�0���
*����hPLؽ�p���{��C�#��5Zx+Y���
4�7�A������%i�)�`!����ܠ�Lg�_}V��o{�-���e[����XCj�$#��8���>���u�qO���S�Xt�y�MB��_M�v�A!XZ��������V5^�D��p�W_K�y�5�
u�	yFa�R�>��x�P��s@���Fzlf���Vc=d�� Ц}�3�}{>���%�?�|�N���Б�W�Ȕ���j,G�C�F�P�����7R���)Z�cʈ�1�x�Ƨ{�x�C"p��	B��M�N��ڨe�9���L���o��󒻫��$Ӏ�JE��З�-#@c#�R���2�AY�5�(�:�LN�O���D� n'*t�]F`�@#Z��2���Y��$Z�}��B����3�EϘ�Т.����f� ɡ)YTcKFr��l�%&��5��Ώ�zJ�ٻ^�8Tf>��Ħ���e�?�Ԋ���>�����.a��d�u
��vx)�e �Vu�F/9���5u(��W��oTu�󲋯iA��������lߛ�٧4���b́X˵a�X�ĸ*I�P�#� ���q%��^�ƚ��W.�^���XӂP��I���C2j��f!a5&����}��X�7�O���鼉�1�q� ��-�U�Q\�[_c+�9�L���RM[�q[��}�C�y�ug�K���R��x���T��.7�R�� }�O,�n�?���������)��_�]������*�w�g�d�D��bg�NiqU�� ���!�����8����As'à��)D�^
�-�ūV�[njej�q*=�9���'K_`y٫���V�ſPy�}��b�S�+E��7��k��m��Kݩ0�P��j���&^��Q�s�����G�9���'y�kh.ʑ	�or�c�ʠ`���W�d׏����E��t���t�̺�	�Jot���;ǫ��Tv~&�����i�����W��� ��!Z6���%nC��y�b��v�@_#A���N6�<��Λ�]�W��閣�����<��i��[�0Ӓ�kĆlε��G����NG7.��r�G�뿪�`3x�������:(N�G��¹l��-����`%<_B���k�]�6�BG%!�)����៴�?䏬n��:p	���ij���nw4V��KW��n��1��"b���F�eo0���Y]�<oB�V�%��@�P�Qx^n�h*�u�hO��Ե[G�Ͳ�4��`%L�/���Gq4|���:�%t�2e����1B/Ҝb�30X�1Ņ�W��a\���s���-�W�^�`�����i�A����l}5����[7ߴ'�RM�� Ԩڦm{�K�� X�; +�|�ãY<,e9|eq�l��/(n�Ooj�gY~H�m����x��6�,0��]�@2�lto!��u$�������u݃��{�
��U���
�-'hn�L���Ӄ{��O����[��qR\�-���r��aLC�o~uB�p,�o,LQ>�$J�u�xzSQ��73aJ>�������>������(X'�
g��VvV�J["�冚e�7�o�Zn��ÿ�z��H;�c-my�����,��x�t��˲�	2T^�rB���+�����44�,Q�F����^1c�H0(|>GI�����b1R'c?}�]�����j��xjr���6��D�_(7�T�O�-meu��s4	A���O��ߠ��8��HК�D+�e	��^�\�ɜe�R�A��� BY��L֍%!j�t��frS�CaY�A5�6���Ӌ��?�5��%7���<�҉$������Ȉ��`Y9� ���WXi;�p}3��� �T���2.��<���Q���{�p�&���jZ�տ��S/���r���,�C۵��a&(�S�V.�1���7�`M�Րl-��a�y�������vΧ�ܔ,�N��L\�b	yB7(����3��p�VlgA~eq�a�7?p1��ѣ�#�C3\�n�/�Xf'� I�X�|�r��49C��r��C��6I��R��".�x�Ih��5�m]А����@�Q�M��&C��L� ���{`����qk2h�q��]�8��ݮ���P�^�䑝�5����O��p��k��;����&�� �:`�kq7�?1�&��V/��S�3���(�q�7U�Q��V�|�6'Y��&!��*��j�ˀG'�#��+:�Ӹ�Pbҭ1�����ޛ?dƔ��s��O䵔	3��J�FǇ�O�>�J���W���hkL���V�G\h#� w�+�c��|���'`�-ɵ����D��9�����$4�+�-x�v>�R&m���+ǟy6��M^�U2��`��KnG,�ߘh�b�ї{,��]������^����%:�9O��Ue��}�J�UMٯ�-�_ɛ2�\� D����^�DU�[���Ԝv2;ݖ|c)V�ܔ_k&�*�^ۧ%�/VC����h��ޭ:��[����2����2�!PÑ���f���Ȓ�<(T]}P�P�\V�tQ��9���Ap1gM{�T��F�A�7��g@��W�i
�V�,����}�Q�}l$_��wԆP��e�+%����H�Um㺼��E�Z��1}o襕ﶪ�2���Pʸ�Lߦ60����ZW'J����Eo��������X5�(��`R]_��V�� >#<�-����r��;$
�w�V/'W}7cÇ a]�����g�NѰܰd{���*�7�X����i�x��jW$��������Y1�#�x�I�������rܤ;c�� \U� ��S���O<����n׈�������������	y�H�'�D7�3o��6�ҥ�5�$�s�?RTg���-�"�aZ�xk�z6ξ'+���7��qGt�k�/d9�'P�?����e-8A!UK̨��� Tg.�s���&x���g-���J�"��n�ʤ����]�sٌ���<��l*k���s��������ם�#���=U?��' �O����a��[�F�J2��[ZԢG�_&�fO��e���QN0Upq��Ez?�����e����l{�,���� �a��`9��i�-�<;rZh~V]2�v���8��$��{-eQ���i+'eí�>�_��#�!�����>�$�"��M�̌w��AQ�|}Ş7���ѝ ���?E:q &c����_�R$�	���z"c�0����Eo/8��&�ݟs��pNHC=�1������t�h��̩����~F~Ok�5$M�k1��r`��h�=5�P�z�q?�Z�[�8��u�
�M3'�Z`!��a�hpٽL$.�➜ːF-�����y?N��;��t2�_g���Y%mn��X���Ks�刯�
3��t����o�V���������~����&�m�r�H�PT��O�Y����%� x�>rS�pE�����-�[��#z�K�O߀��F#��=��O�-��+/Zq묍�d�0�3z2�
�01*?���_�&��֒	b7�yRYTx-���\/�%9id���#K��
��e?�����'��j�&�v�@���D'"���+�=l�L�j�o���#�3[���}�˥(D/� �8=��O�?"��z�e�66�ۆϜ�Nʲ�Z���8��4Y�ȉK�;�)��W\TQ�p7ӟ��9���n%X[|�+:n�.�3����5���>�!)Mq��"s��d�+�O�6X�G˭߲/��E��A;�����������&�")��
���"1�#�	�h�t���ʕ��s]h�;ॆ��,��Ƙ�? ��+�UPs���{ꣅˎY��������JNu�yN�fWB���%׺��2m�T����2d��|���LfT��>dy�>aw���X���F!��6 ��\������t��d�/���n��c�wēDS7�Q9DFQ����`e�ӿ��ݽ$y���V��; �8yp??���G*��z��)�)�R�}~��oY7�4���i��h�߼��$8��Z�z:=^����3�9<&��8�;�I��9�W��	�"�z���4�B�L01���;gnp.3t�� �"I�F���f�X�͘��N<Z���=CN,�zcՈN�^�	Nr��e)2�#���j-���jmK¹�Ձ�8�&�Px�k(��~x{�6���Z`�#�&ݳ�Q��_>lۂ^�2W�9끸Ċ�32H�Ŏs��ÿ�е��X�6���7�e'.�Ź�:��Cة��t$�q��q��N�=������n��!��'E��{�y�
"Y'�N����w��������ɜkD����^3�S������vÓ��Vg���F��D��2*�\�z�kG�&y�����zx�tIv�Pv��2d��0F��rƸ�7�
��[��M��,I�Z2����"'2���X�Sj��}�����QNlrc'�M�O�l�A�Ց�m
����qPV��l������F�͸��~ճ"������J�{ޔi��]�zj�f�P�2n�b��;�s�_�U�� ?c�_Bdm�a]�1D�:q}�Sz�,P ��oH8Y^_�#��&9�jm��v3S&P&�r09�X,�%O��'s$0n��yd���].������bl�<��� ��Tqj���_�U?��p'oj��WrA�i^�g2���c*<<W���I���؈�W�o|����\j(=o�p!�O�39ސ����]�|�U"=�PO!��{
��X�!nR<w�\�(O����<�~Ai���0F0�ث���R�|���0gޫ�����H{wt<�sQ�7֫�"��H�?�rJ��'�-�&.��f��OP(�:ǣ�ͻf�33�0/�9 ���C�g�m�����\�Bʷ�;Z�3�j������tB�(�������"��)P|�4�o���/��J�"�$�\��!�Ӿ��i�����n�\G�y��� ���t4�a��>��o��덋�U�Q�mڔ'q�`D�9���-*��a�S"�x�w;�i.�Fs٥tV��KS��ǲM_��xqrE������h0Fml��`��JJ�8%�F�K�89M�ց�r�����hg!3y|<����A����ÛIc*g�I/s��/�7����:D#���BU�� W��$�*CFT��=�4��P��[�sȲ}��82�&+�!S��i���\PcCޡH������瘩����w��x�-Y���l{c��|9�����FG�e:������aw����~��+ĆT���%�.�j �S{C�̻z�tJm�#P��%~�oՙd��&���~����M�R��H64EC���IW$$�"�����lmQէ�e�|�D����8��^�4c�#��"$���6u^� ��-�����O
�s��t^�h��\B��覠i]��MG'��7�"̱G��7�)��ķ���Ѡ�P4d��.B M޹���_V>���9-�s�^�,�x7�BȀ`�w��gL:"c?GWa�����z�'��Y������ɡ��ִ�l�y��d�w���9���}'�����}c�<�����4/��'k�`h�����W�$����#$���x·Ƽ���9��޶jd��`Fq���;�σ�M��E"JNT̅���+Dm�xd��' 1��ǫ��(�
^5T���%��Kv���@�jx���Q�L7����0j�����Y��7�Z���i������楋��i�R!����|o����qTE@	��	^��!"	w�xuEb����O
�Wv�S�p�87ø0\�IF����r
Y7�M�J���*��[vz�>+=�]"��w�c�EC��{ W��Iq������J��b�;I�͡W�e�`�/�������b[��`VueT���'����N�3>N\zY������o�36
N�Ēӯm���A�B\KGn5ty�TI�9�à�i8��g�&��y����ul.���Z>_�G^P��4��N�6U�#Y��������F�ez���@��ڛ܄.+�@h��$��4[[$$���_���0�p�
�dUgm���T��� ���]��]�)f��#�H��3j>���o����n@���"��4��0[�A��Z��P!��j)�:�����)t�n`q�h���Ž��V��Ưu��z �"�����./T_1��@a�i?�]r-i�}����sKCZ}�3�0x����W��`�v�メhR닀23�ó�-G�.+����	�X"E]�{W�h�E!��m���_���ΠT
_[N�L�xN�(�U�G�mc�˖j��x��a�����`u�9Yv�5����Itטp�o��J��v�YO{���[�s{�5y���ηo�n��������T��ΐ���"�
��qa��
f
�t����9�P��*T;`�B�`���͘-��j�%��|�eX�RxE]Lp H=\��a�F(r9r�CPb<�G8�}2���j�F�,%�5𷦍����<isU����aHaŒ��bx��r�O�5�_�PoS���%�V(T.�1�x�0�ؗ�}m�,�\:�oӢ�A�z��7%�[Mz�,�:�C����v륪�4�LUw��s�e�?�&)Pu���z�n/p����B`�S����.*$���D�-�_�l��雌7J< �.��Hj<#E3w,��pFg|�w�� \�y+4��čַ��eb?��1�H����8�J��y������W���3?}����|��ռΗ�D4�1�����*�ߚ[�v�{z���
%����~|&�n���V�Ͻ��R�ڶ���Ȑ3T���*3rƳR;�R��N���S�X��ʼų�ȧB�_ŉ����ąl����Ǚ�lV(F]b�I�:�6aJ#-���\-$r��'�46�-h����'�[�7�P��Y����+�PT�ĉW�o�H�5�~��~�=����ۦ�U��wj�iu~�$��\4q��%��Bh$��a����Cm��:y�w�7�����%�!_@Y����vn0�)�h��ҭ��Y�8���ޮDM��3��SIn�����Iʝ"O�$�|U,wV��}и�q��l$;�����:]WT�w'!ޮ�V~l����V�w+�ҽ�Jd���n�_��Է)�PM�s�������^��go�ʖ�� 9ۢ�>}`a�p8ƣ�f��)��J1}��rSi�>YJ���I��F+��nfl�\���k0Ղm`a꒫!c��,CqI�ri�7�J��i~�����n����wtC";N角��#���'�8 d�I�z�^e\oܒ��g���Cq��y�2ϼՂ�ﯫĀ�Q�7V6I�}���
bȵ���۸&S+�ɛ� cR��`��U�K��监� ���x����k��q����&/���A�6+�7��fK�A�<7����5%��@xK8���ꈔω~�T�34����b ���l�|���q�pY��8���i�3�D�υ��&�p���;�`u�i��Ei���v]��o�_Y��=��.l�1`+�Y�4��(�*����0C����W8���a�����Ve5u*�><���	�� ~|J��G���U/`�HٱΕ!{������^�*P�µ��"�/]��
:��}&�[�iR���)4�M��U
է���u]�Q�F��OLѧ"h4�a�^]��]���Tv�jIa�Z�?F��Щ�Ƥ��nNcex^Ts�{����?gIj���⚣���ZN�ƹ�;��������TY�3 ���