��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|8���e5�I��d8<��1h��}���:z��n�Z@�8B�:+%��Hx<2r�����OuT�m{�I@Yr��RB���*(�!����:|�wB(�{>�3h��nR�܍.�V���_1
iP(?(&êI���y/+S�u�b}���?W����X�\�d�l��<�&��M�I���_��؃g��9�k����b��uBh�ДI>��72-��/,��AR�bO���p���A�^|����C�SQy��%u���H �,^����5�^���IX��OO�4
5aK�Mʙ�cf*���0��9V|!��KR����"���r���P*��l�;Dau��d��4?ހ��D�:ų5n���k�u(�x�;N�~
;��;YKE-�݃�Qz���������Т%Z��Ȧ�q�_D�z;�Ə�Q�w�[ߧ$�=�x$���oՇ̱�I�)��� ��"��ev�!�Mr�{�;-(�-7`K����P�[Փb��c���L��-]���,�W�T��9������pB��-�"��ژ?ŕ���]k{J=e��
*+���w\���8�Lv_�b�s���!�Î 
Lܐ���h�Kop=kI�t���#HK����/V�4i`~�T7J��� �\��q���]c�V4a͓0�9�8� c���?�"d��7�6j��7�B��[�{��֍μ�uV��S`^m_�Pk��<{���3�c����+��/�O7�L�����#��R�n%�Bb���n��2.V�x�f�,k4ƨ��7�Ӟ�+č�|S�M�iglvY�p�$9�2�kCq�s�7R����K�c� Ĕ�Ë%�K��v�wg�x�,�Z�V|))������_����iv��<:Ɠ��yt�p�؈ھ�Ȧw�kC>N��'x�#@�`e�v4NҀ�N���]�
�޽o2��x��G��N/�jdo���|i�&�sj��2���n�}ޛ�>��x���A��bC_�Ȱ�=��	���}�5-�������r�3Ħ�z���!s����\�{��q��hz�i��y��=�PQ�a�H�Լ/-�}EI05:�P�1�6�H�՘������Y~�&n�Ӧo����[�V틢{S�]�ߛ0EK%�=�����ʕ�ű����3")��h�Ȩj�7�&��%�lr>n})}h�v �˺���H�r�H[�1��X�Am�]n@����OQ������Ώv��C��n�H[+V�؏s�-����z���EK�]�C�	��`>#4S����+���p������gW�\�)�`���
!����i��FJFĘ���\��eI��cW^:�s�%�K���?��ƻ��/B\.-�@�Z����]���P{vd>-1�-P�S ���
iE�#�,s#3��#�'����~W�Ξ�����
��_� �k<>�K�)�ƅ���fu��)[p�୭�Rꯇ=S_�,:a3Q���>�(����K){�r�j��%�r��T�ג������q���q�钴|�`M��_R��^�.6����
_@�'��ۯ 3���D�%:ݯ�IT�Oxs�����3�)"����ΓV!����Zi�Tt�O���I�ۯd�)�A2t����uΗ\���WF�hɖ� ���X�Td�<
MGf�4E'��=}"����\��u��𘱴>�uVje�AqH^|�=������g�0\`�pUv�^�6!ٛ�����=q���Jr�m:�hn-e0�e�"�s �>[x�jԀ�6E2^��0��!f��M���`�IBH��+����d9W��s���-��	���kr0V����u�V����-q'���1:�`�*e�y����E���!��k�X������\�9��s��b�c Ʉ��#4�&�9%�/�ٗT�0���D
X��j���m���78�^��X����d����uZ@5�X~s+�����:aL"����<��;���?Ǖ���1:��PF�-�!}rd+/Q�)q�(��}7�e���A2��@�w N=a�ȡ�I}O�q]<q���܉����PD��M�i�φ>��[06���T�Z��5}�5l��4gel��"qI2g(djI�
��s��Y�Nі�����BS]d���H4�s���9���җ��{]VC�ک�+����� Fݎ����j�n��@힇'� �#��oa)��@re���x�Ln^���ңB'='FZ�o�i��d�x�������H��ދx��@�C �Y�90���*:ϴ�m�{��.Pg�~�_H<�/S����뻫O1�L��/����#;B��oTn��56��n�"y.���=�J�N���p����	�eDcoYd ��Fg&��T� �����V�Rf�:��2tt�0�{��S?��ʉ~�K��v��1y��ذ^#W�d�}�������^>,Gaf�MJ�D��JvnW��f���?�:LH����zf��P�6����4��R�{O`̠���,���CJFݹ�.�G���v=��z���z���m&������L�r�_&�-�d�{Hs�h��Z��6�5B��#�.�ޠx�4�B����:�,;J��>�:�ɕo,�ƒ����9��i%,�P柝���q����4Y�R_%W	����F+N~U����F�/��T��=Am��A�0TC����#�h骿��ld,�<��y�Ӏ�"NyK���^Z�!)�����΍-��H���SQ��R4*:�U���fa�x�9u�n��;��U�<�b����(_¨k����JxZ��S2�)! ��{s�b�×
��ۨ��gLJ�2T�H�<[�j�R@�����w��:o8����P���/��_��8��\3bXx��qd!G�����q�<�B����6��J���F�;f:M2�ڞ�Ԯ����S����"�T��%㙇�¶�n<�Go�Mq����7��K.���)iKA�v�<S��c�>����$=9lk�� `�&�/$ك�j�x�H��T�r^x�����������띦�g�][S�b0U�Cd���ȥ"��:b]�=�}�5��ŢY��"p��=��w52Eq�E��d�s�>�A�k���A:e� i�T��=�G8�����PH��m\�Iq�'���@��� �>Nް-�3*$�-p	">o��6�+<]�afڡA����:�K�vkB�Ŏ��nܹ��)�$f���l�Cd'&��\��(��%�C��ĲA���>���{yʛ��z{@V=�(��f�$-��=��.o�h�n�� wֲ�P�9��MT��LyNd���r�0MҞ�fq��:��i����[����G�M����l����2U��r2�Ŕy�ӔΑ.��5*�T���q�����W����n2�����l+BJ��I�\��a��%�p:t5�˹�mC�e2���u��沽rRR5zf^��ޚ��s0��-�§$X�}�N{TX}���҅�f�9.�~��.;Ќ=�B@�v�o3n��W�ak!�r�u�N��Y�w��d��3.��X5�16[�����¢n:F�h�妢�ƴD·<��$��k��q��<~{YA�!�v��e�r)�k�Q�	U���H?l.�4��vI��ˏm�r���:�%&���1-�$��M�!�`��
q"�{���I��G��f�mCN"+(���������
�6u-�.�,įɭ�'$�غ��ROm�p��X��pp�H�4��D�bt���s+���	jd��Q�t`�!�I�YY���4���'N���l�˶��Hm0Z^���U�OE�ᬗ/�T��n�B�zSQ ��~hI��gTp���K*[�蚭ÈIHXQA�Ll2����.�yU#Y>����H��XQ5YH���rے�V���޻���G��f�2{귖���FtE�T��P�\>�n�!�;��9N����G{bk��,=�ڻ��~FJ�jgm�<J�1��:p��������h�ݷ�Q�sF#&�������f�֎��դ��B؏�������u��uD����_Y�ᢟ�ִ��Kq	�|R�	��(�>��"H�dvKf�c��:��f�a�ʌ7JԒ
����1܏ۋ��7�ؾ���1�
<��`�G�_�G������=]���ٹ�ʦ���P��:�zz��l�>�Q�<c��ua&����o�5�vȃTVs[%�9W�p��n�hp�!��<U<�����?6�ȜZ�_u���G�q��&�Suf���m�'F��6PbpN�	��\o0잕ƫ�ǜy7b#�e8���.�T�,y�_n�I�������Ћ1z���p�e�'��ڂ�u��N�qƺ�'�&�3!A�ز����H~� ��yɸ>�Is�cZ�BB��ĩ�;�>��������t�3��Q-T�)��R-�(D���,�(�.}��h{��9*�i%�2<�����!S?ha�~H�s��ILg  ���{��q��pꑧ�`SD�]+���i{��Nf��Y7�5�͉k�>��b%��g<�����臉�=n[��01*o ��@S��x\��|�^+�w��7%��s�D�b�s���}��J�0�^P�������hba��8W]8%�~����,GmY$�̥Ig�yX�۔��A;��������¨c)�4��<.`{-��y�ya[8})�P�h���@��<���s�+
Q;�ZX��2�*k�!1Y�Ov�e{� r�P	`�i�b��h�w����1��6�an"�����5� e��p#��ダ�|�c� 2�@���P�v�,o�\O7����B̿��C��)�h��q��l>؋қ�K��ڊ�0xe�uɽ'��p�-}l��,� I�x��J���'f�vG��R��=�rM߻e�3�_��ؑo���#�������_A,��� ��(��������kd	
�y:��yQ�^'���|甹���Q�c?�XN����%�(�`V?��w��
Ӿ��Y%��H��s����,G�7{JpAr��D������H[���j���0�g�(�8���w$yS��S��B+AS�9�a�nL��P��F�66�r �W��O�LP�����5�R���w��%?���$���@31�pb�\ Ӱ%:�U��T��x�p!$���E�%����,����2ϒ>�c[�Y�4�P�&m(^�K���ͪ��,���th�:a��b9����[��]˟z���S#�ܲIu|r���鰖[��H��/���n��&c��9�"�>ʽ�t��)Tv�[>6�w����m�y�r�ܜ�D������l�S����KjcZ��;��]4G��.���,K�X7��	$#�Al��Q�,��Lڧ߂���-

��v�d�H�1a�ca�(QO�tY�� �o���c-_ɾ���P�ٔtm �L��>�1s�@���o���o1��h��S��R��wL�D��^�Lf����N��K/+�?�; !RA�G%
�h���!66�ݚ_�SVEOh����-���\�j��۸��0|HH����	�o:�b�
*��f��0i�
�!����a	s��Nzu<�H�2��TN%�<�1/�%0����9DWO�"�Y��´�|J{���w����}	�k⟾��b�R����0�8�������f��,��V [Zٮ3D���"��'�9����z�\�r��n���a8�'i�ٕ7;��G��09�Wr�Ҭ�QS���o�&��bv!�����T��^�X/�a6�gT�40t	��RL��i}�`Yԕ��L_���m|Yb}��j��'��蓤R-���86[��v���/ʴʧ,�VJ)�H> D�\]�9)�!�nH5
߸�zN�h��
o��c�t��P#h�jK���-�ش��H�;ſ���[�BJ��i����i���OF��D��aeB3��+�0xx�2G~���k88a�Ge�D67G�K�sB���Ҥ�+����LA\��{UmgS�K/�!zS��qk�8˴��[�42�f`_�q_3�c�F���B'�+�.ָ�4ɟ���Ǝv�ov�s|'��RD��!=6������q�'���g�?��ˢf��w-^-N����7��"��sO�g*�`� h�L�8���V��Ξg�o*��d/d�:�22E`�/\H,�N��A#�#��C5����m:G�j����M��ȼ��%�
��8�w�2E�w *ý�aHp�� k���C�`�J].���c����o�	f,�9����I)�@�M�
��t����RN�q����r=�v#��m�ױ�ݺb�V�#��la5�=�Nr�g�� �i`4*c1>1w_�כY$��q�E2T*[����~W��WL�DQ�08��rG޴Wِ���g�i�ugLs���A�D��<�A�}��o!�t�P_k�[>�8ˑ:��V�#�J�J��>���в)QY�0�9��?\�&����������nBĹ!��ր�����8S�2k�%�v�J� cu��M���y8P�?�kE���,w;���Ya}ͧݖ��j��v�1�JuTd}3�f]I����_��6�_h���w������I��[������J���Kt<�4�'Ru�mCxͺ Eٸ-3�Į�?�$�~��R&+h˗vjH�F��6}���Un#�1��W�n��Nip�>�G���W�v" ����Ѷ
[3#&�����W��A��aN�'� (+�g3��F�KǦ���/56�o�smƄ^<�P|�
��C$�)]RȊ:��2i�X[�l!���0p��-%?��nד�W��>)r�
�4��)k%¯���]^8ٞs�a���a�`�*>�{[���:'��C+O��[�L�Ҵ{$4G���b;�导��W��"�����s*�"�L�8��&�
�>����[�C�`�z['��k�c�C��;JN�*�&�O1H�h���5=�����ۍ�!�
�H�V�.��!�¬�e&>��
�*�����.�:����.��"᭖!?7k�� �����%�u㣾���͎�w{`Ym6\W�������S��۾�= ��{��&MTfsRu0#\J�F??:v�q�T_R?�WP�B��)h;�ڴ�&
�����c��F�Q�!�W��_pp+X9���ۏ|���sR��j�Γ'Pȓw�K�5�
�61nk�'�BN�>�9���-^��
�0�p�D8�'�X]��1	�Lk��b� N
b9@+oz������:-A:s���)��Ϩp�c��y��}
�R��Jw�����K��܀�"$}x+�|�?����L�����˫M�(�_}6�J��sWwwZ� "Gp�"�>���V��y8�=�e���r$��+lk�D�CŖd� ��F�)f��;��ҷ,�n ���ݥa͟n-(�A�=�!�\ԐK��	�S����Hl�cN�	�p��h�ڸ��:���G��S�A~PBM�@6�lhG�M��*y��E�K��K$\���Җ� ���e=E %�kP	=�|� ϋ��L��uM�e���T�P���WF�gDL|�s"t7>��̆��4��ЖC�$%�����r��^K�>�����u��ʒٙx��=�����c77��њԂYXQF�S�7��ֻ�"g��dCgRM�1�+~�STo�O�r=� ����n>5�b�� �?܅Q^�4Y(�G���Ǽ��5"����3��������,�$�Ŋ�X����w���m�oUZ�!�gǟ�K�$?1������^��`Mi({�D3}ɔ%�z�~�Cw7~R�*��G�T`�͈~0[�<��g�M���ϋ�u��d�k�R�x0���te�D���%�[ŭ\��ټ^����0¡����!�O`�C:�ԸS@��I-�����ہ��{���SFl�f� ���	EL_�LԵECu�V��7������X��>!8_+��2�k�ʨ�F{�u �[R�]A,�g/�3�A��{����+-�T�aW��'�����EP�N�l	7Qt��n��Ϛ�=�s��l�чy~���dy
���얋�z�"��8E�շ�"�ǿ4N�gs�h�B��ykG�_pd���N��VC�W��\�jFH^IxpeR����7�6;UEgꜜ��B�B6���[;��89��\��I�6��aKǫv�?W�e��J���E�&.;,2*(9�5$p��1��[Ct��zf���|׭��\g1Vd�u�&gJ�$����s"O�!O�Z�	�ğ|d*�,!��}�\�f~#��ּ7[J�t����g-_�FtL�5?z9��ՇA �}(������)��R\e�A�����F�F��g��J���~r9d�6Y���=fZYv�,��9�V#�o��k��9��y����Y�kE�jX
0/c��+�́�Ч��ؕ���.r�����;U��<���t)��oL�s`1��8��Ke����w�1��K��j���%�$��h���s ~�y��
� Ѻ�t߿+�Ɛ��a���fH>��<��aN�W���B���]����A#����>�놭7�)��{���q76�i6�0��Pj�>���k�^�/!�.P�����]G��ͬ'I��Ry�=��^�:�U6�!�#��L��ϫ�����8rU��K�y��-�Okx��>T��t�3��e�Oδ����m��~�/�=�O��1a��ޥqM!{:R?�䙻�o�nem0����	���,5h��IO>��[u�(�����?��g�Apǘ��l�4<��FQ�E-;v�z_�Lp��$��\f��C؋h�۔���%��=���a�  ��w�a'�XX��=���)�cOXb�ف��C���Ħ>ֺZ��p��R(�-��.��":'՝�Rw��=�S�_�R�*آ6�dlkx�����S���1�V}���ꢚ������� ө��)[���X�W@�m����y#��a�x&�[ң�N�%P 42S��.�1�[�����TS��E�������^&�2]���Z��e{�sy�ͻ�%xT���cyJX+��wҫ�r�~�����M�J4��� �t2�@'�͗�z���9^�Uz���'���SR�C���o�B�9_Y���ų][τ�Es�|���"
�E#H��ْ�����C�rl��nbZw�ÿ��U|E��0Л]ˋh�&߬�N��\�|N��Aʸ�˥�XR� (�3�sV�u�z�؟��i��-���5��O�,��9��Тj�h�Ra�~�a���Ji��~GW���;�_�����m���Nbk�gt���X,��2{���������R�>e�G�;Z�8ry��
ן ё˯Oq��ń޼�b;=��}�=˷�FQ��#'�P���IRk�j�!f�)�'t)OVᄻ�H?)@��W�QYz����h;>��-.�/_)�>k�e��G�N��t#�q7���k(_�b�}2xyۦF�L��}��%�I�~��%�����#��#nY�m��h�u@�Ƣ�	[�� �S-!�QGx�R�u���u�>��Jr!ߗ�K���s@�(���V�M2\f�T�����"�@�l".7�?��U,�E'�V��-��B��H_+������r��hΊW>:oZ߇�c�P����S�ԛ�G�[�f΃�U����/0Vb��L����O^8T��Z���򌟡U�����2����
�)����gf$��W{�.�z�0k��h܇�UwW�Yp��w����7�ز��*m̐jmo�����9(w�A�H�$p�.}��V��MF|��(�OZ��{}P0�7��� ?2@��7�Чi6�kv��Q�a{�sM�W��08e��J��2�_P
gFo�����Ǿ���)=o�)>�[�����D����.T�� V�������6�䋞�`�������&ϟp;.�����(r4�j4'sґ����n��{R�a���ݒMu�ͫ?���X"��v��h�HAM(���Vaȕ����F��{|�\��1v��������TsjRQ��]������A��4���m`H@���̢?�}`G�5Uʬ*�M,Lq;68r���ʐ5rM�.�ftD�J���D;"���OGc�#g��B�w�����%2E�iU���3����$�݄���i���Y���bm㪫�3dƌdx�.V33㭽x�+>�h��dM����5ϕ��I���5;�d��Z��R+�on�u��~�k}���HW��V���yDd�y=�����$Ω�8Dx*`�M{���ẖ�	K�=�}	�-]�l�	Nh��B)<�	��rU�9�x�5y�Ծ
 R>=�{P�f�!���Q(��r�Bg"�4�mL��)���Ο(z���P_������IO/�&lh�n1���	 }��OG�p{�a��܈�К>�Q����NU�j	�q7�6s_mc��9�K��ڴ �5��OVt�[/�=��ݰ�T}8H'�r<�4雷8U&6x��䯤��NH�J�J��C��ͺ}"�T�$�z/�~E�J�X:3�|�����P��p)ُ����jV��[�<b@�b�3�%�b���(���sd����aI��<��@Κ83�b�y ��j���$�艁�z��ʞ�e�]nB�J���7�ݶ��,[]vN����B���m���$
C��>;�lU�������GmamT���ӝ�R��_�%㑉5�^5T��֮k���?&^�'�ڟ��].��q���G4/�8'�VV|�d���f�G\os�1���xn>S=�a^��JlAE�6J=Agf濈 TL'�!5��t��-������O,˅E�Ί)ls�};w��D^3{Ԧ����_N���:(J��`��3�x�T܏~�.G�u��t�丢��P=;�������!�M�4��3��~M��/,�c\�x0�՚
#����h���ɑ�j�l|Y��yQ(�>�2-9�G2���w��L {�h�*�3����tsf�?yL���~Om2�ຠ�
�w�kn��D"�Ùĕ�tG[�n���L��M�/}l���+��;���zeefx����7�{����4:��l>E0���[�`9�~�{j��t?���q�i�ڬ)x
5��Cs8t�~�'&F�J�5Y�Z����<g�VY���|��x��ǜ�T4��
QϺ��ܸ���5�u�!Eȯ�_��cr�o1�ڳ�cI���;%�B~��$&�O�{~�2�ی�בw��~�qLq����f�Ŷ�h���;��]��:�ə��O�3A��jjӇ5e��˷�7_C���|�ɝA���J�A\h��9���dꎛ��l�ox��5��ϯwo���j?��$`,Mp#�O�����WW�&���Ó��.�І������/7^SװA����ϷZ�(-�h��F�kN��Rl��)ʂU�_�6��:�VA���L6�W�+|/����p�f�cW7t��	��<=v0�sҒ�N-@^/$V|�[]��̬�j34vj	?#9R�~$�#�.,���z�r���"������ێ~���ȪE��d��v���ư���u�����7z���Pt�H`�Lt��~_� �6ɹ�G���2��7�G%釚�vH�gR��M���*�:�MK��~dN��XN��'�G�-R�3�7���J�. V��,+΅�4�3a���n�y�r�e�Kt9�f����ķ����2M$`�qTԃq�죕��?l�y&v��������R��*,���Q�2c��%R0�w�/��I�%D�����A�e�Y������
�|LV�yB����m�_o<�����r^���I�g��3f���N@8>�EU���5�N�19���Dy��%���I9����t��Cm`�n���i�����73�?n�v�f�tT���+,�b�u�/_��� «�XT]G�*���?O�> S|;��0(#8S��r�'�*Y7kD��˵)�p�TR�d�O��i��H	�b:mN�Y�6S�
џ����F�!�vj����cx,g!�7{h�/�mє����:M]�����y[�S�������i��۫+�\�]��[y]9���'?�:�����{~}��bPvpl��R �������`e�? �p������]�����jP�Y����_�4�Ͷ���c�+�g���F�$���^L�&���"��y����) ��@��c�tX�r��O���ݜtH9OK̐H��ߔ��) �#�.y�c��67zo`BE�?[S���5V�ױy���;ґeY�[�~�-�k��w)Dܮ0�o	-,�q�])��2�W:���?�̼�ɬ��(��\�*�nGM!7�C8]�0�R��븅(q��Kl�M��h��ඳ��9_�������+���)H�A=9�}��R A�kr��g��22B�RU�o�Q?3��E~nz|���Sơ��	'��k>�R+�>�Rԯ���%mY�-7��Q҃3�ZbE�%2R[��?\����CN�?a�Jk�u���l�Y�����*q��	�0 ���h�K��b��`��,��Õ���PƳ]m�qB���(o�V�Z@��7Yu�?�k��^Jǻ9ڀT�./Z�ka�,S�Q��+���ݾ����p X(�Kp�"�*��#�_����_�+q����o�)���6��_��Tw�:r�h �r����}����&�s&�5���y�p�T��،d+d��5�1wI��i��ʟD�ԛS)�"ˆ�rd(�W��L�B/�G��<���˪�He�t������V\��_k\�q{�^�OO�����M�m�з6��o4�a�u�TVMi���v& ~�;�0/*;�J")rW�g.{D�@�L��mx�fҍr`h]�U�8̏��E��ӂ�˴3U���AӚ������[�~�ؽ�O.�QW�_��}*��Ȗ�s�u��:O�:"���{��*�}���1H׿[��Z ks����7HXKX&vU�S�bq��F��&Ո5[Ş����:��7��y��u�)$Z .@]��7Sk5G��N8)�i�]�?y���4 �������Fb϶�#{��KR�F+8vz`����E5p@�%�W˂������<F�����$�m�Q��n-��Z�ȣ]E-S�_;m~��#�4=�Ӱ�Z$�ŲL�f�Q��85��ˊ�D��41QUt�=bO��~P"�@�D�������cVHm���R4��(g��L}�944�,��HOh��q�Eb�v�2Z�B��U�"�,f5����������it��;�5cJ��z\:N��إ��Uy+����_��3:�Q�3�q7���$��?�@�y�r�-˪'��֓�PJ��D�?\98���]��u�W�qQ�U�t�Ƴ���Ɇ�7L�J"��<�~��i	�P����c03����=��D�:��#܇4����E�M{��~��J�P K��Q�X��vWn���4�������%��)���� ����\�!q.�o%!���^�Y+8o��a~�rA��rJ�1׌!���$J�I	���9=&%(�_mWU��!��[� +;)��!;8�ba���8Ю�-��t�h�c��]�6F���~���J�SmM_�4�M�,����`9�pB�o'�C�k�c%��Q㹛�=�8�U|.��o�Ɛ�Ʈ��`�N��w�W�w*���d��� I�e{�WP0ל��� ��%5�����l��Ff}j1��=⚀@�ӵ���Gn������n	�[Ȱ!))= ^Ds��ղ|�����S��O���%kx�~��&t�:�5�/�k�����@�)�B2�˝K�>����5����a��jR"0^�>�z��e*?�pw���2k(9P�Z�?SD��q��an8��DS�!U�%`�������7�r�}�Xݢ�!Q�$�=�Ns�8�K�Ң���U.� �d��H����b6�T���d�D�A���H��w��ʡ�ۀ@��M��g4bL
i���Ñ�X���x|5�mܗ ���5)��4���x7�O(��|���� ����1�!gέ��3 {fg�#;ɀ=v�4�]>�t�\�UMέ���S7�0b���_@�,uZF�� u ��f[)iG��eaJ�'c�������\�;�H�mD�9��)�
&���Nn�)ap)Occ"��ƛ���(��N���z@b_@"J��J�(�s�A�RK�'������`WaHz�33a���F
�] װ/�G"$���a)�f`P�%0��?/TF`U�W�|;�A��1��,RQ�#���%������!޷ 2Y�ƀ�����s��\�S��V�.���T�b'��zNxw�O]���n����F��n���_�QO.��V�^������ɮ��,׃l��>0W���,���H�1W.���jƭ�0���F@��Y˥�y��AB_f�Ӱ]+*ڻ���i��-I��:�������QH$��>K7���阙ht�iX��ӽ��	^�E#�ҹv��`ln�9c�,rc�))�� Mf$ɶ��|�u��{�)�rbw�ku� g)y৯Bz��j��� ����^.����̭K6�"p�Td)�6Q3�c�"aW�5��P�:����:Pm��ȋ��8����JӦw[���]܁x^��0�/?�2]-Y��-�g���Ͻ��4qq�(�i�c�l= m��U{}�F��w�Ǯ��Q���R_�kP6���zv�=2�����ET�J�e���c��� �N�L�" �&�+���FS��A�>�K0)�<4���(7&�~W��q�2�+=�j��v�e���,@�wٰ���L
�sC۞�>L(0!2�
M�Բ3�p�<�;#:1KS�j�ƭ1<��#�ךz��?ܶ^�+�h���n"޺D��?�@g����Y�nU+����������3'7��lx��p���k%{�PCH�#G��� =���(~���4\t~{��*�����U���&ܿtĊ����A�U#0\|+~��Z�Kre�	�a�'�}��IX�:(-��j�) ��Ɛ���j���ש '<��]N�jH�]��Y�n�³=��Ƃ>�]}6$?ǋ	�zEƳ��䒓�]��h�x,B�)-U�L���1���b�n�%<�x�lmb$ 66�'C/(��][)�����B���Tq�`�X�7&gf2�����6[H�˔(��NO�2>��I�g7�d��3���)�^�KC���K<�bݘc����y��=J[��#>�?.��y=	Q��͓���J�?di��m>s�6������%��.����V��OLb���T'�YWW��t_�ض��Ʒ@B���kz�T�@W6Gw��V� �.�z�s�4�
e\��!t��?�}��s�t��̥��2v.������D�&�:p��o�����EȂ��q���`����+�̺�{�܄r8S�X���]Ko&N9A���?�+���#�� K���N�� ��o�}��{�	��Oo���-��M�l �U�{��4�FPc�QV�����lQ��+��6l��YBp=��)�̄��`�u~a�� �� ���@Ѯ[���&��j�}Hې��oNKd�at�c����z-�����1?c���18����T>8���܃/Z{�"��w��l����������?�3�2٢9V��@{�%_�g�x���#׃]�{�x���e�>*�C��
���#4�Ҝ�������)p��U�������#V�"�::\n�:΋S��O�B�W
A��E?��a$2f�H ���u�4�$:��DU�����!|WWN�i�d�1�t��� `{��ؼܐ���Iu �6��k�8��೏{-+�?�2� i�1}��㜹�l\ ��%����	E-��'��Ha��t��� l
�֙�m�e��++z�XDG��w �Q����>YZ%n��t뽍���<1@Bv���5�l�~�c��+�a�����ձb���/����\
��;M��y?l%ߡɀw%*2�e�v��(-h���XY"!�0k�j���0��C�v��0����*}Qh�R�7��2��{U�!o�����m�ABNj�q�64z��J�gk�S������1L[S��s?�ZMpR�;��N$F�k,�?Ds��O/*��Ĭ�"��� ���%yV�s,КC��N+>X��gj���0��Jk�� ��css��T1B��}ʙ�xi��m�Y��P���4c!B��v;i�X�`U:8�֛��b�x%w��s�~�㯭I�J2刦���,�tS`�O��'���V���\C�F���1t���C�B?@���5��V����G�B�p�^׭��}.L�D�U׳O;�9��6H$�H�r|�y�����
�x���ICT'��[RR��������9=}��C���x�+㲷A^����|H���ǎn�u�А�����_)����$Jev�#�Y,C܍���Ax0_����C1�_�k��=�}�����N\��9ҷPEy��"���v9�j�
af_C�q��~�����9D�ӧ�r	EZ�[h�<����&��ǿ؍>�{}Ք��ƛ�{v�����ʏ�se�#�|���f���.HG�{���c�}w����JF��I��|�v��W|4�ػ!��l �o�j>ڍaQ�z�N\2Pc
����W��	��z�M_��-2�}E��(�hi��L�R=Ԧ�Lq&G���/�Ձ�t��a@;�p�q�ac*���X))�g	���AI�s�r���aJ�Y~X��ٵ�f������x�2O�2u�\!�6�u�,iSÇ7é��ԏ�"D����Mޑ�:�\��
\Ï�_�����-l���L�� 4����k���K�i5ז!��P�iŘ;{@>'-2�-6�����<�^`ۄ�Y�E"��g̕���sS�{At)�Jh:|��3�����B���R����m�U������"�Cމ�������x��&�%�+��\�9ً>�c@yKN�p�Qm�T��t藓�]Lw�r2������^��9���֥�Խ��d�ʪ���MϿ��d�����5�p3�P�>�N��f%���"(���*f�<u�c�*� <�4����0��N�(��p[�XY-i�V6�z���_lqk�I��9b~5a��F�7� �n<&^/,H��)�����	Ug� u�좲�J��ݠxM;Єi' �L鼛p[v&�6/Lk`��q�q�?��g�A����Ѹ�.�����>��o<�X8���Y��n�D!C�~�׋~Ma5z��
��_��aNCM~m7�]�NtJ�al�fcbQߙ�l�U$$�/"'O=X�,��u� �[�4?��@���-�*�7�}�e��soP�;�A
�<[��ֿ�Q�>B��n�{��Ql�q ��s����b��`Է�EIn�h!���Fe��GL����%#K���M�+��i��7�wms1�>��������a$K���|��|B3w$�G�����SƟ�_N!�C�^ʵ~B��}��'fҾ82��.����5��twݻԤ�Y5��mځR*�q`Cs��g�ڔ\���_�Z1" ������zR����\e�%tL�P�Ӡ��y�Ώ�2Q��XJW�|8�b�p��WҬ(�,�>��<���oZ���q�8��ٜ���}B����+�0��^�e�d(�F��gB::�j*oo3z,��q��f��&!�� ���vV��	��HBN�C�S″LH;�}����a�_2�ʍ�'6j�GG;u���a]��&��,���I=)��=��o9�d/����-�_"������f�p��6u��H��2M�4hA��XlGR$��E�d�?�J�Q��%$G96J��Y�X�L�A퐤���f{���&Ν�v��̿�pH�?�CX�R}Y�$x�s�yE˽&;���s�hE����4VDH���ߕ��t뗄��i��2��� �:j���I2\�"�.�*Q졽���1-�H��|N��ETa4��-\
j38'`���=�i��6��vt+��ȼl��8��}Aо��j����m�9�����K�.���!g���sFb&�azw�X�f
�4	�czC��K�����>0���!���?ӖI��v��SGr�Z�Q��2�HD�,
#�� W6�W���Q�G�!l��ոp���)^	ۢ��b���R����&�8��ĺ���+,�s�K'�2�m��~�P�׮�O-+�@��@���������/~�`��C!�5bZ�2Ai�'�e��~̔���v�4j@[K'%�k���v�čAE@�,��F�_�~�r�hp�#ƻ���˨��5,t.� F5�7�e�p��~�i,�F�����^']�<�Ümu�ʟ�Lm��l�6{Y�M����W�F$�Vz�c����7Ǘ�#v��Ű^Fr`�����NCѢ%a�'7Dh���֨���1[��쇺�Â����i*���EWT@�[�غ���z\�lI��8�3R�����Br���α��q� ��䤰2W�VyZ|��k��{��&����x�{�?,e�����'�5C�����Mi	��$�g�����؝���L@�q4���P[��L����t{��)'��ty@��Ac�46�ɳAFE��(�َ�:�n7�"��/�#�_;37#O�6䙏���O�񺌺�.!M�r)�C�٩PN���Gcq��8��&/����1B^���7�g=�hA=џv�o�о-~��y5�f$A%o0B�,���?���a(�z3͓����q�,e�׵GtU]����� �l_t<f[Q����R�N�_ �j��/;{�g�U�e�{��
�?1}���D��N��~xg�U��P�B2�������Q�O�"j;ih9na� ��C��ڈ��c�Q�v��h�d�����r�V��ܦ*x����ؘAXJ�C�ŗ���t�-U�LȓA$����2�G~��j�7&7z��ՠ����V�צ4qM'���v^Ysח<!䓨��^�XYg�\�'�������&/�1Q��h�h���.Ҡ粋%<i2f��B�.6����_KB���!_3�p!-��~JyL�$�r��N�i���W@,�l���z��
�?5Z5c��z���
���9�JL$�,%^�R���܎6׌���C�>��w��1f�=A���O�z~����O�9���J���_�1|%���]k����Q���{�S��z� �����D�ܘ^ٹ��oHu�d���f�U��a8�0�g����zsj�I���72\炊��ϫLn4v��S�Q�ZTq��\����E]�y y�P���lx��Ⱦ6�Pk^�����v3��;v�B�T�����;���G-v:�;Y�d�ԉk|>�kf%��ׇ�+�W �WKܬ�\1V���#��S�O�H1�䓩=�>�U$��ݑJԕe�$ )Zh\�����^s�����"�1"���|��&=CQ��Y�A�� ��Xa�8���q!Zd�ޔ���'��{��������i�&�l&�v��Z")��uk|H��8{8TPJ&kM�@,�@I��S��7y�no��b*�_���҇^���)��i���xI�U�)��
_Ai�_�#�;�'F�����s0\Ə��p0~���-�:#᾽I-����aiR�1Z���4��[>+��������WZ5Ʀ�;�SQKg�L�ul#�����<��*X��`f��}w�y����s)�P&�G%�uT�%��VNT����k� Px{n
_����=طP2�@3�󢎻%Ѱ���G����Q{[�1_l�����8P��%h���Y_X� �WS������8�7�d�Q�\�B���˿�3�xH<�F���<2�T����zn_�Y,��V���a����~�lHz�6h�EJ�N� s\B5�Yn��u0�p���u��fG�Ň���r�_#���n��	c0�����U36]"���OT&����x��]���(� ؁��-��C%m�?��''A䏅=����\���a�JI
豾7cNݦ��M�>�,���='�|�K��ȭ� E3��]�-�!�,
�A�ƞ	p8�2�:��,Y5�G�j(U���(�i���?�l͢4$z\�Ӵ�8�f�D���@G�#h&aӭ� ��N.��X��ɓ��ɄވHpKq	a"��V&Y�SXb�L[���JϬ��/���G���F��'��3���t�`�GM��w�|���!.d����.�����/���K���y[{�����'|�h�t6%)Ιm�^�X2h*L���oˎ�L�:�;D��/+ ����O�Z�U�UV�<󜣞$��*�c�8���<���9
���%۳#4������d�#~�`�g#�趰���`�=X_���{�>���y�i����z_����Iy�['��$�p�t|W�|�uKM���y;�S�*x��:�xR�Ũ�N	���&�R?_X�)_|#��ZY `�A����/.X���$ƆH�	�t%����
(�e�|LEA��<��o��,���QnwcI�N��Xh�	�#�	ι'F�9�E�ݧ�ɋ/����%FDΦ�_s\�F�V˿���eE֯�Y����)m�u'���o����}z�~-.�5���O�:Z�q�Yӱ`p~�F�ٸ�-:|d��l?J?j�2�04.Bv􅵽�����!�[
��P*�?�?�+L���V|��\=\��{����W��b�H�ec��/������a�ݖ�e����6:�^$��UE;�H�ah����6�L xgD�!z���^�9�m�M�P���L�|��D9��͇oF��)3\�(�-�6��n(l�VGJ����s�ru�cC����K��bN�Q�iL�p�5���~��݂������:ܪ�y)�nu��D�}�ѷ�^�)� c�#�>G��J-�n$��@vNl�qg	�LӴ�D|�B��y��@rQJ}��?�#5꩙B;�m(�у����8�3�h�
�h'&T���uQe}���*�t�.$�7h2r	
�'n|O�\�,�x��:\���7��嚅:�I�`���J>�=~IN��*�1����=���>�k���xj��"�s�.y�hb,�W够MZ������='��*��)�𙖺�������H�I�D��`�Z�x����oZw�2ɴ�pb�>�x愱�$ܗюṋe�I,PV�IQ���&�&�*�Ė# �)��f E��?����⼩ �5թ2�����*��J��z역y���UX���]@���K�p�4F(w�k�?���ƠX�p$�ѺN�L���[�ǒ��w�}{��l��ёԷ�	b��㡖�Ex�N���֥��q�I�l�N�ϣ���S�����ż���A��pTl}C��q΋�/�5���'N���2d�8lo�2�2o��OT��x�PQWe�e6��:�nfU3/;��'��)�Fb�Z#AѬJ�[���A��Uc�;��HYնΌ�/�)-�t���(�&}7�,�1��p�2�gѺ�H��.�\�ƍΩ���1�ص�v�tX|�QԔ�)�\/���\����}K&�x7��`ވs8Ҝ��r��)�u�d�p�!��*y��PR���\n	;}~uq��@�����lo��nQ)�z�`zbΫ�=�5�R��2>F� ;z�>i�^erZ�=m*	U���X�Y��v�d�]�h�b�tu���ufV�ݛj�.S3(���缛F,N}�D6�����,���L
��<����m����qR����{�;��e��e�b��������i�W��gW<�G�~��?S�XM�*[VE�e@���k�sW���]
P4���;�r�:��B1+1�Jo"�	E�`)���=��$UmB?m�:�a��.ʼ�?s�ϱ~|�Z,e�f ��G�� U)�=zG�)��!��j�[��2�qʄk8`� ��E�&?Ћ�ߡ��&�
e�<<;��qib�9�)��6���/Z��(�O�!|�I��:�J&�Pu3uf(��s�K��m�����S0�F�����lF��w�$����qE�a؃a��K��Jt=��jz�"�B��Ŕ�A�d���~>@�� ��Nݛ�$B:=l�Ko6Z�+�{�{T�5���a�_�&�g��+0���j�h�h,k[�bj=��k��n�����)��c����&C�O�q�_�dm��4��<���b�񝔗��}��-�y��e�؄�#/˶K�.�D<h�W.�zRlR��8�B@Kaʡ��&O;�;�R]m�OxMP7�,M��$<�<y��N���6���儅��(D�>$�p�]�3�����X��4Z>δ\V��o=�'�c��Q�t�9#���NZ�??��G�ew�FJU+�z�����<-�½���{�e~�]��J�
���̝�?}�95��j h�[nj�D@��1�&�j��p��h�G�J����*���W���Y]|:�`(Fo�T����o/d)�q��N�N8�F��׋K��Uz��I�N�b8�-�%ɔ�����j�S��B;
p��\��L\���n��З]ӥ����Q�n8x�X����o��⠡�L�"�Q
}T���`�iC��Gob�'��(ܥ����Z+m"a��h�D5;�f�)t��W�3�f� ]����c!N��LcP�j�o�Mz���~	�r�h5�L���D0���k^Ԫt� ��V�.�B������	�ꈚ��5��~�����e�!B%��2�䂭��O�ή��p�&�ޛs��Gp�n�gA+��y�Xh/�S͉��Q}l����������]#���Pz9>�$�m��Yq�����W��K�����oK������m��n_^a�2���Y��t��K��d�~x��2Ǭ�[�lAE�Px���|<�q�3�� �@��4�A��QXpК6��v��P�΀� �h��q�� ����)3�zĈ���ME�L�y��o�T�^�,Z��Qa��٠-�0W �m�o)jև$s~�������޲s^d؉�J2��5�Lo���w���p�Tv�r�ve MK�<�/_`�Y�Ð �a�L"�܍�O{raY��i+��v|5����f�ԵCY5�����{�7�Β�V�n���K
�Y��K�|5���y�ŃռW�~�}��BT��[���A�}_�JD|E��J޻gb��G�ƉmD��X~a���6ຈ��<DD�㥪�e�3P	�M^�_;3��~Y~�D�<����{s1?e+�	�ED�	9��k9��%⍩}~���,7�>`�d����ib!}�<�L���'����]�%�!��BI�Z���>*�ay����e��I*�2���_Q������]<;����8����)BaQ��ɾ�^{��M�ز<�r��O����P(r~��֞}����K��Ƴ�r�1�!��a}{�$�f�
�:\M�]�9�x�:��SB��|���P��8���=��F{U���}��Z��0�}(_b��7�7	�T�)ŵJ!ezL���<e+:��\œ.8�BjvO��L4:�i=i�����U���h�'Ӫj^��-�(��d�\lp�h�<N������#Qҗ�T�33� 
��t�ո&�5%�!�{G@JFg��:�!
�5P����h��AO�Dm�܎Q��B���f�B�1`�Hs��^΅��D;;�Y����Ċݹ�4L�4m	���pE����B�Q�M�v��3.��P�4pE�Z��6�}��z��yy챇͋�>����CZ��m�֡Z.R��V���`D��iNݷ���i*ʸ����j���,EJE���ǉ 2�^�B��������{;�5��x5�jW�@�L�|�t���)R������?�z�cm��> ?.yf�4��ܘ��w	�	�=��D&�����&{U��\��'[�aП��f�ԝ��VMe^�b�̚�v��(� �����$#��ܫ�k�H�y�K$m��A�a�� �%;{�_a��¹A+u����8�q嫮5���$@��jχ�~G��&���@s��hD��O��D�@5�m�V�A'E�? K���#߾����̹��4>˨�ز������
6�iJz�p�n\O�:���0�|֋��:�l��ޥ'#&šM��gn`AE)O9����$A ��+&��W�&��%P����t�~5�F(�U�?�9�wL��B�ge�fj��T@��u�"p���� �|��f����d�y,�Z�)��#�m�!8�-�`��� 5M����X����z�I=�$��;;dF�Jh vI�,N��Lp�}��J���C���f�����t��s��Z8���l�~��)3��z�#!s�d��E�Ǖ��+��^��o�����eP�wIO��A�n���O�f2Ua��X�`�P�
��ܬ<%�J�@�e?�(�\#p��m&=��Y3����n��4��Īv��9���yI>(����m#YY��#��Wb���<��&�I��Au��k�C���hiƯ�$���*��.�`z9.^:P��Z�J�[��4W�G�� ��y`����������tѠ��yqw�D��K�:�nTJ�JVS��݉�4G���(�7��(�ݙ�$.zgA\u36=vnn}�IE<�*�TQ���)����gᎄH�6�N����jx��8�!�k�*Z�����(�](�����_i��k2i=j�u��^L4'61ũ�+�r���?�
f1�|�`�]0��EE��~�ajzqi���sPMf&��O�h�@Z�΅(I�"RS��������[��45��х����ybo���M�.�B��8�����?x�Z��:���t�d p^y��9봵 h��&��δ�6lĬ�7,VP�o���w�հ���0.�%J8�J ���֖>ϠVy,��x���9��)��J��_)�DGs��Bj/3ܐw�y�&�j���A��{giB�s\e{G7�~�{���!K�շ[�4�2	�;�厧QK}i��-��.T��F����k��[/�U��[
��C�B�`v��g×�-���ri���\V�2=�M��(i�~���7l�+ۜ6*�[���T����m��Mc���)����|U��|�TI�l�,-�F(��wC_ɴD� ����?��C(tٖ��{m�@�H>��> �HsT�Z916�2���[�v���i�m>8ۗ�k`}�P�/`���K��#����wϮ����)�GN��B�� ����'7�Ao;;��d�
;GS*y*�z��,��d�"-�콆n)S�7��R
�7;�V:�2�������j�	)�^���x�������a��U^��w��!�J���F���J*�t�E?Qv�wb���ּ]�,w]Zfnm���|w�o�B��N��<�sx&�-���0�Z���"w�]Ц����]���9[����$���Q�	h� (��>Qu�!.�	%e۸-F �u�r7{���{-���K��L�h�(o�1�"�sx�����D������kV{ƶ�;�|����S���2� ���]p^P��h�2+[��$KH*�;p�i��V�""/ߕ��X�	���(�JsB.�-��j~��P�m�:{\�`E��MDe��@�����Ee>Lb)#�P�[-�"��l���j��6G�&G5�s�tѱP�?���Z��j|�IvY���O9�?�-�t�e꛼l>[l�t=��XGt۳����g�}w�dd��|7����Ho����Tvt ��\���A�u$�)o�1��:�u��D��J�l�nW��ߟ$�4LQ�eo��Q�����Ϳ`g�5��F�o��p�m��wԝƥ(ǝв��,��*F.�:��gE�4į�l˸�؍[�2��g9m�Lu��f���2�V7�@.��O^o>������0;ka��z
�ղ u�h+��YG(*.����qXے:���n���ٻ�0kᵿI�i�w�'D�C�������<S�a�2S��,�6S�����px�9�4d�&�c�B7�%Yi���7hWer�Oe��W���,��g���W�g�˂a���(U��l�c�J?E#�A��R,X�g�%��_�f� �Ҡ�y<�����<������)��Pm1�B�,�(�z8���Qc�_@O��d��Jw�T����!v�jPޜ�Caѹ�aNv�a۠�����]
�x�8�O�jn��}y1O�:Ф�ى��{�V Aq���>�� ��(�;D�bA���1u�GS��6/n��\����߭yT0`fz�.�y��C��<��Z��/��]��unZ�@�&|��*&[�l�r$��?�Ot�æ���ܦ=<���|�����u���e.�1�MN�۴��4���~5��n���A{"P5Fyؒ����[�����o�߸tY�����!��oO��OY?<�na�t(�< ZWP���+0��i,&,GK�p�U��p�+��~)�)	�X���,߽ƎaZ�gKKw=�%����,
"K[��|J�n��̢��r�pM�<�e���jx����(�&zV"9v������%!��NիBN�������OC�n��3$C>�'Yx��1�
������;]sk�p*�u�'5=�0k���wFm[������+����n̼ZĚ���.�u��<"�d�n��)�9Js�l�ײN�8b�p�t��W�$^���