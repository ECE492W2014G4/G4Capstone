��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P��v�"<ߞ��&'��k%P碶�R�ӣ�sĞ������FY&-揍�2�v0}�B9be�[�4��=����`q!���Z2M:��:7w� ��hZ�0��!L�e�}�K|���٭�y��?������^�	�#լ�LE���?����43f
����
-c�̿NS�I$�SQ3�5�W�R���Ǡ�S��>=��#5���2K]�Y�)}ϳ��ep9d�������,?#�/�4qW�72�:�йAr���T��N��giyUt"e�CP����TQ$ҽ�4A:
�/���w8�u�	e��P�S'-����y?(x×��{�x�g;��fґӋ����{"��l??�� ��ߎ6�i����O>i&2.�[���ِq�ſH����I��p�4ő��Էn�*$'%[Uj��Q?��T�q�ۈHu�]��Ʀ�� s���Ԣ�Zzi|��iPF���P�{�$��|��S��{�c�\��,2�#�T飓3>ȯ��,��|9�.c:x|�I�y��j��T9�l.�e �1}Ve��2.'V1\'	Pw̞���b-2��d��aH�Y �J:�浳p4oצ��O�6y.��h9���T)����ŧ��|V�ti�(�ёIij�oR���H����($<�cEK��,l�#1蠙�2��
���B�o!􇶱�6pو�.є{x
K�G=($b=�B(��,J���0�:��a7�t�Bpq ��SE�������c��h�n���.4:�~���<�o�ˣ���F����d4}W3���b;z���Fy��Ȯ��G4��`�倰a��lޤHU��z��~�t���mq3���u0N�F����ߴ�<~ݧ\*5^s�1��k%��F���#��c6t�R$�X�^�0�E��@O9c�nqk�d���fu�cۅ��}t�F��K�O��|�쉶���4�"��$�|�aI�"�,�-EsN2����	���*C�����{2ߪ���D��M�Б��o@��t�D�Ù�^p
3���
.��UJ-V��<W3�T�I�_���տ���續Oq���6�"�ܵ|KN�9�*�>���$%��P(X��$�M�{/����&�r	+�`]��,0N
�XF���tu�D���k*�Q��b�W����R�՛ZQ�!����pƚ�_��%�
ˤ�,m���$`t�Y.��q]D�'�/ `�'���͢Yh�~������^���q�:p�:���s��q��k��g:�)����D:��3�$�ͱ�R%�R �%(g.��:���WP�,V�m�����a�*S��M�3�9ħ2�v��� Z{�T�H!���X��e���C4�K���p�6�:Yҵu�۞3ءVuI�ѓ�b��8�s��XK��rD����y
����m�C��Ʌ���V*WKHyGm���[s�����ɺ𑈱R,	NX��wr�z���"�J+ �)a�x7��>8
i���Mre'�E>����Y��%� �u�����G;�䏆�Ɣp�0$m=j�����׼�5ȝ&���~��I����J-$�מ�rc��?I
���'F�����7���1�b����߉�⧋�}���MH�$V$��v���U	S<�*�J����eP�a��%L(���Iw�~LТg�~A�2C�*O H��Uc_ߋ��( փ�dA���]S �YF���Xg`p��7��=�+DUb�~4[v�<�X:�%���e;�T��VةU>=�h�Ր�yx:q�UCUa+���2[n�=߉D`���&��Y �5؀t����)� �֞�<�M\&�E�_�2�Xr��\�m;��i
s3[��FlH"���p�]p�P�h,c\���\�1 �szg&鷀<����O�>���h�DgH<�.��PӵZB2�¦���1��hYa����*;�G����m�Q��Jbh�a��n�5Z��
>�-i��
�F�F�/ΠY;�.	��k��H��igN�jx�ׄc�((�o��0K�J�1h�ꇵ�`�QM�����Bo�!Uh+5F��!�_�+
} 
~�U��zN^�fW
;�A�~�K�ls(���w���#8X]'*�>����*S\�F���}���E.�p��VC�1&�� ����a�D^3R8�ά+V����1 ����j�> 	�CU�IԴ�Q����"M�\�,_�>�U��i���^�[]�KV停�E���pZ��DR�z�6�:8���=�W�� ���˩G���3{�&�A����L�oY�C�N60K�o&�TS��$Ao�K 	R���V{�Ŵ�TBQ�6�Fઇ�r���J�ޙ@��`��Y&�M9��i@�o�{��iVu���J�4�����2�(�*w���>�~K��}Tю��O�Q$,D!���ձ�Ժ�/l=��I��:��!4�*-U'[>�b��#�xoj�Y��%\�m_9^MT֧ӗ�/�PT�<�����nx��O�P�T��c-|r�MC��^����[�fM4�q���:��o^����B���'��� �&Z"
\��U��z�u�7E�4M�6 g˥�Y鸁b��h۸ॄ&=]���Yi~K5����v�!s�6��æ��	��2������6Oj���=Ǉ(y��G��AY>�Z��8iy���L�R�򡵡-?k"11��l��J�IR�z�M S��#˷q�6�o�1G5��y���DeA��|��t <�b��h��3�����)rx�7�5SA';�T��?�����K�'̃W�$�*lW�ʑ�g�8�Ov���4�qJPc�w|�	�9�t��z��V
��کl !��O�΁��49�R�A�ތ�^�,���G=!�� <[j���!�b�:���b�U�h��O������H$�\xBʄ4�ݠ�!������(�՞|�ǜ��������� K�ÌsCA���cm0�G}����q����v�f�2�!�<B����P���S��70�q�|����
�
h)�_���<t6�Z/�
�/��
���K�Tw�L�Ђ�Aѷ�d<��,�X�p�U���u�W���"g���ܢw�Y��a_oL���)4�w6������׽ZB��U���BC,B&� �}��y_�1�T��,��b��E7�\���Cq#J�G�")f�����~������!ϯ���|�J���)$���:��-���_Е�$�+����0S�w����X��9iq�L�� �R�F���bH^
�A����D�=��Rqa$�c�X��s��Y[J�W�H��
<��FO�����j�̓ �w��6����g��}�|C���_*%x)fu��n��$�ޡ��r-zss�Xd�)8.��cn�GHO4������\�m} ����e;$Zj���>~��̚}��1�.��OR�M��Ik����L�|�XN#�|��(�a�G/;E��*���O�2��Z�3�$�_6h��)�_P�76�`����v�k�(J��	�c�lT¥�]g�`���yQ� d8rp�O+Bw�e�){�,��	�*?�' 2��3�fǂ���3�b]������ef�M�R�%:��������|�1A�+<8x�^#}!�J��)��+t�/���u�پ�����p�l���#��C� V]�T]�r�C�E�c�*C��~���C���
m�Y��	0���?�U��'�.+�Y@\��20D$Ő��o�	�(_���I�0�x������(�.m8��F��;��r�* ��j���g�<1�j�p
��:�9��K:>��:� /�����:�a$��C�I����Sڀ9�1�Rʆi��i�X=0�Za��ob�%�`%]����.����-/�)~@h6G�Z~������NW��s�
�S����'G��cšv��5b?��n�.���	�٭Z/[�fv�}�B���n^�<r,M�gs�ōԭ�X㙀�;�~ �?M��,�����2k� ��B���NF�*��p���Ų�5�ZD��ʭq�߰� '�"{\�b������څ��P)ң����q�a@e�"��Hf=/��r�J��P��/���[��";/�]υW�B�]r���j�'� ���\�h?F��:Gn���U�m07�ӓ����5߀��e�gF��,��J��,��Mn6�E_��#X�߆T$�#����]��q�Jb���|�L�2�g-a��+����P����^ ��T�B~�廗�_,�.�[�BĐ㓒^m�i$ =����7���v(:����\g�Y�Y��ݚ��a�#�h{�CW��D���QX�Dֱ���{clc��W�C�XU�?�<�k�5��sj�]%�0����zI�[R� ���D3�������h��[p�[	���)re������h��P�[���c�p�w��^�	�=^6Tw�A�w���BR��e��GhX��T����7�~3Ԯ�zz�ۡ
��bh1��>��W��nRa��k���t�q�����"^�ג�a��Ϧ��F=��O?�KAZх�ʩ�` Lk2�
)}�O��;���,�n�O�����^ي��P`{���.I�u9�$��-��W��Et�>���s�]�����a��w����b����%� AݟTܝ$݂��6m��珘0������_��F��*q�/��f����Xr�\Sā��|'�VڀT=58!��T�����ik��d0֌�K�w߲{A\&z�7��Ћ��ܙ���e�!$�A}��]	�<�@�I��R�~6l���C�W�y��i������PZP.�T_����K��F���nY]#���s��b@�N��	F�/���!�Z��H�^Dq4
���Ȟ&��b����o�=�$�K��̘�vt�?��/�9�r�4l�Fc�g��L��7&�r���Z\���iU���\�&�	n�7�m�ѺZ�_rvc��uͱ�*�\��֭+���r:����(���(���[6���Z?�z�CB�����L��`���J��)(I�kڎ_A���b������%�n,�<'F7�V�o���|b��<�PH������a}�����M<� ���+��ʮ]����E�s���xup�WK�_��$�;(�2�4�U�t��t؉ǥ�X0[�l�nr0��*0o�ع�p��;]�*�sw3��F�	����ӳx�Z_~=9p�
+`��9M��Z����Z�m5|�����sȝ�������g������B�)_J>`�О�B��X�^�8����ؐ�1�H���8Y��.Ð9�)ϙ ��=���jz�|�{筿���1���M��੓b[�rE'�Kx����ܠt#9Y�QB��[���䁳dIRj'k�ES�Q�ӵl�%_��Ӝ�r4#И�`�y-�#+�P���[�P1�8DVw�T�?ܪ��p�{eزq_��6vn���{E�����OOB�x���bukN����i��͢vlj�����n�Uti3��\��[�f˷���Ƈ�Α���n�|~M7�~���SUDL������z�b[��o6	j�QK͂��\M�hIXQ��c����WcB#�6�j$҆ ��f\m�Ct���h5�eo zl��lch@���lv�1n!s��_�X�Rh�)u��=�r�e��}� ���0EY=u"�CH�u�R(`_�fL�HSpQ���S�PU���5MX��(�@ʾ��xG��nFA�i��5B_N}��*钫.�uh~��ٱ�B�*��L�i{~�~���L
u�$*�H�ey����S��� Х*�ӟ�������9N�hK�>;�Kύ�P'tP[29_��d�c��>`�@�#�'Cӈ	���z��)�^`<�f�&���km!��S �*�F8�'g�sz=�R.�@���e,��Q�g����@V�.T�6pm�%ĜI���>#
��,���5�/ͻ���G�E��5c��ӯP�����b�\�5�6d�Lu�ն��<�F'��ds~��f���bI��S��$�@�aw���)�!%��U�Pz�g����lq��j����-�ntR�e%\WC����%	ʹ�!z�S�����]��~۰C�Z�0�X�5A�%��D,���-	?6U�5AĂ~v��0�W�<*��TL�:NW�A0�<���������#;���X}�}�	��u���_���t�gM9Q�*;�G��-}�o8IJ;7a��3�g�{�m=�b��P������HCD-�}�W})�(ĴM��j��o0�k�s0f�^�:��X�&\��Z��τ��Ѐ�Apb?��#�	�� Iua�zH��װ0���Rl�� �͚;/����������?�_c5\y�k
o3�ؖk�=�I�D�h7Nu�w�P"쁮��{���>0EW�s��B76!3�u��c�Ǡ�e� �R)�~��_ۡ�FQM������b�g���h���؍l@v܀T#~q���_!�k,vq<@�Y��2��w����A�;=�w��͙�fk+���)#]�P۫��Wи�i[�� O;�H�?<f5�x��K� ��B��}	�jk狀A����l��� ѡ�@;�η'��Պ�D~�b̆��2G�XG��vs�%��dDc�0���TN�ν&�/������$�����h3ZQa���޻i��#xn���.�0*�w�B��2ak�l�V���O+�{(�iU|��B��43��;q;�h��[�y�R�}�2�y���:$V�ɾ�a�b���2iGn�Uy��7c�i��<��!����O6'�!�^��q�L�gѸ�����d�F���â�����[�#h�(�Fv��}S���@HR�j��&�&U�ZL��&g��Va����{#T~�q����h���w7g��]� ���3HΠH�Ck"=��2�{�\�|?Y��a$��w½��g�N麹Q�X�)�f��
�y~���Y�aC��6��n`������	����{�=�u��L��ʔF>nܦ���G��n�<҅k O��?�d��&��T���7�������_�é�=��1^N� �i\������Q���U@а͋}���RK9Q�w C�{F����T�V�d�D���=8]$8�.nl�o(��í����0頀�Uw�Q��D�9s������nTi�y�I�`OO��/�]u���+E:9i&�˟��%�.��"Td�6�������d�j�ٓ�C3}��j8�D���#=��A�U�;��\S�7m�Ҋ޶b�:��Ib.�A��_�@��B��Y1�n����$�	�/mo�e*���=W�u�*������:�N��ez��	6���ZJ 
!F>�_cLj�$���?^B����B�����)�O`��J��By� �X���+���]g2D�m͑Q�6���)��گ��{������Ǩ5"����u��W��(",����i���䃕�]杴a4Z���i̡�)�6�ЫV�����[�>	6]e����kܤ�ؘ�M�̼\�ko'�A�̏;��i�����
�z�f1��r/�h䜉�ܻ��I�ͷ�[�`�h���%I�[�
쵻��8�D�77��P.l�Ͳ2�i�Ƽܺ����ϝf��r7~V�r!c�>��[D�6xO��+�(]��6��������2R����-I�"q�!��	p�i��x@���b�[�z�����K���N-��R����Hܒ��2äA�ת!cq�%�j.��H"��J0��!`g,��_]�:�*?���a�1�����p�|��5r:�.�c>B���a-�G���xH�}*�⅊�2z��p�|a�Kq���f2r�l�"e}���}]UR���s�$�d�!��@� Gc������c�-��qy��+j�*�1UA���v5Z�m�+��w�O��2 1��9�k�D���@15����7��M[\�:��������i[���2�ޔ�;
L��-����yFz�-����Q�aB{uƃ5f�� œ�p��W�|x+i=��hn�+M�ް��ud�g��P�+��l�[[�MQLz �#�9�T9�gL��";D31h��y�[���U�ՙL�����H���wU�^�A�B?�;����
I��'��_5f��g�Q�m�y����N��	��2��"%ot?����~�ly��;��[[�hd�Ս	�ikO&}�:\�۱*
!ϙ���{{B�j`����\e��.+��Lu�ʋ�DY,��٥
��8֫=�u������YV4�X�HB���7�\!����N;��9�4\��eZ^�����U�AP-�/�o�G4�^��q��_@H2