��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P��v�"<ߞ��&'��k%P碶�R�ӣ�sĞ������FY&�EI,�8CFy����Il�6�q�c'���P��_��J(��KC��6��
�Y	�Ŗ){z���,-����^���&B�Ѐ$���9Ǌ�/�(D4�,���6,7sS����w��c��ˡ�v��fK�儣i�� �}դ��L��"�_O������׺[�TL�^��89�d#���g�^�6My%�[G�WvWˈ���(���E�� y�nG��I�&7��C��u�ڷ��{t'c׫ʱ�����x��
*ʛϏx����5�K�����u)ulU�� a3< �muJ�F�wځԿ�7BsL����+�m�>%	��lD�kbC�}l����d�;]�nѬƳ#�m����%J��(�A�'I�1�TnS$[R�[�Z���u��gL�O�8,�ֈ����X���gG��l�@��f1���CR���x���In��T�*�l�s%�x�Vj�"�CN�ݸ*C՜�F>�� �I{r�%��A�u�0F�����-����^o32;�P5c����t�Sv�!O�X���8۞5��DRwWV��%�?|����u�\V]�Dc�kc�;�wA�Pl�|�H�C��\�3�2��l4�0-���X��4Ɉ���䑯�ù*������䯭��@L&�;9v,��+D���S����]�2zō�K��z-Q�";K��e�a�P���>�{�����7M�?�\/�&��s�N��4�][/�/&��X�+��m�pq��2�PCz����)�ܨ�"кB����DĴ)�ί�ɸ{26��(���$�.��(b���V�Q�o�-�z�L]�^xa"[���j�(N�췴���o��1e�R�Tw}���w�w����:�r��آ�J���x��wM��[~q?���΢�~���f��z�!�Ӯ3��f���`T���8M9�d5S`�EpZ7x������( ��H�K����¨�P�?I��@��4� ��_΀�	OK�[:u)��K,�Ga��`���d�U�K��|"%	�!A҈����J���/��5`),�T��TZE@�q��h��.}"�i����D@	Ę��;l�̳g�Xd����}��?(�>�&' [6ln���''����sߑ�Ʒ!�]NL)9~�8q�˰�v/�o� �w�SF��C�d���6��� ���}ך�����zhV�C.|����Td؉����Z�/K��C7����}���9�U�.��>e�'��Qc��{R�x,l?�S��:lVV+ُEqWP�l�9H1��Y�P�W~����o/��ܐя�'>G�,~?>� ���,�>�4v6���z�5c�w�o�p��sa�#�%�:�5�r�Kڰ�*�È�.i�Y���72��_�mp��d�֮LIoeK�׮�Mܫ ����w�������G�2l����]�����sR�T[�-�ZW����12��z��e��*K6*8r���E2���En���/�a��'� ��ݙ�?���N�n,Ef�T�):M��y�F-������p=��eZyZEZDk��x�����͐.)%��/�J�)%��t�=�:l�>�hٙˎr�cd�!�WG_�a���ϴ|,��Xa�� ���Nͨ���0X�^л��m	�*{N�y+2"�����J�R�2ˇ,ލQ� R'H]��5�o�~]�@އ��
iS�LM�Zt�=0&&P	��� W�3�K����K�>u< �-��qp�M�`h`;����2?Û�͜��j�� ���gt	�R~j��R����Z��^8E�J�t�����;Xf����-�\_�[���H�vs�����R+�y���}C�{2n�u[|�oc�-}�O�U�2J���ںT=�$�QΛ��&��X��N�l^(�C��YlT٪F��_>v
p�!U��l��&�8�[w'�n�#e	�B���O�tU�W��m����5�/=����>���W�T�4��n�MxJ&�������!�����$c:kj^��� �S�5�.�X��J�@��˖���@B�(����$^���fE�c�헤&�~o��E����P2b��x��c���E������ ��jm&��~w~-3ӌV? 9Q�>cc����)��6�Q������vu�	��Q��<��j�|-�o�<�5�J��8Ơ��1<8c� �=a�ạ#`b����&2,^��v*�Ъ)��0�!�I�p���9E�?�ӎ�G?��=�b:~����M &$_���ϚG�D��MWKI ��p��N�,o4+����\��Y�]��f*T��`z����s�ocCg�"󣤬���Hкe*�n�>8�r�o������A�����4�Ҥ�^�+p5����@RͲ�Nx v7���Z�T��,��*G�:-ú���~�+H�I������@p�Z�3�չ1杁�hȍ�AD���z%ϐ�0�0�DS���H�P~3�e�ӄ{L<ϕ�?� �2�j����ה�֪�m01�"R�|���?��X���5�690U�V���f�t���G�\�j50��X�{�K���(n�#I; I�d ���nbk�Lb< ܣ�K�e��ޖ�<5����,O�_�|�Î�ыU��&�ūW�1�ECC��=j��J�Gb$�|��/C�ոe?��>_f��Yhd�_[e�:!8j:��u|W᭒����fx:��,���.
M�;��T�߁q�L���7aq�O��y���k�3^������L�K�L���U�M��������@V��	��zN�J�E�!K����G����@LB(�� �+��pށS櫰Z�"��S�9�����C�2���J����]��˚_o�ͺh�SxFA��k���̹�Wx �:]�9S��~�f*g�ɳ��Zn8�S�)u��Q�0�r ���iKĢ(iX��e� ZX�A�\גm.�5[36���o�`R{�%�����v�Ik)o��[pVNf&X�	'�Ҩx�'����Pz,�l�\UV9��5zx.Gō�kɌ�A��^�@�8��n���N2	�x�>9lے�����bv�=YD����_O�C�6�çD5W��,	��?�)�y��8v9	���Sǃ$�,�e�.b����p��Kj�^Q��#�#)Z�0�r�q�b��*\yWf���-�Pg���P��Min�C��ɸ�?!����&X�#a/��/�,M�>c���1 {�U��|��5� � �s�k�^[�oVYD|*C�#У�l؞0sr�T0�n�Zr򫾸/j5|��mJ6F ���G�Aǹ��L��<�aut�!�����m��.�W$�kq$���� �ـ�W(kxi劑'�I?��G߉�����i��g�v�o�7���%�/��{5�J��͌]\�hQߝ������]ȝ�p�]f��ۣ�k����� ��r��O�c���.͸�ɴn��o(m1m���h m]t�v!_��_'ᅿ�'F����r�ܾ\��X��aP�� ���q��J<"E����?����}V��8�@�6��-6�Kc�^�n�`x ���?��]�ݼxuvᖡu^;�%iZڳ- �:Nc�t�º�1-A|[�l���O�T� ��U�^����[���8+�}��8]5�;?v��,��ĴJ��}7X�VE����G)�: ���� C2�x��d��; ����M�#^��?Sc�R���jB2���'(�D&�F_�&Y��$V�y��z�<U�7���%75���#��T�B�]��ʴ�+��#������yA!��#,�O�}�N��NP��7�M�Rh��Y��GݬO�
N4�
������`��(,��slӓ��m1��&�4�a���ow? L^q����[�8Cgh��:Ӫq⬷�޺�O�&y��*:6��g���^#����oYΫ_>��`��SoѢ����<h�vx�r�zL�H8�;�I����~lq�����P%/���H�ݒW��,��R�ɓ'�ʮ�o�l���ތl1;!��dEe=�O�2�\(�E1WV���
��88Zf�&z����c�E��͏Ñ���[[�S��r���0=�~ /���)x��;vNn��5�%��5/�Ч����FݦF[T��� ��F���Ơ��S"�z������:^ŋ�ɱ���Zg��{�D�W�-/~Qe�H��w��ƙ��i�����/��}�Je̜���K���&�j��_O�_k��q�=>�|j"N����U�Y<���}G �bZv�a�)b�\Fm�r4��S`�t"z��49}�X�w���g���x]�H�!�(Z�űN�=�rw�"�eW�� ��NI��+c8V8��f*�˙�d}��0�K�#�h�,.�r��A$�^a�I��eZ�\�91;`�����������A2^k�|�"Ó{	Ps��`e�1|x1)��K��Ϋl(��V�B!�v���F����js���a���jX4��������D[�.R�G�\��޿x�۠��X�o�T��f8�8 I�Pd;�g)��9Vn
w�q[H���ʈ�y�>*@ڨ5d�U�n�mK��j�t�ͧ� ���K|��]�J�f�U>`��i�#�ԣ��w�B���2j����(-HI�Jڒ��p�ߘ��I����yr���W�
� �-�G�*{�p�ΨF,Y������nF��V$^��~r5�A; �+�-g/��	�T�(��E�閯?�(1�G�W�ef���-�a���%�Uk��"ϙAx�)��٫�Ƙ�/����J����'(i�@LD\�� �-�0�i-$�u�|�,xC�N瀘b�FPD7�E������CЇ�F ѲnwN�pu��W~�u�j�@�P��b��sG�L��A�E�D �|�=hy�=O,k�4��B*ƺT�np��i�Q/5�rQq9$�:����@f����رk���{ �~z.T�G~�r�6�XC�O*$����,F�㓁��8�NJ�a�̨S3�N�/�_Cׂ����T��C ��,5D�?_?P�?�xR�@r�y�ֿ;���9��!�̜څg���u���B�mN;��b�����,���G@����y��E�k��y4Z���;r���^�+��v�C����]��>13cVE�/+�>V(�Lq(�tJ�6Y�T4�Kzh�nπ�Km�5k� �3^���;����|���wrmr������ٮ
|�X�����>��Ť
�1L[ �u�V���7��օ�v�s��k-�=ܬ�]s�"	�>k��Ia�Α���;��tX��߃�\��F�^i���Q<��;�5����SZ�3W� �ؓ� �i���2��*oѢ'��N���~���?ֿ�+��q�s�@z���!��ܛ�b�$qS-���$�S&�����^E��,�+J6Y��d4��
��M�^\�S?�ݨ�Kf������(
�N?N��r]t�v@,���=v�Cc�G��AzQ��ÊZJ�0)����\��E�Ƌ�����lh�#������>�skP�X��P�=�7?�>�<�!m��H&�ҋ.&_��W5�%��+!D�E���ϩ�n��"�)h�~l{�5�XD�a�������~'U��\%�=#�H�6�A{�́,L|���n��eg.�ee8�7PͭםF�R��I��i�5����uTO�w{w�ݒ�f��|�Zg�(�׏��#Y_A�W�_�[��P��U��+�Ijn���mᚖ�S :�b��<���k��Ꟃ�C��H�v��;;��B����~Ύ�uS�ʜ���M�� ��c�������M6�X���G�C|h�HB��
3�{����OI�l3rm��qH�����
�v'~i_F������Y�7	�G6��r��z���j�z�$�L��ĖBEu�!UJ�&���`�7d4I�p��	h��Y��S��$��m2���n=�%�#ŧQO�@k�}�{��g7����o��c��BP��L4��:�s:E���Q���h����Xw����HJW��.?��h�)w~��>t�d[��49z#�i�J+V.U���{��M,�:�l-X�Hx`��/ҼVM�Y<&,�E�yflA	�5��ZJ����MkK��v��
�y!^�v��
��:�� �E b�$T�ǰ����F+�sֱ5��dzL)�G	E�fBe<<g���ΙҝL�D�R�mf��X��vׇUDF�.�����N��_n^jP/��[w��'^%iB����h:~��x�_���k=���(E�	���ʷ�6m3��H�;��V���Gc�@� ԻA�)�H[��t�*+���*�G���k����B>�ӭX��#:P9T���?7 ��=7̎ю�JMI߽��R� s�/][��x��\�����Y<v/�9[�	�w�W]Jp�M.(F���Ey���걲oI��6�����jd���x	0bC��heX����Gj��ȫ��R��*��j���;�����1�����ӆɺ���fN����l[tGp,ʪ�����:���k�\��9�$�v�ZG㯔�8P����)������T��,󵄎%Sǜ��Ė��
���8Ͷ:�3"�q�h�cD���b� �6�d�启�[�K�Fej���ЬF��e�d��<�'�&��yo��řrz��?KC�:߱h|�-U,C{��(ő�H�|N �A��4闋@_���g�g�JOG�P^l-����~)|c��e_�I7O먍w%���ظ�����aU��g�B�yإ>zm݅A�]����&� �/��E�z"�I":Ye������n�a���k��89�v�"�jN�� -�a�fN�ϐ/f��/C
%e��AI��1U�!Gu�'#M��<��w�g���&�cJ�%��&����:#+�s x���x()Z��-��f"s����E��aR��O��br�P��Ƈ�������p�jʇ�^Vm/�S�]E+\�6���<_�C9h��*E��� �T ��ց
��6�oֶ���Y��U��fI�En�s�3�-���M�V��7GuG��`��(v��#�U�����6~��4�N �h?q�{f�8見p����G�S��	�����|���x�Ԕ6+`;�ri��w{��?��U�S�#��b;������?4�,S<74��;g��^D��|"3x.3�����uG)M��!T7�ѵ0���
jJeq�(*�G�2�Җ�n2�^Z;���ST�m��1<��k)}Z{��8�˪�OR�R������+tΘ����S]�P�T>�F.Tׅ����&ӌ6��m�1�YH
�oU�/^Vv�F7�J�y�Rn�)N�?�ꤿ���k���ۏ.�M��L�y�&�e��B�*�#;j����f��Q5�8�7N2V�:������fk��H�]%a+�I���l]��t_o����N:j�D@&����y�㺢�_�����T	8�\�z�i�B���+n������&Z�w�T���<Kh� �@_���ʗ���o���w�7O2a
Q���x�Ǳ1��=����u m��v��E�Pc+��zn����R����cQ4!l��`�V����ca;n
�Gg��;�KͲ�r ��	��'(�\�<�XX���9�A_��8'3��j������:j�_�3 �s|z�\�i�1�Ie��!����/.<Ee)l,-�~�V4�9�(�OC�ƻ��7˨�HzԳ��bB=��
�t�v%�:��qT`��dOh+lA���g}��~����Lޏf����@S�a��fO�O�vF�zT�|Ǘ��/vO�)�,���A�����0�7(��?�e|P�~��O�߅yu/VY�"X\��K�=�DxX��\���?<{�-M�饛���<5�{C��{�$�d7�E�z�n�y8턫�b���LR}G��'��6�P�I"\ ��Qp۫$�KGp�sʠX� g�IX�3QmjqJ��}��+V�y��yƸoR������B=$#�	����n�:8<(�t��R%
�|���70�P/�_��}�}�TZ����4f%9�!�~v�؉�̉�	۴�۟{�>��d�@�{r3%��Y9S�%���E���r�W�$F�[
�L��<(�����)���O�<�b�5����T�?�L���'��:X
T���>!��M�Ӣ��0T�Pk���kEp��4��l[�}����i�|Fxy�@UL.c([��r�?����ܨ���h�3�6����Æ$涍p��<�/HC�"��������. �V�AQxH�!O� K�Dd����\&�/�ĥ�4F.3�5�[Ɋ��],:�H���p���y#V���$�RboP�׫�ܻ9����E��w��G�K��ኃ�$%L�n{�	GW�~�"s��rn\���R�MO�3b)�mE����-�R����Gi��{��n˓�o��u<��u=v��#��x��}x�X,K�l�ȽV�ʔ<wu�CC�Ɨ���\"�����lx<Peʽ�w/�+�#xiۙ�h��微�j�i��o>���_iF��^�"�T-��T`�����'�����d�"~hd�?���@�Iܞ��@E��P��C(д"ko<'1�䄣{?�Ž��Ʈu���3�Y��b���YJ��p�B��_�/%��[��Լ'MRk觵H���;\�A|����u�i��,lX���Ө���ճ��оX��t�׳�CH�)L���3�xԄ!F�n��d*�  �����U�((|5-0�����g�=��Q)��e:��?�Zѳ��A�\����=4�����#"Oh��7������<FO���S׼V>���y��鸾�.H�r�.(n��N�'	\���6���%Q|%����7H6
�x�V�����N�~=+���uyvƙ��kMbg�%�s$�8�&���7����G���p]�?5q�5*f.��\v�p�]� �0��	v��˄T��*G�QB"P�����N<�W�;���[��C��<s��J*g����T�0����{��Z.���h���4C2^�:��K�w�g�m��$>ղ�	��DxYB�<��`���� �lܧS#P���O�@��a�0xGtG�o�(a�۶����M] �q^��9r��:�E�>�ώ ~��p3���P2=f���)��oI��jõJPs�+��2���a�:�����O��������E��k3���)Y+������J���9Cx�ԡ�����g�7Fz�Wc����ǉ˵-����|�0/�� ��B��E��Bq:F�:�Nz���R��V���n�(O����m�n�ŴB=&�V��L��P%�J�QQ�8���;/o���\9��|�#1@����8���ԀP,Spc��Ϻr�t��}D��wO�p� j�#���P#��	ڒ��ZBd��7�{�������ؓD�A�\$�iw����*
�x��>���&
ƈ�5�/���N3�r�|����m�Y�J�Q����gg�O�C�$�Cސ*�nҪ����q�M�J)�ݾ�,O�!рW�-A\3G����0��LB�M��饜/�h�e�b���'B+�j�"(<Eţl��!��>���A���9��� X/}p���a�2	��2>t����J�pn\:]Z�o1��dV�н&�A��D����V2��QA�0��=<
��c�����ȚV��I/!=](��o�
6;��Ln:��;G���s�#�x_��R��좥�C�ױ��=(�r�Z1���TtE�}�[�u�����ѩw��&�s�*[i���9�[�ҙ�?�N �jC������5lM�g2�q��T��j�k�wޞ/<�?��ɍ3����M�Cʽ�v������ý�6��K���a��ڦ#�T���cG*�e�q�r�/籢t7������C��DL�:1��i~��m� ���'�����	�>f�`)[��gq�s��l�ѯ�ni�0_�d���p��0;��#7�Ϭ�C��#��&Md�!%P����ݘ��E�u�8�N��Q��=���7�)ݩՇ�'���
�����M ��qG�OG�aT�M㵫�W��H��KG��(�_9���:8�#�6 ����߬�0�x�+៽��%����1$���I�p�Ћ�r��i'��g���h[���ѹ�*�  M�����UYM�>b�]��+�*X�����D����Բx.;�׭��QJ�jr��EAm��uσ�n̻T[E��B�R��!�����h��ǿh����-�Gˍ*v�1��>F:�LTL_7��)~O��CL�/&���'q��,�SF�u޵��[޷��d|k�b3�e�=L�7�rI�O���w)���5�M���t�_�c���@���l�� zI���T����T���0%�r#�W�����	�����x)%![�[:>
.a}��wm��y��O��Ɖ�b����_s���2��&'A#H<�nn�s6R�� ӹ�ΉN��e;k�;�ޚc���bQ�:P(��c�L`�g[�:A�ݩ%����x���=��A�<N]m_(�}�ֱ��D�X��$����D�X�dT�X\�C�I..hY�:�{�z��c< �?�Q�ó��c�\6mAy/���eVT#��6�Ǒ���p��e��Ç��T�WL���*%Q�m������g�v�`ͮY4�`<���[ߢ;p��і���ǒ۞;��y��^�v��p�<��
�k}W���o0�e�E�NH�:�W��#C����x�7���}����V�M���¤Ѿ����B;���@��y�Y(�'��f/�����S��{��'R�u� �k�Y8�<���g�]��0�홠!1᱃\��cS[N�2N�M�$��ZEPʈ~>�� �cȞ�
!��\ h (J�-���\�1Jh]N7��
Ѓ;lă/��J�?�Enj}0�~����í:r����W�76�]�|����k̬l$���H�c�Q��8��1�e��~��T���h�	`UG{�G�
��{�+��&�ˬ��˥�ݞ�����t��J��J3W%y���|�ӡ�����YQ�Wv4��|p����$�-�/��,QNţ��b��R	]7��z+����D��,k�C�f���+2*\-�!=��ь|e؇�B��+JH2	 ���қ,��җ�+�,.;|Du(0ea�A���چ��̝0�om�L7������Js��MlZ�x$�G�-��E�uo��t����׼w@�싆}�`�)Z�5D{�A�>OM�M��-�fn�8n
y/_�Z���I�7��׏0���y�j|�`s����+���v��:B����͞N�T�&5�൵��BVj��Jn��{d�J��_Z���g(��`O�D��H�:o��a���0���&0TN<�*���0�L{���TC~G#m����T����0O�4�7f`Z�-���y`�w���k�@1��v�AW*�E��|�i����{�%F�гL�f���T���z�6��7�j�6����%���]S�=�(��Ъ�+��kj�7�%�'
�2�#�+�����֪�Ko��Y��Kx���[
W���-rmp��.�r���z�2;KW����=@�Rn��D��e�U����T���w �rJ�!55���\�cc!-�L)�����o����36�������]��=q�o�:.k���
��a]]�t.�
���ui﹡6W(�(��t����.��u�_H��'ތ|v^��h�H}p0�k}�(�L�.���^�	�pK��R��]�����Gi����z�
�"Mז��j��eNH[+'���Z���r��5�;�:�!�W}��L� ����Y,�N<��n�AĞ�p�tQD�og�bbz@hA+ǌ7��'5�/=����⽭��MǔO�'e�q�c� γ<��Y[c��جw~��u@*�$�%�A�G_U�D?�E[����,ݿ\�gT?`9��J��(O�RkB�i�`�~O�7%�ڶ�ynue�cJ
cGCd9�����O� �xu��R��p�wW�-.��	��J$P�������oa=p�ˊ�*��RM����X��e^��n+n�o�J�yc0�PU��8+�s���� 6�3�9ª�+*�o���W��+]����
��"B�� A��N|����?&�� w�q�s���KvM����xO���gF1=)d�*;�M��@�*Š0ݞ���Q��-�1K�*��N���^��<�ͩ�o�:\�0�����m�d��*��ڌ�J󩽮x�*�SM�w�+�E����P	�r�R!e������چu�KV��m>�`gcT�N���QBl�wR��C鉝�d�a�x_M�����u�[�&ێ����Ԃc��4:�X�6���X�f�#~�3\[M�ֶ����I�Jַge]��=�FK m���$p��˜�R�o͚�:hY�)b��w�gN�� ICc>����\�,�e���rn6A�T�5Qd�s���!�}�*Wʤ;�c�.U	9�#�ȓju����G���Cq@Мk��?:��FY�q绰wk�CD��Py�m6�W�;�lQ0@��c�Y'%��K�6����3�|_ۃ	!~V �dP�EN�*�ڵ֠ ��v B��n�Q��e+9��	�(�g��⫩��ګ���Lx�R*�U	������9$����Zي�%M�T��^)�8	���^�1�z�C�%z$`o諕� f
%��݊!��.�nO���~�M�4@~��	z
��_Yx/	��X�v�߳�$�?v;�{���(a"x�>�|�9���׺�@��(�^���:u��<uAȯ�� ������r/�ejA������gj`t[�A�UP,�7|��LƳ�{̽>9��y����o�M,�㏘cƻȋ���w�@ A�t�>����FX� ��_����6��|xL���y�P4���V�К���1{!��b�̏T�tEW�Q@fۤ��������$_��׶�b�HY�|�km.���{�%D,;l0F��[���������##>g��-�g̎��f�K�4��t^�ϮT;�m�c��*�����t\(i�)m7&ʔt�0�� �^�r1�خ3�p�<��VPq��$Z̷4�5��E���r��b���OE'	孱Oq�2eTr����N�M�����^5b�x����6��Ί���,�%�O����¤U����Kt�x�ю�1��v�[�Fx)���QmGu�u�ށ���WD�
+Y���_+Ȭ�Y';)��W�� �'�6qY��:�\�x׀������ާi�[���\�E�2��-�H�9O���CfKFe�ma�L��$ f���UepcH>R9m�]TbRWA���5�z�;EE�Y	3�Wo�1�P]W���>�����S�8�
i63���=�HN,��t;	�U�^�L�$k.��ed�>R��j��y�")�J$n����(u��i�e��qP����(�n.��W�G�ˢK���d�=dc�1��`$���鄖��A���K	z�s,(��@~��E��|��o��LAp</���&�1ag�0YKq�C�*��'��b�E�1e�)��.�����R��F�]�>N�.�]U��x��W��ǫ�j�"�-��,�����`�a�9o�N��a�U:*���:ϐ5�Ea'`&��y��X�d!Hc(Vy�\q/�Dd�A���](��d~���4�����q�����ٳ�C,+��/��w�L�&�vi
����y���v�"��d2Ik�%���A}x:�d��4/�A�ϱ�yL@g[���?��zk���h-P�I���2Q��V%�a�s�1�Tx{U|0&u"vo�m�0#�["��;ƽ�-w�փpT�O�mI�|E/y�ȷ��:qAmvw���r p	��w�OT��}�֓��sȠ7��lW��0����T��g`��J�ɺ��6&g"�$x��?�\H�tS��\� M��*�%y_q�0q/�x!�9��~	��TN��l��.�#s��T�z�
px���[Wtk�Y3��ZT�{��_%Y��ƖWϠ�Q1exЧ����Qv���X�mK�P܈0[4��FA���w�!Y�x�
�W�F�d�p20���"rZ����$E�j�싲��=�(�R�&K?�?�����#�b�&�o(t�⦻9
t!� k.������
򠺙��Bc�Գ�x��oh%R�S�X�))y����u'�<'���GK�mO�7z��zvjj�(�X"8��J9W��@V�!�U���R�0�-�`r�҂�G�"7u&I�	����pw��lI����D�K�k^n6�X�2i%�.�~Z���R3��Vxq�0���w�����
�zЯ�TU���F�0��:	�����2����)����y��d�o��R^�G�H����_��c����tڻ���E�|VO�<23��d�s����
��t`x*�J�����<0�1y���WG(!������8A���@���'��%r�kD*?,��p#Z�PuJ,�N"��� *R.@l6�GA�������_3��'�~��)�e'�m
�b����?���4Җ�aV��� ���������k5p��	�P}<�eC>���vNj-�7��r&QR�jJ
��&�t�\��<��qvu��<�!�:�nx���*�bf`�����B��yTC����̖N�+��MH;9Է6R�a�o��w��ܒP����&V翸{bG�]���Z+K>6�o/�/`��� �� s�A��+"�\]	����A5�Q	��o�e���6=��4~��o���H����� �[&U3�sx�^����W��<k�o,a�Ҍ�P�yG�� 	5�]�/���jy�d28%�F��@�0a4
ͮ�gOa)�O�rv>�����
TIhā?��b���~a�9،H�)cSr�m���I�U]r�\�ϟ��V�]���"�/��B6ruQ�'ۤ�򖞕�Ex�f�|�ܦ��W�V�Q�������$��[7��c�N��7�'�$)"�*�FO(l*2�(�<1��γ>1eC����:�B����R�.�n>���ze�����0������-��f� Og���:���-��pY��6;�r"b���&�}�>�G�F �u�w�����=�K��G�:j������Ɨ~��I<2ra��?�P*s��`Kw\��Mݣv:�`W�G��~�Ġ-J�P�`egXȐ��aK�,�UY%�F����F�����v���4؎�:u��2pm�a�ϗ�0�����Dɋ�Ɛ9~��@B������}c�/�(ͧ�q�$4��i�����}�������m�- v�W�����r��/l��?B�W�*�@�(�gp`�śy��߳R�`%^&����m*�yw@'�c$#�"��HA��2�͏�h1N�nXU��-\�&��sz��x��B��XΑ���� F��͒�&C*�`�����8"��ٜ}z�X
�g/�r��6�`�R���ަ�RN���J�7�קn��M��eɕm���|���q��n���1P0۱uT+���ܐ�b��O�B�Efv�u漥,�>:�T���?�������EM�a0*	������=���������l�I"�I��Nث ��n����,��z�(s�4�:��.�=�ų��3!��e���8綕�-���&����S&'������������z��M��t/��E� \Ň��ΫV��і���I������ :CA=���P.g���"��͒�Bcd��=�~���g�}�kU%�KR�Hk�R�w`��L�u|����2���D�l>��R�[������E�^0=��f	e�"��Qw����ڵ~א��w�qTUq�RH�+�vN��٢z�6m}���6S�Ma��,hU�A�e5{��ݶr�H_:A���k�����n�^�˳E(���a���Sgչ4�1=�'���0��L,�b��d���41�$j��I�1�\4Q�}gֆ����׭4�7M��E�vK �F#�.�=D&�w�v�3�u�1�����IӸ�e���U�l�@�T��=r���?�T����_V��g
r�ڊY�0Hc�C�Ly����3��s3I�������=1nvK�b�E:�7��JW�@�{���lXO\etܖK�*�a��bW���?P�ef�{��|�t`_��iQE�Soo=5 ���CrL�c=�8���.J�
�
y��m5���#���[�z��6�����A��Ə"��P� � �0k���T�!��@�R4���l��ې��G ��Lȓ�Fe��(!o0�P�[Y*�$E�� �W��޾�����*P��D�PP+u��_S�IZ �ƛ�On!?�^����2`Մ@)0^�ݣe�.��˶�-����0�4=EV�|ҀH���WEg�B)��P�@��fH��*�K��
�Q���D�b���!-IQ⡅Rn#�˞⭟�4���^T֛
�)�d�Hut�BY��<�WS�رD�^ท�Q�#əT�`g���־���n��,�L�m�T@~��[)M��&�Sy���vC�7�|�¯��u2�w���i��=ŏx���r�f�殺�������L��	�S��L�9��ۯ�8Þ^�������y��(+�܁�wҌ�4u��Tq�b��`f� ��Qs�P�G��F	�ٳGlB!��L���B*�:��Q�$�I��ߞ֗$�$��c<o���Y�Z�T�%�԰�H*�Ã��>&�ۇ5��MG梒��Xr����ݺ�1��aO�Q�q7���0��K��P�d�d.3]��.�9��^����	k�*���J�1�ΎuGcoK�m�7�'`+���N�ӎE�����'|�!�c��&3ј����2���(c2�����j�C��w�3��Zb%���*���iA�C̩a�3b|�R�sʪ߾#�(��mN�J��;��V&JE1E`�z@��>�2���D�;Y�Y#�^&�c�z�,��w���}n��ew�*�jϸ�ɑ�T#S�EW��]���/�y�y_QkS�x��q�ɺ((F񺟡(wN�f���J��s�RhBmT_9�*b��hJ��_)zо�J�?/+�\wѲt���l{
��%�����K&ߒ��jˡ��Q{��i����i�Y���:w�R���Ĵç;�h�������1�����ZG�;���`���{O�Ժ i���$��H�y�n�_�7��ȟBB�#�#��Q��#��+π�V����u �za���י��J��z�伩4�V��Sr+�c�oo�%Q��F��PՂV(����L*���xʹd��&���1��xɦ�z�7)�8^V���@��9�FӭQ&qX,a��<�����RA�6y��[��YE��k���m�lt�y��l��(/F��SU�7We����$!�����m,��7��f��;\��jj��������.��MWgx:d�1Z>����e����@�#�{K�b���fi�y�S�u�D+��)LV�-�n��*����d s��
���)��B�^֡���w�Z�ۣCD6�d�YNz��� C���]4i�` �Z� �+k�jy����q�=��k�#T���Gנ�B!�p���"�؈�HPآh�c�~��p�,���X�v$U�mIp��� �fa���uYWH����y����ȱfK�p*I�����gyͷ�3���z:��y*X�7�ғ[�D�wV��0kϋ��o��[�'���S�xԢ�ض�ξ��@�O�G�g�?�`ZUFVp$�%8�20��y�KxBǡ��1�Շ��+c�I��%9P�s"KrW�p�L�.��ӽm������A5
d�Ky��h<�� ��+S�w]m���`�v�F.��jw:Y�s�^�&p���i��R`N��}%5�X�%;b؇�u�5I=�Q�ٿ�xȰ��H��������A� W���y"���)\J �2��=��9Z�͖�֒�+��3��T����=XB	��v����9�2'�{��R��¾F���.����S������J5��٫[�fc,;���ɥ�6��/Zg��+'�2��*��;��p�����wޙ��:��J��5.g�Hv:�����z���D�3���f\5g��cb1,.C�sH���3�ed�fj� YHJc���+k����4؜�L���(��HMyy�FЄj�6�&�Y}o�yT��~�yĶ�{��"Ա�m�8�p�Bxs�W�s�%Ȫ�l[�s��juC��Q)	����7�MUFS��Sg��i��ϫ�>s�K����n\�\	1ȟ�ro����ړE9{��mF�S��k��WA\#�&x2_��S�J�3փ�lv,���g�̍�@6�W3���c�+*H�(Ԛ�BQ��x<�����j48k�Y�u|YUz�����c�W��5��������}�ɥ���I}��V���Jc�+�Ę��b��zƜ�~�9�L΋k�������1��=}�DZw�zq��0�J���X�-��Z_��|�|,9��3*�.& @�cAa��#����6U�����0M�(6�Y�㱭�$��3���F�XgӢg�Qf���aL@��)^Dc��>���.b����w͉�b(�W���_-E��SX�\�K�c][����Y��4�������Y�k�&5��Ker��c
i���>.G�EH�:�
@�e����lb�/������7�֩�}|Ii�/>��(~�!��p���Gn������ b���R{c�q��
�q�����3Q���xѕ�t�0���RY��A�S>��ʉ�7*� t�(zǼ� i�H���瘠7�;����6��sC�̎�i�~gm$J�w,����҈�xh[ʏ�
�n�Tv�k�T�,k�N-N�;\�p�ڐ�S�:�r�
�hV�B�ܕI����h�N���.����7����JK&�lƎ��'r�3O:�ZJ%�ȑ��Z�_�SZ)���߆�˹Ty�bk�l���?���Md��6K���ϖ�����C�$��ٟ8�ۯ�fຬ�[p��au_vu�.1�Gd�|�1�d��<,�z��+�C��`[ퟕfT�r������rc�Cقh>z��t���kET����1SQ�-�u:�����m����?"�k�ĵ��s��@�/��J$TĽ�za��:�	��.w�5��]����量h܄��t�����3�uȩ'²��X@zV�~�tۺ��I�JE(�C�+�)��N����BP�2�p[��xs�>Y��1�K9I\�cR*�	�*-dh���7�M٤�����*��	
x0�A��L��଱A�XF����&�"X�w��]�?���Af���~��eQ��G�����0�ۓ��f���r���}�²�>���=��mWC���%(W�����\�����]����3HG�ubV�B��ӀI%s�-�+��;��	���&RWܽz�r�#�Oذh��]#�3uq5�AѾԮ��e5i��5�4��v�AV�S;8$�������� �ｚ%m�-!u��+�plk�1�a��D�&T���K�ħ"}v�����o4M�8S���:F�x3��a�$*m4"�ф�㸿�P�ES�6����^�æ��F�j��lY�=I<��sH�!�;�������5�:�W����P}���k�/R_�<J۵��}�S�-��5FJ��8O"D?�_)]hQ ���ލ/�E�ߌTJG��!������@O!j���!����<��݀=�/IZ��A�nm}�u�a1�	/������޵YK����A�E��?��Z�ԧ?��NyCȬ�P�{��.����T/���D��[j�Uy����T�F85ږ��P�Z8�w�~�3	$^�g��P����e���2��ڟbh�fԊ')�nf���0ͫ�ϧx ���B��&lj�b�\��� �?$��b��>r����`C�9mn�`����D=F�����ǭt����:On�[	F r8ik����5T�/����vR����Qm�t,�Q�+�2ٖ�N5"�b��?;����o���ESX(H�8f	�+J5��1m7p@��R�ݱ~���Y�Tv�����N����N	��{��"��S-Gg@Xzv�p�������������?�� `�hs�LU_����*����w],O�?7&-���e����v�{:��:&�6�����7�[�:�ӟ4�O�7B�I��-���x�~����5��x��uL����D�G�]��tp�Й|��܋]?I�`:�	�ɣ�ݣ8ubA�B����H�c3lГ�q҆�{;��p��j�ƕj-�[� �"���b\W��W�D}��?]֭J�ߙ�?�X�jb,��m��\�l��<���n��xFi�y֌�k�bo6��Z*��CT8œ�P"����`��t�T����k�h-�#���O��_@���z �B�Oo�T���n`z���Z��l+�9:Q�D[�_��@q�W!_g �X%���FN!�g"�G�Y]��zљ��C�x F��`u�셗��%'����rə�(���U�UJX΄~G«
������yK�{ε�x�~��ɴ��4�;&/?*�O�Ox6saA#�������K~l����M��%��S	��g%��>n+!D�Dl��\7���ɹ�� ����Q�;Bp/��ll�r�|�	8|S5��s�IV���^JL��w��[�h��d�]�䐀�I�{�u}U7q�����U=�6Q����ν3�H\[Y�hw�^c�ם�}^J;�����;���s{�z@�	k��/S��U3�=ֳ1���2�wI(L~?�'��n��)��$����Ұɏ��	\8{�21�"'�-NE��T���-��VeV�^X]��`W�Ƒ;@"#��<D���l@dr+g�"�?����$��Y1=VV��ظ�o?�o�˸n���;ےK�]��V�<ˣ�L�s���nP�ƀ@3� N*ps���L�#�܊C�vɋ�V��)J�v=4�T��to�jI��)��Sz=�f�u�Պpx�=�W�Z�H !떢�tߢ!rǆ�G�k��B���Z���l�������n4���D�|A�B�H��;k\Ъ	hČ�_�����+�@>�.׿����B���{}�WvB�v��x�GI{Mq�9�-��Y��Y�X�#�{�D�����FR
��>pQ6��i֯�VXc�w�x'�ޯsR4�$G��導��t�>+d�-@�����eJ�s��W�[C�/ն�����N�d���O�x�S�frg8��ۮ�ȎOZ�xS�D~��e�����@-+�e}]�\l�.q����w��E� 1�D*�Iq����XE�V+�%4𒿻���j"���3'qX�a����U�hG���j{ e 5�T�x��w_�؏.� .�T�5!��rٲ��kBH��&��F�%	�RK�j^�0�X�H�V�N5�\)���ys]s:�0Quy��u&CVtYMhՔIPU��1���3��Q��e��B�7�0,2��c�(���*�gg��^�wq��D�&_��!�����v8����]~�3�KZe~5��A���s�t(Cr>4�> ���«۠w��_4`�S!�y.@���=^-���m�ά��s��R��j��p�]����P@������ƅ�{����`� �{!��'�v*m<���H娡�Щ���E@:���\�͊^pFї]�a٥Eӳ/N�-j�B�Pi����h��af�D�Oz4�\|�YѺ�ln����Kp��#[ztiL�&�E��>ʌK-������_���s�I�=�4���0T9q�g^��X���7j��=��}�)@�N+U�[�0g*� �4|Q4��o�|:��L��jo�`:��ա�r���x��2(�s��W���E/��o��f},� 1ag	������3��8���^�����"�!5��D��
_�m��'n&}�B��e4�~h(��!�aAp���M�f�|�Td���������?��"y�85I���i�RI	��D�v��K� `�t�"/��1�]��x�|?q��\K_G�����!�H�u��(x�#�"�`��Ǉs$ˎ��܃�z���1�aC�Rg_0(:���#
�n ��P9�:ų���K��rM_��#k*�CF��V�|!�٣�}�4Eֆ��� �屾̄7��n�&�ǌq�4P��e���Y�Y`������T����c�?o�P�����u��?��l���5���V�em���I��
]>Ź��-B¥>�,���ZG8�����r� S��}�쫔���:J�&D�>/Q�	��?j�R�뻓�	�Dw4�^k�ͅK5㫘���]Ϭ�m~���'�u\��n���#�M�ˀC�z�����fϊ���a�d�pJ�h�ʰ#%�u)�4���V2�jmv�,��G*�Y�]۰m_u:3{��O`ZK��\����̘�Oh���N���r8��\��5�"�
�ρ9�Cq���jѰ̮]�~�nv3`�xM��L;`��T���GJq`�"2n��a�9_���[�}
�ٍW�I�R���}�x3G����M\��@� > �Il��Z)��B|�j�`��ؠ[�
�3��@,�Oj��
0Q�_@��"�4:N5�l�mөn��N�cQ��8T����o0�r �,���	��P����?1��ęJP���N�2�.�=��f�9�|�kﵬ�Ia��e�E�^�������H������� ��S
�sb�z�v�(-��t|���$
ٱxv톙�s)Ь��{;��Q7��A��:�k	.�s�[�	|ԏ/�4��M$��������
n0(W�a�lk$%-������hl`��G�u���4�AYe)4�qG ��S�=�o��fΉ�g��_�A��CwN(ͿSM�]#np����/D{�{�6"��Oj��'����}@�Xv�1�+k6q�V6���`oLN�I3��˱C��u�y Bd6Z����'��rZ�$nh�c;����;M]^��`�)��uXR�U�ٔ����I�J�����q��Q��aO����y"�ǌ1V�����]a+��pA�]�!�;��ɘ�����>�ҋc�6bi��d�E��uV��בĝ�[Htn/aa����SwsT�;�&��*bG��~�[Ȟ��t5� ��(��"���}0��� 'd=�+��[e�Le�c�U6#���FS_]�����ѧya�����	"�]F�wv6ؚ�e`]5�b#�C�L�a`c =F����X���,��"�걒�����"�_d��+_���W�8�n�;�*�����j8Ya�$��@b��I�}5�"�O4�8��ZE�fǯ��A��^~Q,T��ɐo�0���J7�s�T2{y�P�t�H�q'�b�_���K����zJ���.Rm�����U�tmD�a#i������gg%
F��#?0���������]Z��.�1"�B��2���}wm#Z�c�nz�ck+s]Ĩ��&�2��[Sw|t����iM�^ǲ�]E<t���KͨVa����=�Nr,����!�e�z��4x�v���뗆W��8���b�v���D�:��e����ռ8ВX�s+�45/������`�?R���%[eb�y`u���`0eά�ŷ��)h������ܬ��RC��U�մ2�(Q�4b�J�6{@�{O~�N� ��Hz,J���BM�y��=̙u�HPW�ޝŝ��c�+L� Z2I{��A�a��SV��-���s���3���g���Qpɯ|'��fe8�%?�ݵ�g��.Y��x��Z,�iύ����Ң�6�}Y�#�_�g<ϥ����*"y��4j3j�8u�����\r *�cX:� ��
�>j��1-��m� �21(875|�1bDk�~o�q��ZD���ow���ü ���ؘ	�mN@�ᅄ�}EK�;iyq!��ie�SM4�������v�qD��/��I|;9E�r�bHi�k���ԉB 6�2������,ߴ�CSӬ����}�[��ʥ����ﻈ�q\�r4�M����d]����g����g��ϡ���69v����!u�&T5^��{���:���%��'���B\���T��颊3��	�i���v����bn���R��d<���+���v~v��; ��{��K�������*�yP�5�(�g}��w]�����U	��rh�Rٌ��4r7\Ǚ��|�> U��5���@�^�!D#��2�b�)F���-�uh�}_$��n��|=��m�s� R��Nɕ�:*$+����Bu�g��Ge+�B-��m&��ҘŰ�Jnp�F�8>g�>G�A���>ơӚ&ӎD�J�]D�����0��z4Dt�0s�.���o�.���Hx��;=�<�*H4�%A7g���mQ�®y�`;��$9?a����T#DKH�C/��.~k�&'iY�FT&Ub�4��lH5q<v���#ڛ7��=�ð����=;���<�BZEpy��pX�wq<T�eHV�ԗ�W6wQK1D�]n��x^D� �j�t�wѵ��%�@Ӌ�sZ+��������0@��Me0=Wb-*��M�>���j��E3:͐Ь5y �n>� �&���?�0�I��[��G�i7�AUQoƓ����AŻ�����8�v9�亵뜲�`�uw�B$&e#�śUE��W��_���,r��$ӄ�u,����Fŗ(���G9_.�,�U�<l�;:���W�������|N�K(�Kl��%iJ7��;��r�,�֤���}}�$��kUN#��d��M<�Wn��Xa�-ګ�@�gL�
�j�����ٕhV�v���\W��k�Η����|��ؿ<9ƅ�eO��Ҿ0p!�A;yՉ1v�F�j�\<�c�g	G��Y�<�����B�sU20�`v}�?981�S��"8���0�O��q�u�X)�ͣB�28��o����֞���!�_�Tjetb���)I�Z�KGx��삑� �"���}蜾� /��aO�K��鏄�ͯ$���L��W&브�X\ʩ ��Ӣ� r{~�H�ft�q�ϖ!�Jg��p~2��T�I?y��U|��Ȑ�4�sI�MI����8��53e�!���Q�!eI��_ 7�Ё�_I��#���R6H�t�̲9^�8g9�5Ǳ��)�\[X�(�,�ʾ5fC���tmh�ݢ�*�k��B��������*DPѐ({jŃMt۰���Z����v��W��*�~H�d΅( +MF��s�0�$-�� ��Z�̐���Ώ���<|����^/�&�nf�ܧ�(�y��g�D#��A@Ʃ�[�Q݊�#��;���v@�}T�.1@ȯ �!��~�e=�8hT�&4��GZY%�#��v�	$׎�Vo:0�1�\��U�+,t1uq��i<�����E�`�w)ė�,O?ig�b��`z��{:�D��1���k�m���Rg,2O'/'�%�Μ��i�3���6+4j��c�'iֳ��\�u�Q`a1�2�~&}y���R�<*͑垒۞.y�����s��Ա��L�i�)[a�0[0h���Z�oᙜ�=D_G4�H�E�;�[�*�0�US%y�)�N�{9ьf��ĥ����1ȟ5n��!�"�T�8� �A��U�Do���U���'W&i��ϯ1��d�����6�G�Z���\u��962����h<����ԉG�,��ڀX!i?�,��N
�f����>/���9���E7@��\3��e!�[��ǒ��,��7>���ld:��Lz.y�N�A�}���
A�e�O����ϱ�K�)��:\'�
���)'~Z'�*�[�MS�"��%^��g��C0ZU�|�xܠuܽB��,p:-�j����9ƹ�eG[�[ۋ_0��:�U[��b-�#%���=יlV�������?�3�Y��!k��N�o���j_ �V�+�lU�� ��<��ra�}������[�L��7�6�8�_<vu���$[���|Ǆ��T]'�4��z%j?�d�{S�g�i��&�K�?t$8���_��F��fq�M���KLM�1������9�����٨�@���uE���7^�]���4�)ƀ�H�Z�G_AE�S��U�k�rv�-�;�:�v/��jaޜȢɕ��ǜ �0ޓY���}X|"N�M��V��";�����;f��s2M���nN��������;қ���?��^�,��?Xe�a=���"i���؂�N�sb >r?)��������v`t@@/c�����hY��}��%�dOr����o�o.�ҝJa�l����-0��+Z[����{��<*�Rұ�-!9oiD�	Đh�X}~I�8ӂ�b4���)lm�tE`I�Ӣ;�~ϯ�$&%�4�La��*����Lq�]r����;�0��D�`�41��ǠdkgNF��@Q�7�ш� #���ՄI4��7�{�4&?0����	���=�-�^����-����C<�s�!�p��2e��$��9��^��ܱ�Ӧ�$=��w
C4�E �*Vu�t2������c�_�8@�iS�pl�Y�O{�Č�L���z����F�$+I��:�ǻ���[i�#G������%T�F]�]�Y�W��:�2��c��=�S��׍t!��tyǧu���@��
2��O0[	)�"i@S;ɽ���L)S_����t*�B�$�cB�Ce��MBFL�u2���-��7-�l�p�!m=/�9^��QCdӪ!��m���3#���"�h	
�h�@��H2���4q뿵|��
[`�������۞��]p�����/��X��<@7�E�4�$>��s��l�p���[M�h	
-W.^O"U��=����d�Z��ͪl:�
וY����5M��ꦊ4�uL��D-G:>���|9B�{�X������g�׀3�Z���9���=��?ϱ�+/��e�iDg��Uů�N�Ɠ���NШ��{�FxKb�Q���Mʍ��
�Ą8D��;���8��-��ؐV���<,c������&c���<Pn��8b��.t�9Q�X�����c�^�mB7��]1uDy���V���E�[}��N���=G������L"vAw��4�<q�غU)���E�7^\�ϼ��xc��Ј�p��[9��p��;�({�}�u�kB</�U|
����ږH�E�K"��RNm���S���AD���WZ�ju�ʻ8���KH��%�_[��7|�g��4�O�q����Z��쇻��F��CY�Ar�q�\L�����ޠ����n�H��<�����5�	cT$i���m��ա�.u*v���F(�["[��y��`�P	.6}I�1�����bw���h��?i�V4' Vw��C�%{O�c���W3+!6*�#������Bb�&1���I�t9
N)�@ɖ#��QT��I��>�<�$I�
�JF[�ckl��F��.^���3��<4�p�	#����o�\��ð3u�k��ވ�T����Y܇���`w�_�(t<Iq��s�,� r�z����ϕ���K_
���ׯ<�	�UDb��7��ZK�E��^x�ӯV0��Ѩ(�(z�N�x��X��dr����|����H�`��-�6�������iN1����).������oVχZt�uؼo����� �#Bt��i�/=i�Rȟ��V�3��T?��-/X���-����{����<N��,X}��s������tmcb�5v?�߻��!��P�q��^�<���d����
��j�y^��Jz1Z���N���DV��.��`���_�n�mX��dry�B+�e����x��e�k�
<��H�VB��_83�+(�$��7�[T���%��J[�7�%=��igvƌ*��v��c�.���FUF��q���V��W�(z4~w�@��m �@,-��pG ��O�RN��1�5d�s�@�jk�S�o+�|U���9/��&G�1���X��O�t�&bT4�&����|A���c�������M�AODff��űh>���3�}���J?�8O�G}l�E����N�c�8��J{��g�3R>q�:�_x�2�Z�T(��z;6ž����&��<p����v+E��m�h`[�y6��Oz��D�J憯5���ѹ|p��u�@y�2�R�`�r�X$��rY;�ŗi1��~�(������E��v�q��E0�7+�����6���#�l���n�	���6���3Bu���`?��:�`���]?��|m��O�y笎_5Eg �鍈L�+���7|{��<Z�1�M9D+~���1�tD7��`D��|�4���uc#Y{Z�?-�RjC1�	3!��F�R�"�?�S����k���Q,N�j�>Э�a����q�Z��K�"���V^(�3�3 7�8a!D�
����#���M9���+�/��Ȼ��M�"���6m�-H��� ��v�@�������@O��⹆���-��l`C�� ���g�� ��9>��'�_�Y��˧���w����g2Q��"�"f�ڜJ�/ظ��+����B0�y�y�X���/-{���#4Ö���ۣh�͝�ٜ��]sS��Y�*��-�o�B�B���c����$r���?�RE�v�ɗ�4e�^;�Bܤ	�k��)x�Zc�\�����Ic,�.Zׄ(�T�i4���ڨ["b;`�&�k.Q�]�����a�|���Z�,�1%Y�I�Z����a	Yv����!)>�����Vw^P���[t@	y\[�P�I�XKO��uT��oG����_b�2�0�i��=s^-�^�7(U�����kv�>	����������$V�lIh�J����ņP{�U|9�6ٓ�7�c�X�Ldn}�j2@�����C�)Y|!R�}""/�G?R�;ѐ���� �d���x���bd��(M,`��;��(6�f���h���i���2䎟��g�UmA*�ռ긼7A�~�Vt�5���0�{2/���E������.A̢�Q�[,f�GA̝��T$���
<�����M��[ÿ�"�C����_-���^�֜��y����$���7W#z˨�kV�F��n��I)��=��Yp�!�MP����wq�lm��
�K8��Η��n�h, �C�5Oq{T&,����2��f���lN�_��T�_d!��A�P�Ņ�s��we5FC*�A?b��V�ʱ#�s"i+����Dz���҅���rB��k�$�%�:����-���D�`|��Q,�(�=ي�I&C�N��wk�mW�]G^�;x�Q�m�w�z9-K��
	�1�>�a����Q)\��[��C��振�H�� �Ww�r����r��ĕ|�I�o���a_�.�0�ގf���Ux�wx�9�4!F���&�2��"�Ʀ��	y��yęh6LZ0m���+A@���3,�W͇�)��Q���p��I�;jJ� ?vl�F�_ر�	]7���A5<׻][������O%��g��O�^Ʊ79�ԡ�:�U14F�g���;��69|XL}u��KM��E%�(d�K�:ޅ�$b�	���4t�w�NNk����v���7{�R����n3�)���JO�v�LX����������W�y=z�_n��)	�(ԅ�Ǩ`��t%o��Y�	 �M�P(����}%��,�be��4�Xi/6SZ�V߅2f>_�?�x̸��+Q��������Ӈ�4ܡ�&��r(%L)i���?�#�8�r-�h1[咕�2Ts+�Z�N�gڱˣ��륁*�LD�pF��uI/����y-���gv�e�-n�쥹|��60��2���(�o����J��Fx�	̀��.(��v��y��L\�J��i+�m���8�R�!���AV����ܙ^g�.�MD��r��@�N����d�v6*����%g��dW���*���׌��˿'a���w�P��z��D��=�Z%3��%E��L�J�rĜN�X�N�{�qʧ�%/��fL�?s�k���QC�� � ,I���S�~����>��|K���.�j�������p-WX������ ���'T�`J��Tepɠ�r�M;.������+~��9ԩ<���lh�q{�H ���J'�MH7Ƨ>��>�ͭ1��n�-��R�#*���S�z�Y��	�v�)��TSn?_& 6c �p��b.`Ͽ�CM�hf��9941��Z�9>l�n�E���N7���G�]��/��$�9#���6�af0yBح�Wn3v����ƙH�<@��]�/�%�`a�|s�ꗯ�m7p����Ɗ�X}:�)ۋ�Dg�g4'l�r� A�82���������yf(��-��5��6�"�l�%0^ڭ�]�N|��
��eՙ�K�e��/���r-n�D?]7���j`z�bS�?G O�T*Y�]�o������6�y�bF�?�.'a��
E�@�36�|F��)vFf)	�T\\�C	+�N+W�ħ�@���e\m��}�}>l���ԑ�jb_s�l���j�z�j������^����t>��Z
�N�1��� ��� O:�0��>����F��r`[��Ր����.�*�Z���C]PR�8�%��g�oo�e�Gw7a�3ꚫa��H��t���|Հf��!��%=�a�X&��,}j3I ��u^|D{�/�b]#�� ��q� �nN˕ˎkV���z�bk�('鉽�j��%IU.��D���y�F^�k�j�ۀ�b�z�Gf�	Q";�O�Q�����a���|�w@�C�g;vFol���*���T��8XWP9�rī��D.�S�'����rt�u�����)Z�s]�5&��f`�<��R��m�U��ȉ ���l����}�Ѩ�@6Lw��z߱��̀.7��iL���4Ok�o6W
ߤ)��ݡ=E��Lj0 }ub;N\�� `QvBғҬX§M�����N��!�["]�@��'H
;��c�	y�������}����4k�_���T/�F��Qj>�9�j3��"�w�W?%��C�g�����2��!����B"ß��'�W^�t�1���z���M��w��0YB�� ��і���ې�&�8��ꁟ*�%���Ȳv��!�1�`a���s���5���|tb_Q��i�7	tuk���S�t-(��)	�fC�[�-k�;ԆB������6ä�kĞ�6�2�|��=�)x8�%���O��� `���!>�E��ya�"�{������Ƕ:#r�c�jf��ɸ<��Ϛ+�clh��N�<��:����ѣN
X\y�tOvZm�R]`#2�&	%��$��z����)b"M�n��Z��$�������ϱ�iOc�t�( �J�cT�ʨ�1���?��w�ݼ����v,��t<���"b���5�PpV��{y��F�x(�t[���-sv���0��fA�$��k�u%}�B����U�+[�2��Q�:.@FH/Rp=���V9r"֎Eܻ�&�'����K�22����3��N��g���D9��4��Z�z��l/0Z�o+U���5�>\f	�7���pv�� �J>H�yWz���]�WOR� k��+5b��!Ef��<���pؔE˞%������A�>��:��_Fi@��A�z����MCG�7N���y-6|�Ҡ�B�H�sH�6U�BE�p�u�W���0�ɢ2�љ�C� @����a�u2p�ddF#���nU�9{�V:t��ç��L��{<Y�Ϻ�b�9	ڠ��f�/�|���82���u?�;Ѣ�k�_]��?e"����$��[
���1�dĦ�|;���af����#�Z������8��L�b�<��z ��M |�9�� ��<i��p󩪓o����
@��W�bA����_��Ck�g@C���܂�#�}b�������XmzG�������5E�糣��	�A����ZW=V��'߄���H�ǋq� Ԙ�,�� ӫ���kWN��%�%NO�}��pf���8���Q���f`�Z���ϱ�ou��zOEe9����S:�B@�Zx�*OA��Β��ѵO�:k&�H/�Ї��gr��__\�")�����yT�,�iO��s�ީ�@�j��Y�)�)8�K,��Cm�	*�<�K�;����!����VI�YX�R�[)-8a�%=����ӕ�����Ԣ=X�����&\C�������΁s�*�!�6��&�De éQyv��̭ �	 �b�, %��;�p_(N@�WCs�QL�i�����{��y���~���Fx@�o�9f��O߼N6,��
'Hi��j2���u����t7"����@�fW�`
�~���,�0�����c$�b�q9�;���rw˅�V��,���:�m�����㵑��u�7�R�[�u�`岈����m�V}���*��V�-I*�@5^���M����P���c�IX�	�&R�z&���(*=?�GK,� �����A$u����a<���T�T^ִ�4Fw*=��Pp�[/���[�TOt����G��YC�)$���?	������ujF	�=��@�J_�ҡJ"���-��4%�A��<�M�$�F3�YFJQN]jS[��~�c�¸�5	5�y�B�WD.8�n�?J7��T<�RY����sX!n�#��jP`�`����E1f��u~�{h�#y���Q4���������3��t���q��i2���"חx:�T�%
Wu���>�M���8�A��k� �X�� ��5���LW�.��ߖ�E�
�Ϋ�;�U�i��[v3�d���(Zt
4�>c�k��B����0�c^&�녱����/_v$;A̷�f��
+�Gs.L��f�5L0�Nj�����1�x��R���d�OK����I�?���W�@�n�N��b��p���G�z��[9Sk�~���)7��P#[��GΡ��/q�T�U[K�rf9'���Rz��
i-@��	�u4a!T�q����[`:����gVȮ��0dWm5�׶?8���\@t��e��!�����N��=m��쮁���e�s��^C�{�_'�R���ew~ϕ�< ׳)�Cա1!�ā�!�\�uC�g6��R��6���ߥ������'�-��{V4�\)}m���NPb�Ղ��xN%����E�7��mr����z�)��]3#EZPx������rG�m��-��!sʹ9p�3`zS�3K`w���������S.�n���|2)ʕ��`c���F��=A�� n;��:�F��� C�n�o�XUm�SD��2峩Vt�qj�$X�*+����3׫�N��"@`��Ǜ#��[��#�% ��;�H�j"�t��N��9n<���h�<���W֊����F2OVQQ��9����kk��|OC���K�oB�.\Մ���{���tOk�;�wV\���D�o. �*���9��i�O���t	G�!z=�
3P�P�n�����j�as�Fl���W����������P^ �@.^
`�"p�V���E��h;��GUV��I	��l}C_�@�~%�(�S������M�K�.r�a*�I�$�B[�D�ΐ�/�jU�ZC�L�����x���?���|0��:�� ��M�r�#�������u{����5��ߌG�8jMK(����HƄ���R�[p  q���	Mq���Z�s��M=E�)F�0��Śe�p����	��-V�Wn�\��)wu��54B>��_�~� `H���[[n��hw�WO��[^%�T���8侨��{��m�Xe0�m���mw��Sʋ�`<Z]��4{h�6�3Z�f@.0�[~�%����Qb�8a`�usk?��f:|�lyA��N�u�4���>��d�ǂbo� T�3#r�p\���V㈴���ʮ+��o|�0�����AwV�*_�D�z>������m�4�h)[ќ�7fNϡ�eck։'WR<�x��4n4�]ؿEs���pJ-(���4��nOpU
W*_}%n��r�2��/��zi�RY@�	Qf�+U�������P~�}�0f��1`�|0�%���Z�ʩ	zB�-h�ڰ�ez�'��Lp�N .v6ǟ�&�)�,/!���N���Y(���n�(�C�o~��f��>y��#���FV�{�{_Q��f6�s�S�yi�_��1c��}b�.�~�l���H�}k����3���Kk�i��y�Ήz2�s�q]�d�/�q�9�h<�r������R�ж��_�X�w[7*��$��=������>֒:��r��u����AA�GE��TV�Ep��c�ʚo�ү�	4�M��#��D�{�jd8��u	���^�+��p���8��8+���k�����_�Kf����a*�,�����]�}C��3_�Z)���
��'��v���)�Ҭsʙ����Id�&0���E%܍%1�R����Iꕖ�Yʃvw����V$Y�3�=r���}k�"	�Jc0�|/N��8ֳ���(@���X�`r
�t��aċ��=O�*v���>��o[�/�y�
�#�2}�������OKӸ4y��|n������9��Gt`	�FNʢ^��b��8��YrDl0@��nʌ<�9�k��&�J�T�댻p����|��7(�����;D�8 ��N�ĳ!1�JaI#��S���ߚ�$r�T�ù�9TzS��3�3�����q�6�aV�q���J�Z��R��m��l]�����|���fYN2O���{��M~3~q���,Rd����c�J�L��?� h=!ɤe�usC��s���*���F�Iw{L?i������7�L��A=�����ݒM���;���2�=�
=��-eC=��HW�OFVq홆&q'L���<,_�W<0շU-�Q��JA�[�lv	��Z{��E���$��@��R������)й��(1��0�#Y8i����.ޓ(�t���EfO�!Q���S�I�t�CA\`�n��u���mr�F� ���<�TVV �v(:�1���ϔ	L��P6RL���a2�J7����E��o�Wnn��"K��m0D��8�1��V���V9{e6h6ɇ����NSNp�ެ�!fᡡ��43��%q��*��V�Sue�֔�)L�;��4�G�i��PP�a�#�ũ�F�m@��㬭���{���U֖>��|Ҷ�j�K�c{獬��Е�[�@'9Iq��g��� =N�7�G�z��L}M�Z�k�s��f���S�	��z���D m�U�rC}2�)��O��3=��,:7婑��HL^��j��1�I����Mu4Y�e��[����=3�g��~����zp��#X��&ǰL��r+$h͓��*f��I<��}�Gg����wysAk_7���N�k1iR]�P�[�ަ6�?[:�J��<x������J�jG��L��u�ݺ�b�t���u����fм������d�=���g|��t�/�M=ܩ|��7��lh����c��p����G�3�){]�0����T� xb�/�/�%��(o pͿ\|&�����!�*sqɤ���D�6P��֢&>z�D,
���B4�ٞ��VI�ե��b�!�t��H�Nk7�,���YV0}}�g���oE�&n�6��-�gO|�4&*�؀p�k�~7��s�1,tW|����ZJ#�����U5d�����uۭ���G��I����5t��҅Ix��J,�8���5�}室�<�O�D`�Tx�Y[���fgi�å(�U����Dx��� ����hĒx'�i�rd�'�̻56/�f��?h�
y��� �#U��1Q���`�Oߠ�&
/�����j��ƶ�O�}\�x��trD�����Br(� �n��ԁ�i`*,�,���M���Z[�:�X%y	c-��F��:�(,���Q$=o�;:���[@κ���
Yz�,�n!)8���H	㤮�@�	�O����{�MM�
��Â�#G�Ʀ1X�8�Ba�b9�#����I����\>�KTq�6��l��p�A4��T[� ���?��k�^v"�4�E�P����8
/  ���E�`�3�+S& ��,�:�{�<��x���C��+������o�$���R�̥Mf~�d�O���2�O;�pΡ��' �����]M�W��ۊaY?����ҳvD�J�P��J�	�%X咳�s�|EvCV?�	�kmB�xfK}N��B
�㹞T�6���|���v�a)�Uk ���ւ~C �P�$>�֛/�a���9�Jq#5�jX��>�h�m����]IX�X��N�F<(�_$U�<���wm��abگ��t}HW��h�(�
�3<��3�K������Ǫ��2����{�@N }O�3���5\���p�ђ���PA��?����s��5A�Md��o��q<���Ћ�,\�h4ݥ���
u"��Z7��|:#��$�nC�Xy�<5�ۅG�7".�q������e���s����H��9�(��4H�j��¹����L�r	FD��<S��M1���3�sB�d���;+6I.¦�R��~��^L$�5���A`���:�V^Ue)M���j�nz �c�)<mk���K�vb���O7]HPU�����3�G��3(���u&���N}�Sy
���Xs�L����V��â!I����[@�>;��^[��۴��%J�כ������b35iC�D�_vx]/����w��o|��C��S�t���KC����u���l�ݐ�d�5YZ�b��g��I�*����(��l-V�N�6"i.���r�����p#�čhܘ��/YC������<N�f���߸lG&���X����i	���z�d�~��oa0���JDg�WƗ�UL'����鸞��|��%��h��{����4_������=*�	�+^+Oŭq��6���l������^��s�6a&+J��;<�QD�~�*}A8�Y�6lE�q+zd���6���H���g Ezw�@� ���ІSz(�)�p�	���8}���B�*��!����Y;�)D3�Gx<��h��T���b~�|>�B9�T�Ɋ�9@���tiM��^��%���Zp��*����Hl�c�	�ާ<[:�GG�NLZ�jj���Qq��c'��:��,x��̻�#X]zM�}Ec-��O3y��̟�'QG��t�͂����Q��$�O&�����߅oD9fO1�t�\�^|X���s�Lm�գ��Q�}|5� e�Xd�f}�6DTni����)�����Z�Y&��F�?���#��j�����~���v�&���I�!^�和=`m�Շ������тr�����I����U7֪&8���e�)[�p�U�1��wf?��g�D��_Ro�oV�TE�nͮ�Y5vA�����NA�m��1�w4��FT�@l�.!�
s���[�E�*�
�xS|��18޸�8���R��PRTq?S�n��56ù;�KQk���:��N30tfț,bL�/��?AMb��1�臤ՃN�l�Pw�Պ`Ҍ�#�fe�غ0���;<d�e-YA�>s���Êf.�V�t�#�	�v�uYm4�0�\I�F��$Bl1:�\'
_#��Q�����|m�6t�_�P@Nkb���KAy�(�����~��i�T�:��9g24
��R�Dr��(�Q;����l�?�-���.�.A��[�Oeq���q.*��p/}�v6b�r�0��!�5�9���E@5�C�[���'pw5�}��K�Q�����,<��������+F�Z0��1�J%BO���XD��a�ݮ��*�KuYc��vY
�䀉or�f�ʰDŎc�1�����As��dy=�5fۓ��oZ�����E۩:�g����׹q��o�{��$0��X�/�(��u��C������N36�Ͷ5`�@ڮ|y�����88)����d!���ցv��x����Ӹu]����u�l�σ�G7�[����{޽Ŧ�ʁѕ4�".��'5��f섥>�+�ǡ?ˠQb�|3:�9�M����Ѓ�$k�"~�)���-}���?�/��l�V�7&���		%�r�[[h	S�0' 9�4P�h"F�E3������㸈�$�s���d.��q2ۻ����jx�.�
���F`�,�g�ϖ�iß:�Nk<�>R,7&tjL��{������LN��7�=����N���._y㸅��_��5*C��7��U͘�Rv2�Ot�@g��x�j��������u��-9s�|����,W|0��a����[�3���CtZ�g���_�ЅJz��?����i�����[^�=�Hc%�n��������n���e��K��ww��{���e��5'�h�E�y��f�ԅ���(R�ƺ�r��.�2�1�۱O�)�Xwg;Ǣ���O
�vk�қ�����\�As(������o�d�^Or\tn}�hy�t���| �<����`ܮ� �"~�m�֜(_.k43��jL�γM�*���؅�0�Ik
��)^:˸�*�A� q.=Kx����-�keO��݃_�c�/�ڏ����}�O�ds`���u@��zD�@L4 yi)���[�ȓGu���nݑ�S4F��4��!���h�b6f
�-b�ϓ&K�}�9� n��za�Q��j�T���g�#-���a�傡�,9/ �Oc+t��GZ��c��L��������RQ#��3�Sz���f/B7 ��#�����/�ee<S�)�%�9��S���`�$!2����n�=^=��$�$֗�z���s�B��(CS��Y8��ζ	.̡.-����Q�ϜY
�{&O�V����ȩ)�N�+r��s�wV7���ndn��Q*}�Z�k|7Գ���@gw�}�����#��+W]���'�ϱ��z�.�Jm��2��5u��=��7��鳗?$]�}P�Iwl�;���6��ԘM@ �]��t��M��sN��0��%pq�����A�/%6�`�n�������3�č32�,���@'������2�������N��ZCw��[+h%��������b��|��k\g����{���e� ���R�ay��
ݒ�J�7�<,D�KI�6�ͯ���#	0(`��kd� �ģ�7"}�(�+��[g��eh�C��B�g��r�vq�B�B�i'��>��d�>kv4��y}�b"�%����k�8���'�2�[���f/`���P`$���~�/�;,��T(# �Ss�p��!�L{�˧�xUȃ�XQE��Y�*Jw�؁�3��8�V��t����Q���隬u�=X�L 3��x�;�������}���S���_-�1�FL]Յ��n����E_�������:����!�_�5�;z�U;��~��+&�y>L�%bֳ%ڦ�J��^Օw�7}gT���C��+��N����'�3y� �*)�ȈNI���o�C���j,1  _sZ�#1
���wI�)�"�^LH����%j�]��{�F�^�E0��cOșFk�Ix��]�K����u�M8�����f��:��իq�m�]��9��_�E�OU?ˇ�m'�T?��T �'o=�q"5Π��6�\�P���R����Jz�ٞ�Bk��|���?���n�e.~1D���}�]�3�I�md�q�i��|�\���ɹM�?nZ���t��em	�gY���^a���v�K4J�@��xc��B��[���oᕌ���}�����g����p@va}��
�S�
�a�=��7{`��V�q������D�n�嗐
�_R@^<���'7��-�>���h���\d(��7��?;��c��О�]ú
G$���I����Q��|��=ʥa�����`��k|�}��y��f��Э�ԇ��OSkh���
��Bu��Δ���wf�r��,*j-j�0_/ٌ=�A�q���U �"8���?���;5L��[�;	V	�ELFÀU^77�m����{2�6���H��8��y��"�S�O��	n�x~T���uK�x����H��
�ny�#G(>$0���N�����\Cm�
��J������U.�{�����?/q���~	���v���mR�y�Bd��ˀx��i4Э^��=���a�<N'�K76����I/��h����m3	Z:W��$��c�"3��o&P�dZx�9�e�o�^��_(��*JAHK#����5[/9���+͘
*�����f!��#������y�Z�2<.�D���8�$|�s�}�g�C�0����.!3�9����o"�k��uPG����b�I#7Xz���[OF���S�����!�b+4�%2娡l�Du$[���<�(W�J�.P�>tC�5�` m�3`����l' 8/O8իR�=\�a#��������K�#y*�	��N�w�ɯ�`�R�H$���,]���L�D�L��*m�?�[xg�hX(���Ꜣ�� 6m���A��w��+|�OW59�W����c-QRQ��5Xf�J0���,�si 8��%��������E��m=gAr���n.��E�|�.���Yjd�RX�mVfw�S|Ƽ������D�vM���4�I[��G*�M aA���#y+�9v�S��JG�@OCT�k�����V��l��y�OͧD�	�*/����:����x��!A��?\ԍ�����1)@���p�J�-j��(�g��I[���4�qPY�ao)���ڿ8r{�*� ��.j�DJ�SK7!��Ic����3��@)�#���v��(s�;���r��7�He�ӕC�A��Ic2.b �����3P�2Px������x��mݷ%\����U�;�	?fV��6/��A�� �����>'+}baذ�zH!�m�
����Y��%�|Vj��8 [F'K7[���9����.�WW�5��p���JWgg��]��e)�7���t>F��|�V�pȭ}�Ju���Gb/���R$m��d�lԗF���z�^�t�S���1bvә]�ǐ�M��<tDl�4us�N�'�v�2Kl�V�#�9�ƺS�n�TΆ�	uO��⩁��w��_�DP�)p�������ٚ�����X��4��7��;;�0G~��!�g_�!���]m��â	Sھ7F�\�c�sce	��Z["��������G�'OOǗ�����T!�����v���Qz���=`$+��괂�m	�L��~��H�}�9	�mLb��y$�˅hʓ
��H��͕NL]$>��6�g���򳍙�-��t}��л���N	j���`���C�0��N����E�H�z]�'?��-�a���#X��{zcW6��/��=�A,
��m�!쫙cZT���C=J���D~]D�cU��6�UE`ڱE���_��Ztr �P:��Ճ�vC�O��;����v��� ��6(/ 6�]��j\��-��%��Uz�(�x�ӎB�/UTY�����}�Yl}�x�����܅�NjT#v�O�CW��<#i�g2�բ�8��겑x���[�V��/�U��Wz�u�0��ʚ�f�ǡ�<�<�/�6��o~ܩ6�4�nF����� ���Y��E�T��G��_�ZX�c)]}L��w�;�`��7�!wou��9p��1ܣkG�XGX�mfx�+�Q�-�y!��NF�d��d���\�'uO(E'g�<��k��Жtm��S��;)tm����[��W̮ƃ�
f���)�2�`��KĤ{��m�9!]:+�~L�M�Qh�hb���0��b��N6}�6�~�4�����;�W�P�?/��U��_����!�p�r٦��wd:u'g�W�!�7�6[E��\*�ԭ�5t�U��(���R#��*��:���w��`([�����w_a)�A��-uR8ђ�n>�K7Xy�\��MB�+[Ք]c�WrY��S���(;Ay��r�ivld�+윇Kg�z��U¼_�L��#�š�qq봆�|}����M��k	��[]\.��"¥c�t^SQi�}~�*y&O�'�0�G�>5�7������ev�"�j��aG�-
J'�@�Q�d�_ծ��O��g����nO����.��p������\ r��tC��Z;�\�.�7s/�����x���z����E􋌕��!w��ޞ�u�S���k�`��q������c����Q�\h
%9ldǒ6Tv�߱�w��-��(tFDk}Q�I9DY���Ha�FZ������^�В���79�H 6^�$ɛ��d�w��D�	��a(�ނ���L�[լ�I�.��>~5�Q���Ĉ}F\p/���,���<ZrJEXAq�o��Ⱦ2	�?"��#�:��B�Ǌe�Dԥ������4�W�ߎ+jBM���J���Oec8ƺ��;���P:�ф�Ӹ��l9���3�ێڑ�+h^��.u��⸇�sE�������zA�L�[�Fɂ/
��Z?V��9׌�ARv�j'����B��RA��>{�i�����88-Ǩ��.�pL� �`��3IUl�Bƴ��
_�q�6f��Q�:�-8JV�c�<�ݲ��Ŭυ�.	�4�� �k'a�S�q���l5���i?|��V�ʑ��[���y�w����vL�;,M��(/V+.��z��e3ţ�G����r�=�.�вu!T�PZ7�-��k�K7���P�S��&\�[÷X�B��:۽|E�8��N��<�CO��j�W%ڹڪl�YLlT`no��ޝ���Eŏ�";�j����mɆ?�H�yj�HY�~D���q�}��*�Me�I�|?���P�)s���R����Jyx�
��[����Q�{�q%Uk�<�"\�08��c(��L�}JG~S�<�(i�
���S��W�Sħ�8�
ݠ|#6��W��tlf��ǣd�?���>ٻ"]�9g���s�{j�B���E����5^��E=ғ
�23I�_��_qZq�$�?QB?SZ��R�dVh�>��� �s �BIڹ�̛��>����E�[@;�iP�����'w��X�ZUpˤd�ޤ�6P�F���4ϊb�-�z�nL%e�4�IR�n�J^�R�z�~��n9vg�	���*���V>����'L�Gl��CɎ`��~�hy��ڠ3}]u�C��qS:�P�e8�XwN-���!I;�TV��.�[ǢeԞ^��|$!r;�lX�ݛ��*m�}���� MK��I_�#4(�ES
��'�=Z��!�c 6N};�$w���wi~�eR�"]l��|�Q����I�'���Mc��$�b��N�DyᇳV��2kd���<Ss�%!s�s�s�����閳��v��2�g�a�S��M����2��9W�hSQie��+-�����p�:�>�#|<#�@ۯ/�7>�
_���n���}�2��q�2��X��j�`HQ
�P7�	}��A�������^����FC���n�T)>��)�f�m��0:���_V#���c�i�J�(�Z���̒uP��*�d!�$�ڠSZⁱ�;'�s�X�{��j2�q��ҫ�~ˮĪ��s�!��;�(-�F��'���>��%M�h�VݚV�K��dᗣ��n�����
�Ϗ�,!9��i$I��>Բ��(����qt��1_��x0��a��<Z��v=,��qw��35dɻa@h;*��wڬ�h�X�-ty.&y�:�s�y9���X���.�i��g�'������ �f�H(}�~V�V�/Y�%�$�h�g�07,/�=[��ӮN��x�qf�묾�*�Thu��yf���^N�wk��`��ϸ,Y�$ϴό�W��.f-Mfk����
�hV�,y��ʶ��� <h~M��Ͱ�5�S߳�1vO�>N%�O�	Tj(���\�N|���hˤ Bn�p�p����G��6���͚�1n�h��1 1�I6�ԥ�����f4�㰃���]�������'!0�����6�5��8�#�Ă|�-����T�`��ՍU&Qc��xNJ��u���Á%s�����>A$��'�#�9� ���I��ߨ��1�P��z�|@�.�M�F�J���Gt��,t`x�Z��VF5&���^ۍv��޲��r��^�kgY"���5�b�.iQ��n�gJFЎ�
��F߶��#̰�H�PbZ$�m�z�cJ�z:���t�O�S� -�Y������D�[�����̛ gEaB���mq�����)EE<�r�Y������Nn���zK.�6�[�0Z�{\7���^}fc��&o"�_@&\���PT*��[ENY>mx�q�M�sM�^���'{�V�,�|_������@� �G^��u�:�sLQ��Ab��5�&���6�R�_χ8G(��߱xu5��+�mx�M��U�j�/�f
����x�����Z3�,��+���U2�"��ml���m�y�����f~Am���OR��` �9�쫱�9}V*� �Ƥ��O~��Rh�W����?'G�8q���� ��!pe;o���Ɛf,���!^��1���>�㖼��0�v�-E�I���?�}6DU��T�E]~L�߇l�l� ��t�O���&W/^�9�r���C�-W��l�<����5� ��z����*�ׂ�4~��g�վ�5�=�����w/���5qt׵����Xk��>��!m�����.�����"�gM��Z< ��}�C��1������;%���*���&�@�����OH��{1�&p��Cy�r��J���e���cd��mj�х'q�E��R�;b���Ő�B�-���Y
ƹ�@��;_zå�!I�����rr�7S�j�V���4O+V�3��P3
�;j\����<ލ7h~�f?���Y���_6�~
^������J@C�;3�V�L���߷�"�����*�V��6i�D�\`S����x��*c8��:��˓�G��7�5A�.��<)�dUBM8�dx�ǥ��{Dm�j��anYG�t+Ȳ��{[�`����Av���d-��V�U���޲%I7��>�e�����OB9���*ʊꗌ�5�`�Д)&���|13��V������z�M��,��b)&�/��cl��2�ߗ/�26M�Y�jW�l�׹2Mr��5(b��]��t�Q�XJ�Kd��5`)m���E���V��Zd�wA��uь�j�.�}8jJ�_���\���pE�o�b3�i?�V���NDk�}ln�r���nWy�"	}���!	R9/tu�I'mΘ�F0�=G,h������=��e����&?���o�6��}�H�x�;�q�:<�m�L�;�bw�g��x�~����8�4�6 ���;�����t\~LGc�z��f�&���u�+��[�i3+�l���k��':�]���h��e���G?�U ��i��h��ؼ(\-�Y *-wGS�uX�/�l+X[0]V)ڹ-@a	o�[ m�9���_cD�;� `(ƛ�4M���T�v��޻B�+<'̫��'bS(�m�`E���)���J��w;Aݭ��!_��yő�>-�\r0����(�c>��v��g��%3�6�l %�b��ãtm2q5>v^�:�ҝ�'�ɖ�|L,��	�/��(Q����ߎ��)�fgN�� �v�+�=,��otC��?�Ftj��S����f�o�z/@�0'E�5�|�\V������85�:X��D �)\�ԧ����,5D�5��^>j�@�_ߏ���%`_������s��|4��-,,����=F6l�{f��5*j{�F��>�����'8�S2]3"�2yÉ�6o����	��9+��#-p⋚�G_M�c����t�FϹѹ�G�i;�o� ֶHR�ǵ @d;YKt!�|�$2e���x��q�<wW�x,�++J5��`,�J���K�G���W� 0t��$Τ�������t�fi���!t��c����]Du^lњ'��o��=WN�0���{$GJ�#�5�+e�}��(�Gk_�U����H���Tc�WR�����G��H0ev��b�<�[��gUC�^�_�m.�2�4`����G׃��TK%�TvlvF�}��q4@K��a���/h*. ���Z���c�~�?��ϘC������/��ܯL'���
���8拊��}ݑO���k>���*�Dҵ�2�9Q�͉��[��	���k���(l�Ὑ�Tj"��#E��B��r!()�qصQuw�]^�M��*�W�ޓ���.a�+���y(*tW�"?H��!| ܁���%�b�}��_���!��yw gd� &S�K$�sϫې�߱�ӉW�w� O��.��<o���9��')/;�� 1=�Up���lu�W�i�(�7-��)��Z�mІ���ڳ��3�Fˆ��W���&�}m���5|�۠�
�*�w~���P[;j0�����826.�ő�Ac�3��Q|�;���Oz�4���4�C��Q�X_���b��Q��)�Bl4���W\�\�Z��ed:^��IY�H�&��I�IP�~������B|G�	b��铮M�����Mr�<��fƚ5DDt8aI Ժ�9|�	�S�/�k�cG�o�����w*� ��'�O
�q�Qy�S|I�܅�KM��Ne(?�n/�m?!�/�hZ/�d��t:%����B 
����Lý"C�K�Z�c�N�~bX9�����I�>|?ٔ�<:�[���c�}�SrʗZ��?�$��ٯ�H��VHq{B`�-�M�r�e�!�,Ug��zч
��d��YФ`j�� *�TTC��&��R'	�p^�< 8�/@L�W��a��q��#���^�.�G�5�IY��0��Sꉘ��L�������b�+�V��w���?��d�r.�N�,��[r�d��t�jx���u�x[�em �Զ�^�S�p��p������ĨK���q�ؤ��5��N�-��'E���J���#¯7V��0���>�n���9��t�kL4��(\��e��&�4,� ���8Zo3�6�؉d�YF[�(�b�Ӽ+�l�\ȕ�l���v��ϣ:�D�R��.��i�r暭�5�z�s��A*�2��_���G�'/7.�pN��ԩt��d��G�7[����Km �\��� 
Y�}�C�⛸#�nZ�(o��)�OFcW�+�������������?ü��	n��q{٘�r9���ٗr��ow�vk����f����!���ʁ>q�O�_Y��Ǟ����$v%#�GB�����A��#��1�A�6��3]*�={s��(�fVDxx�jP�2���'� I$Yto�e�Z^neD:����-L�?,���U.�X mY݀YO�vi�R/g�O�u�6�ؾ��Vs��m�9 �j�h)�H�F�3���`N��b��>�"2�cG��x*葜5�m0�Ń����j�o�M.MI�����+D�E�����]��H�f�'�@`�_!ןKD��':d�Ė�oFxg��D��oq/�܊�v�<����yY厊���뿮�
ٜ�d�Ņ�u�dk�:"��G�W�R��"�f��u�o�ҭߎ��u�1ҭ���>$�H��b..3�l��_�q��#�������/��A�M,���˰����;�{<��J�<����U��eò�_혷uƫ_��]\닝����|#��1W}�:��ѝ䗎0��b"Q<���Xf	vχ��ٵO����oͪd��灮���U�K�~H�ixRŨ()���̱;�(q޲~RQe�@ ������1q���6�7p���.�� 9�G5?�ڎ���kB�h��f����*���)7	�����uf�2H�M��T͜�
���x��ڝ;"���ֿ�!�	�"s"�AY��U���mji]ō$�4B�?|�����TS ����&��E��b���*9>+лFB�:�gT�"�r]��^Lj(�r��{�u�Z+9Q��B�ق��\X��{��"
��>��=,�?HI�3}=;n��A@��ޘ���� 	s'�s6�'�-3:a�~i����$Cuѡ�*�\�QI������7��D���U��a݃��M��C��`f��_����F���	!�pH�6���?T�Q���E.h*lꖕn��ųcwa�g2��;T�<ˇU��o4WA#z�,��`W����+>,[p�3&��\*���w����u����J����7�H�j��ii��#���ؙϽ$�2�֮�X�4��્�A*�dv8�NTb��O�����^;����Yz�=A��㡝yb��k��F�:�@��o\րi#%����=q��jF3�����g �zR$��i��Hqӥ9���U���+�����p�f�J�x��c�z�~�E�vT���J��ڌE��^�JZ��AA~�Q"�a, �R�NH~�1bu�V.5o��K٠܋)���oՈ�2u��R��l�U��_��+}�da����IY�*J4�}�j(�1�����<�z6d�Ya.�Κ���kw03g����r(B'���1�M�.5��t���1�8�M�0��V|�2��8��Z�!�d�=�ߦU�W��ha�g'+�Հ����H��ȃgc��C��Il���[��2�w�ݾ	��M���DFh.w~G\�Bn�iL�%�	�w����U���O�I������as⃏�����lk�\��{k*��DD-x�����.$vA:��k��qy��i�� +_�Vt��j��{�� ��aK�LJ�d���nOV���(��=����kh�J��#�43�7����SB6���W��UH�H�43���a\�8�Z�uRY������%�5w�Ӑ
Pj��h�\M+�"�2� �./厶�Y24<+�c�!��ؔ����ޤ�k�7B�f�,����)N��}���b�u��-�ջ��0���� �t��ݩB=*r��
	5ӻVj[)�o����m���j{S�w�����J���or�[\�.���sA���ҫ�P���������G��mM���r�BH��!�[W,b���Э6���񡚼����TO��l3r�4�Rf.˧�;&����x0B>q{�����d�����g��Mb��ڇry�{U�6�w$\e����U�T��m(sέ�W����F	H�N=���\U%��>�uz/�����s=���ʳ`zI�a��Qw���ĩ&���<��]���ߐs�?ǎ���2�Q6�=`ply�&ƴ�mҹc�ǘ0�,"�k��u&ic�+��ڊ�����f�Y�5��%Ś^��Leŭ��d-�B�� ��̩������Mnx[{?f?\���NQ�;�'�V�l�����g�=|z�5b��C��W�z�>���%M&�B��]�]�2�sM��A�H��5h�,�b���P,�>R�l���x��#���m�FV)��m@9�47�x�¤e)�d�&纵��J^�_���LxX��륕��\�� �H��"��5�j�av}3tCh�Tc�x����Ժ$���i� ��2���v�)�,�@�غ/)��9�\���"���ҕlFQ��>�H7ã'������
�]���h�"�_��t�S�G�-�È���t��lɕ�im#��Q�-nE���nP��M�x�g�g���,19*A|��.�2�g���0���,�Ʌ���|��l��}�Rzb�j�ErP;�Ӥ�frht�����F�z��W���M�_r�������9��ۊt'q�a^�lJ�O��v��.(�������"`DYk�cR���^`+,�zTD�5R��� �̳zWȑU��\s��UD��$�Y}�$�8��f������zO7#<�R�+�J�-+�E��"v~��'���1��ٟ	��<� ��i�������@���n�;5-e��� ���5|*c�	ء��'-\��	�kk6Yxa�a����n"	{*�u|;?���{S�Hދ�T-����|��6k��}�,�c�wk�Gv�C1�R܄q�-3���I�ݱ���,����Z�����B$�E���I�7�����`��D� cD�$�(V��0pe�P�erš	D3	�Q-�-������sq��H�ȲW�A�n1$�O�r.��=�c0�����������D�Xi�L�!�h�so�%����)"d㖧����⥫���ͦ��ՓN��>~���&��;g��#9�������FZc���l�nY�FrV�D�P��Ɂ|twg�&e-I��U�r
-f�RE^��E�+΢@\����� w4 �L^L9$�r�S��/3��Ȧ���>�P]͋K__�4@��pi�SbJ�Z��+.->�L@�n�J`7�X+n��:��u���E�ʅ��T{��W���+޸�{^�Єޙ�Z߁�!L�}�'�UrZ�ܡ4_� ��$��������guQ��𰉏�~A��E�� ��G㒅cd� Da�8
�n6���-C�����["P��+T���E�
Bܫ�jX��v��})��؈�H(��Rd:���Nq������*y"�����%EޯC������ �.D�b~¾�����\PHw8�gq9��&F;F%����I������ڄ�hCz{i����������^��{��%j�kybp4��Iu����?�������jJf�.-L;d�z�:����1��x��Kʙ=$?��W��/�<�,�&��,s�?�l��A:!�7��f�������'N�fܟ�ţ
GK���:r,��2-�ߡ���,r�:���ú�$�۫�ϋ� ���v��H ����}�� d�Q�9�,�z<�!��I"�b>�B����th㔱�|��o����)u���ܵ���P	P�j.��U$$��t8�w�qw�ϓ�͜��	��.���h��i�뢃 �m� ]ٗP(���Z�p�`o�q'�QY�l�9�<�۬W栟�� ��H�4xȄ?*�i'�Ɠ��^�����f.�1���j��\W��Û�=S��-'���Uǋ��ia�pQF��:�Xj �va׏���g�m�����؆"�B2A��v�Q� @�]�n����G�3��c3�+� �	&�<:�8@��n�",r�%;n0 4�8Y9��s��`]gg-����,	��|���^�G�3z��zC6W�~��&A��C�g
Y6.�_)�Kg^L�Y�Ϙ�����F��a��pkI�9�����ᢔd���铏���ԫ�������x�g�c�r%���wR��"�֭ˉ�iV�%���b{�J�C�����#����.�w�f�va��i�g�#kٙ��R�0�ǏA��}v��m�u�jY�6��"��*!o�׈���Os��M�����"���/��M1��?k�r+,m�A5��8�w�	���ܟނG����+;��xdӴ��ޚ�vZp(P�<<h3.]���B�4I%С���h���m?���TZ&#��k<Y���R��Vy|	]��<�:�r찬{ꎟn����h��� ~Ғ�������rU~��W���𚁙l�Sb�y��^5�s�i�5iR��*�.oe�*F���2��G�k/�#b;<��>D3���`l�P�u30,��%VBJ�WwgW��B.9�{=½�h�:�m��'������;�.?�q�������'���"z�π/!.�h_��ha�nx|6hJ�D{�.B�#�u���37T�	�Lo�V���,��0�(ɢx#k,ڍշ�<�?��o\|�>����&��,3�0p��4�?����BEʲѶ�!���nw����E���IX}����cX��{�%HDp���ذÎ�(���f*S�.����I�Z�՗e��A3		:Iw�!�X�"��̦ZP�'{�D����`X���ǆ�C�e��r�0GφL�zrR[�H�ج�j��&+}2�q5W��F�Q�t��c��-K�,�X�}�n��V-e)L�O��ϧ���&�팇%�!?K������� s3��F��=Q%� ^���0d�4�nN+v�*9��#�QT��Eurq�|���ץ*�9�u%��Ȓ?���%%=�n�;:��̅=f�cB�h0Vrb�30@�z�(���4�2md�hw���+��i��@��;�$v'NK8G��vĵ�e����o.����-4c�(�>{�o�2>���@@�z $X����ʱuWi'�ܴ+��z��4+FU���=	���Ẑ-�2�����P$��ν�?������L��qV��m���=�G!���j@ީ�&1��"�U&�(6M5-��y�}���? �^7��Ԫ:�+��c:�"g����E�+S�h�.���O��a9��7�~8ch�_,�'Vu�>!)�xc��,{��ۺԲ�� ��R1�6��6I�*�Pm��_���C�E