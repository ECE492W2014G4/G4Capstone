��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�"��F9s�`&���a�oq���F�g�O�]�<ݲ����eCL��D���{�5��8̝DFI��Zp\m|Q��
�}�6C���UnF:<�jΈ�2�����<����sf�k��,jڙ�����2��X��Ss�HL��	�������+g?���N�Ż�����|�v7�{M��VNB
��Rs�゙�Ld\��X�'��R :�J���^�����kMkx�Q���3!P}�e���Z�Y?.�U{�RP	�)��lI{tI(S
7ZF�����O)(}��b�֡�.㒂DF}�[��]���	�]y.^��`.jh̬xUQT��`��¡w� Kb�+7[c�h�R̟R�͖��Zw驼���X�t�[�&�����J��Y7D�ˮ��v�\�j��r3s~�i����r3p9!j{2{��F|e�Rb�p]"����ƳG����q���u����W�Qa�v}�ݗ��k"�O M����][��w@��WX?���m� �~ S���+� �"���B���m����m�R�Ti�r�^��R�-a���4�6m�rg�����e~&��$�=���L��^��V�u�Z�o�����&��d����he����]G�r�4F�\u�x�������s��f>�#r��5F�����pX����=J��b5������۪��$�l���G�4����"�f�^;2�s������ߓ�QZ�������x%��h�$�s��M�Z[�)�^�t۬���'H��sg@I�p��h���9�U)]�]~���d�'AʘP��Z�I<�u$��
I����X�ƹ*O��#{g���.埻��&|�':�C���x)���Ƅ!������i
 ���~�[��xO]dlC/V�f!>?���Q�A�v�>Z��˔����LϜ�ox�l�zf�f��x'��WsC�I�����b�M��DMu8W�ƞ�\�����8�$������z��B��AM����/�$�ࣷkDt�Z��o���Ռ���Y����/��w�Bx,�M�##8�(R�	�,ëml܄/�na�����L�,�`�!#��:�E��ef6����@bR~�0d�}'����-4�׀��R�lX{��a<nw��!�T4����#���f�8�=�o�#2��h�)���\[�"8 �D>����D��r/�ʢ�0�����yl�.�#M2�S �47����_'��Z��Ԇ9#fo0s�sKB�̫[��$��k;�g�R.��s2tm��r@�u�q�������ݮ�6�(,��Sb�f�'.�|g����F�C�[Q�0�{"ǒtq�0����&�k�w�ϱ��b�Uy`@��K�^�6}J��cZHfO� ��of~�ѷg��%y����|�M@�l7�K4n��CI�8|6* қ8f&��.�B$C� ����ss�A��E����)\���a?.��Q
�W�p�{(���� �������{���(�y����1�2؊1	�_f~^0���g1��-�g���[<=�
���-$��f��:� �x�Io$^����޶G�U@0�Vښ1��#���e:�D=�)����!Pb��Pȫ�k��`�Ar�>pಘ�?����[���M0�į= ���G4'�iW&�B�����+�20��_����P��l�;�
x��Q����0��mb�Ć�Q�-�E@ߊ�F��,��oK����UZr8�P�W��d�P����Bb��Xڔ���B���$� Зs�}�u��c
Qr޳�(p#�qv⦜A,��O��|�l�i���>~zh��}8����w��b���S�/��%t��d~���b�I٢��%�st�3��غ�8�����#�;nv?�[>�2���Jk�a~x�[���>�^b.P���$~"g�}�#������"�8����i�YH�-y/�kdE�IoARP�_�U�O �C�!��;!c���^���v4N����m��t�x.>.j�-�)�� 0*��2@��8��E��~�f3�֌���!"�E�<�
d��|�{`�-wxU�#��>�l>>A����>�l�¢myG��l�u�7��	z��g��v�(/�Cl2�nV�qw��F^����
"u7�����ؾ�	p@2���=���jE	9�4τ�#&]��GZ/�ۂ*x��L&���7�([F�M��n�'�?�˺^b�>���Şp�ic{rꠓO}��-]���^���l-��N��|�0㜡feb�	K�t���"��\���u�����O�>��&b��w���2���G�a	�e�VbT)�y�m3MA|�� >���9G�Ӭ�q�w��f�=~l��]-^��\�N��lvo��#�H��j�(9��_3��Sxƹ�}�ݕ\�K�}Z(�{���M�R��9ه�0����Z�KT)6#'����0n8��S�g33�S�tŞ2��4�t��S�,.�R
�	�S���+�����!��˘ƴ����6��T����sӃ���	ѡc�-��n��Ϣ=�N�4�b���ղM���xZ{mlOGߖX.�t[HB�G���R�M-�sth藄�TD��6?�D`�n�[:�5�r�S�q�մK�x��nwwsi6i<{�X�N����x&�: t�0 �f5 @��A�I^kPPE�UBpb�#]%?|���ƽ��>�Lք��O ē�j��,ǈ�~����~$�����Ur��Q�^Z��eF�M�W�*�};-��Y �
�%{������V�"�-�(
��MŢH�
x����jG���<�!7��;���^��X����+�w��cҘ0�f�Vq=
�u=[{�})7Q��>��Ǟ!Y���'#�Ud�+h	�ƿBP�����p;�v�{��ˑ���7]E#M����$�����L�bb��>�CG�og�%f��j+�XP��|��۰��'d�df��4sզ7�ø0�)� ��˘�M7�qw����Ӷ���j���,*��������U��>uN>�h!�E��W��Y�����ٹ�,f����ک�[�kZTu ˩�^tP�ȸ9i@E���B+U�TO�m;�k���ː��#��=ꍣ���4xs����Al�t��Z7�s&����]�ᴌ}or*q�E��._�4Wlo"��[��9�S匱�	���D9��.� !1Gj�}��E)m��[y�(ѿSW?w�����bi��)�3��_�<�t:#��������N�"�_�ᘖ��`ְ��ԧi�5 �v���8�lUR,�����`0���.l �LZ���Cs�������}|-��IdY\�-��tI_H�1JdEx��4�i�&cj���
�I+Ea
�j��9�,�W��.?�i���qk�F�m�0���妷���=p���|{&r�r9:㕛�����b|A��(�7Om񊃽��\�L���?M��T�o�s*=�dn*AW��D]+�G���^��W�iL�\��I U@hM�gĬ���f;�o�g �W�5�k�
.k�D<�=�"�1"���wt��tx���]�S\��.��-����z} ����Z$\���/��W�|H�q���a�o����5�':�^�ZN��O��oR,{br,XN�Mi�K%"�r�
	dD�g&]:>e�C@�PD\@Kl�&VHM@���vH�p"D>������(�w�0y���Wޑ@^" W�O)��c�ϻ)�kOF��>�Y�|X�eO�bS�#�̬e̦�jU��z0�nV�3.�7���4hZ�0H�ӄo%p�P��x�0~���B�5C� ��Z�Tm�?1��]���Y�;�̨��U����s��Vp���񨘤Z�e���녌lCZ�G��C��*2h7LE�I���j+�j���Y���H��F<j��u!��=/���u��ݔ���yo^WȦ��?��2��i���:f�`&���tnTc%���o��D�䚵
��Ҍ
Ei���M�,�X�$M&b�#�����[P��8Y�5��ger��m3�;hw�9�����Q�v[Қ�+�:�3Wޒ�L1��ٟ��1J��:_�lN��x�����z+��L���.��S���M��4J�f9P��>����?�8��a/u�ъ- 5I�W��d��ZQ���_K��ݍA��nn��	��Ξ<��t�6|ٲQ�G���ya��pݣ������g�YR-
�Zh�|k[k�/����宾�/�<~C��z��A����V!b�VJ��*[X�E|?�;�a�v��p�(9a�OP�K%V&�6��1�T-����]eqA��?\3��N5�%![Ft��fS�5N�a.�������U���c^������[����w'�	gi�S�V��U���F�T����1]����17ǧ��1�������'���yO3ߐ��T��ˤ�M�
���a���`3����H�K��' #D���൰z`7��Й�(��5�m����&u���&��3�wD�e%����*	=�q�U.�S�_��xN#���0ڑ<#U�M4ӆ���,v( ����9�΍�o1�E�IlVz���.�.�P��2��V��4���bx�B���T���3.��ZfT��hS��84�Mؓ��Ly�,т!�H��^�l�����]D���-M����_�7���a�z�L%����'�KD`�<SfK�d��5\���.t���XZ�}� wl8�#"��� !�W>c|_��{pօ��@e%}�	��ё��$E[�V�&�kcyŋQf�F7��n�yD�q���vh�c�"V��pYϛ�DaZ�W(-SGa��\+�7E�8%��M��_������oRZ�(T]���Y�4���)�q�'I�.�J��~K9�!��n��-��N��.1�K��7����t��g������Y�N%��R,PP=�!�Po�s�R��2sHVj� �B���5�ڬb���O�B/�%*:=�3���ҝ�6�G\�d�������p��_�}7�2�S�vts��m��n7�M1�����lɃ܂����]�Q�xɣY	,�nH�
��%�X�s��Ţ�dՑ����p7l\qBI@3_�{�h ��V��l� S7\I�2̦��:�]꡷�#�o�'�h����l�)7r�PÞ�N�7�P���D��e2{���ܘ�~��0��д� �_�F�O�_�
k
𶇲cJZ.�3���ڎ!��i;������*�v�|.��f�q+<��\�޵n���X[6f����v�CZ��ڣD�	�7}�i�&X�5�P���OP����&u*���wG����ڱ������Q&�p�����-4R�O����H!��2v����'�l;��'gX�}�:���F�d/���ra�L���"N&㝩\�B+����]��[�������m�f��mډ�L���z�QPZ�'�ҙ>��w�N��`#�H��ʖ���pD�ɿ�+�a+Yf�Ve�A��Id�_�V;v�U�aR�|�t!��}^�b�T���!�j��c��w�X�J��Q�	Ju��G�b����-w6�kz�:ϱ� #��_.�A�Љ =|>��GPC�����D�g~��[�S2)���j�Y̑�\U�hAW�_h��I��2�بm���R�G|go��,L0F�:��ƭ])�l��P}΃d! �T�?��7���Ek�}��=������\֓Q���Վ"��p��w������w�4�o�&ar�����:W��Fd�p�˺J�+��sm8�Bg>xE6��N]���7���L��\M`����c\n������꾇5Y_i�70�T���+.��ܪ�
�s��ë�Le�I��:��5'f��hp���Q�X�ATs�$�X���5N~#�9f��/�i�
�qr��|����Gd�ܸ�ٿ��)�Rl����%�2����ޚ�|:�7�����)���=,�u��AA^�zp�]+ĎLk=��DX�䲭�Ox���ȟ%�QX)%�'���Ўi��aY��e1�3t�>7?��4׉�G�D�EE������YY�ڀ�VH���s��"�L����~�nH���ƩV��-�T�e��lLy�b.D?fTFo�=Y	��J࿰�nfش�٣WI
ё[(ܴ�/*���,(x�Z���C������\B-15`0Ct>t�"A=V[��nki�:�Y~��Y��_)�Mf��Y
+%�_��B/��eb������006"Em�*��L��fr��A����pSe�Bw�gh�A�E13�{��0�Ճ�VI��ʧ3��$�˙����NT;4�&�̰5x���A���d�M�:�@ɫ��O�KI{�oo������7�w���XG��)Je�5_RX�~����Z�����d�)xwyi���S����ϥ �� ��;wov �	��j������c��T�:�)ڍF22,�A�@��gy�$�2+��H��0K�-�3}i��`�';�j&��)!�#y!�u��bۗ̲=u�+�r�O.Ĭ���j���/)���_C˷U<�ò�Y�ܡن�:Pj�� ����I`˃!8"G��xm��TE����2�[�X�q�>�c�c��'�Fpp��'Lw{��>��=�����p�ى/$��+ճ���ׂN%w��Ø�
����?Ѹ�K�-��6���g��lh��b�>G\��n
�J�sK����|� ����h���В7Ө�f����]{�tfbP7\�|��	�#����B ��y�G�̘җ2��U��U@��"N�gyQ A���(��b:���n�HI�%i'����j�b+�#߰Ә�*�2���,����t���!H�p ���]��@)�\�.��Q�v���h���-�L��3�95��=�Du�3�=g��⿩`jf�&�����E��2B4���`uf$l����	�ϛ'�Mƛ�|��LKy�K7��z�[��;�I��r��h������2{7�<����<�X�wu`x>F�?O��ĸs^�n	M��A�5r����K�)���ֻl���r(�vU�s�A$�w�����@�&R���2� @/'��5�����D1Y��ѧ*�|�l(֞�с�v�mvm�5�Ӓ+���u^��}����eh��D[y���K�&��W��rjC�7�Z��&]����z�]��Z}&jK�a"*�jfgq���G`��3�3�w�����,�$v�_TC0�H��iK��D0�����r�q��
ٿ,Z�Fƺ8��r�?:�<&�sǬ[!��g�����>�4I۵��}�Sk��p����$ijN"K�T���̵��	����$h1�r�#�q��3Õi@�������z�Dv�i���𓞇�2��W�R�1{H9��O�Hg<as!Ct���Dߗ��dG�o���d�X>��������Eq�Y��%	�<�,>��E˷m����$!y���Q�
�`����p��v�ŎD�a�س�㞦Sڜ
cn6��b�#,�X��6$t�����6�͈gUV_����.PS��R��]|�dfl��&�maB��� %�&�U��؉�倣>��{�@�#�u<9(r� �~�6�y��m��بU�(-�2#�m��"+��l�W���sk %<�U(�ω9�?*ଐ=��s��� ���Iw{7#A ��*��AJ��7�_��Jx�+d9������Z.��nXV����ǄM����x/����ɮ~�Ý��"���nV^����-ُcp��ʀB����>���x�7���sR$f�x�s8
ˬ�%{q�DR�z"�+3��>��S���Rw�qm������?F<�|� >�R.�B��ֲ!�1~2):�WժK�!��-f�u�#WM5G���⊑���t���';O3�l��wpk�³�x���թ�sRK5L��*�PK��h���i�\�S� ��gDB��q�﫻���ƯOtS����?@�|?~�f��;��잕��2�_�F��A��<�]н�.���t:L�>8sf*)����&Ib�`�^HΔ�˹,J5���$�0�����Z����`o��k�^�"���n$����rb���6ʙ|�^��/WN�J�p�)�U{R�ʉS?�����-��Ak-�֎&�2�h)ҳ6�C��+:�E�����q>p�
��O3[���t!�2�-l�ܧ_��ҐT��j��|��V�(B^6Jٞ Ci�#n9}�sd�bՐ��b?�с���\n���H�c3�t���(X�3q��\ gc���֎�@ka#�����L���,��e�+���NЛ��I�QR��'7ڲ%�����-D@��G�9�?^=�6������$\�*��T�-�����܋
�GQߛ6����G��|R	���ù�>��n}� �A��<�_�u����� &b�~]*(�����~w�yV
��!2<Hi���c6 ��7�����⬄�ב����2\���#*
'���G�;F�=�fvx�E����̲Ŭ߄��uc���я60��p�L��x�ā��Ҩ�H��C�w]���N��5	5}&b���3�ˬ$��o��1G>�o�L8����x��f`(T��4GbM'=��e���q����Ĉ�vd��3���.����<�3	�����_l+��W�B�Re�_�9�y���� i�0d2��`�aw��&���r�c�ԫݳ,���Y��	P�OWic�;\w)�9�`/KH�6�['�%�^�㚰��,9�c�$=�ȱ��G���Z�~n��Ngk,9Iz���f���ځ���MlZڏ�� r��0��>��ΐ�,�\a��tf;R*���/	D�!�ߣ�(V&�����YP�8�C��"=[F[U9M~X2Jf'����W��3}O=Ǖ�XE��Ρ�+K��_,{!���V���:����=����U��H��ll͌Ltj+�r�2]D
m��B��bTE'kb �p8'���寱�Dgɺ��9����)��m��nFg��jQ��
t�T�/�v���w��f�tN��`.�������h��R�c�에��Jj��l�~!���j3;�����r!��6)J�����_c9?�2�Q�s-Pع���&)~��Y���V�3�D�P��@ih|�P �u��ɨ>D��-[�*"-�~!�����3�������i�>r@����m���ld�]����}�*���$��m8��Fk�`L����쫎Jx���4��N3�]�����%E�	'P�K��[�UWV�D�4�U�q.+�J[����}'���l�}B;�}||n;h}�N(���R��
a�,���}fhl:�$���G+�:����^�I��?*ݞ��c���v��lp�U�08ջ���ܭ�&"�|"D��{@rt�q<[u�>�=��i6�y1���,נ���4�܎�T ��C"{x:���?����;Wf��ވ�J;nP}�&+MW�4�L�P�����5g����*�E�Ar���BڗK�I�XQk��id�r�[?Ӫ�����Y��������l��(��s���2R��şK��"�\�w���V �,��AP��!C�T0j]��<���[����?�	��g�
5�Se�ӑ�/��O׸�P��7ˎ�O�Br��p�ʑ���(��b�����L���NvJ>�>��q{|iaG��r�'J�Izx�?HR��Bb
[7`g@�~�&3��)ۺ�������`8�_ԯ�}`�!�2g���?�z}�� �~Z�����v ��:} t�ב"��WA�i�6B�r���r��J�~�пsI�?���gmV�8q��i1W�(6)���3'y�Ǒ�C�[U!3��|qC�m8�T���=�pX!�_ע�[M�H��Op��#ѵ�O4��Sq�q)�pd�C���&g��I��˷gaz�M��r@�%�
��sna������#h{	��M���=�ul.-���50Rs^=�����RE5�DQ�R��� #J�${^��;A����k��)�~)2�q��+���j]��p��©��B�V����I 6�!��7��= �"RŸǩ]8�}�T�2HCn�Y�Cě�lCG�vV�a��Lk�1v)��1��y2ޝ�1Kr������wȑq�?�&�f'���/l�� ҡ<��P���m^1uX�3U9��WI�n���N"/�,����7�hz�WU�^��"��WY���X�����w�`K^�B?߼�xƏR]>�΄���f��
��`GױaS��ogfc=9x?�`�����T��� �X��5y���Ƀd���C6���%tU����Y����<(�@���B(��?k w��Џ���hV�B�k�{FNY��ؘ2s�����"U�� �͠=KΉ���+�C����Q#���B۶d3���%a�)�x�
o"=��U�J�ޮ�mZ���o#=Sj`偱?�\�]'w)��*�����G �q�d���g.{Y{9_/ME��¤�Vu'�G�OP�3JGz%��S�A���OqW��N���>�1�Ҟ��/!��8�t#5��!�_:m�	�ܖ��������f*��wP��ǲNZ׾V ��x�15�"
��Z�(??�C
�w���+S,SY��]��� ��ül�nNou����[�E3tDCت� iU��F��ѣ���n�Ĕ�ʩ�+H��a<����D,?X�g����&��3�� P�Α���[r�me8���;9�v\ۖ��RȺ�jY#0
���
�Hϊ۸��8��u�vv�G
0�I�ֲr�g��4s<6������H���i%K��~Fx6����������,#��ASՄ���"���f8�Dh�1
���&��\��B0�T�}0���
�M�����^et���+[��ͧ���*ϫyY1�F�֟���bT �P�Ȍ����D��a2��n�[�O����1�z"�Is%�萙��NZ�]��س<���������i�������a���h��p�^�EtzGWܱd�a��΋QT>��,y>���p�-ڜ�і�3���S�>��}ݮw!R�@?���7�{����l+��ʦ��2���ޫ��In{:��y ��z�c-� O��ViP���1�.��*'6>I��h��~I�j� ��B
-v=�w��ŷNX����c/�m� ��):ON�>����^�������.������c���e����&������� �5��?Cog����c���%|j�
���3*�S�`�Z�D��]�X3���0N�95}��*�,^<��̐�d�T�mO(����f����7��M�� �O�!ۗ�Vf%�<JW�EP�����r��=���"e�)�l��]�F6�����I&��k��ܴ@�8ג�{�WQ����\�b�$`���j�i�G�ށ dǛ5�%=l����fj"�ls��P�J&��ԙ9& ���*F"���d�[�}�Q�)Jg��=!R#}.q�FP�I0��n2���0�=�U��4��S��|n\*5}��I�*7��{�:̻Ć��ŠN�S9�[��~T� B���lT3R�쪖�g���+�`��
�y�:Ïh9M���:L6|l�M	a[�V�5������+�k�嘭(�߂�����SvJ�G����#5-0��ף��G�<MI
��R�l$��ν^B�ڈ5&ʰA��e�l\G6�O���+�x4v��e%x�Z	Q	�0xj��)|%Sɷ+廈�P0��n��⬡��le��8��
����V`4� 9F�%Z��Ø�W��d�Z?�8�M\�4�Sy�D�����Կg�d��6��U�Z�^���uX�VS�<2"�/^C$c�Q��v����!Ȃ��,9��7[t�I��w:����Z��=�*�:x�����Y`�j34��o���uZ�&E��;�-�P\n�9gZ�jp�X6�J�XM4vi֟%`xݘD���2q�����F?QƃO�fvj�s�x���I�����:��lA���f��jlF����q���y�	��O�gh��sPR���D�j��ސ��M�@��A�l����;�c~�^��jQ�����]\][[Pɝ�j�zdC�W� ����	�����ϐ��o\�#�x@�A�=�`'�j�����-2|y�?����h���
q�B~!��z�&�Y�"����$�t����9�`��#�Z/�dV�	2��M�aF�vQ .J��Ord��xt@�F�Y��)�m�2���>ܜ�y���/v��L�{�S�Y�x]`��3��J]1�=l\TH�|2���T<����z��ۥ(O��|$loi:?���C˾a��!�Yi�[���$f�o}�ԕ��<�_QR��
X���s���K��yt�] f)�����/�;���A�L�����s�H��q����8>&W�D�t���Oa��?�x��x�=�W����'J]u�<�>�l'O�\!��@#�)�+LmѦ�p6�J�n�ӹ���%Y�
��!�X�.:�[�K�ü{F١��v��E�l��O;ǯ�	͎����I�)�8�ZԀ�),�y<3�<��(~haɨWq� ���h�D�g����("3���9)�D9�#�q6E](X8L#��X�w5;�W�[lk@y���-t�2��\�n/��� Re�/8N��k.yB��s�C�P.��$f6�<j���革|��3��Tﭓ��kѿ=�8��5x���u�ɠtvP%�`S�; `��bo�Ռ\��R,��w U��(�ڻ��,J4h��WB�8rjl��15Y�r\��j���.�s���rkd�/��`�Z�G��r�4%|R�7�w�K��!G�#<�1)�M���.t�O�X��q^��#�$/Y�9�CNi�s|��8#
�8&{4�	�e	R0��|^d&�Z?��t�=:�.+�ī�da�vW!Q��.�?60����	��p���L��Ʌ5w�sY MŲ�sIT�d���/|�y��"Z�tTa)k0_��c�/Of$��f��B3��!&q��4����g�qMF�����5C��z[�N�/���L���Z�g�VP@ܐUx�#[}W�~�/�{$��%yy�X ��z+��/���wd6���.��A�\���zzt��N���ʔ$Q��P�&\C	�{˴���)杰}�|�;�dWoF��j��a�]ȡ��Վ0E�s���X8���_6F26���C�!����� ����0��?�K+W'�d]��:��7��̭ĸ}׶I�&�7pe�VS�Lo�0�\fݎ{[ g��s�3�fۇ�P���J�;��F�^qӘ���5�Ծ���h�9#N�����.4b��������=�54�� �đ	��E��8�ۖMߎU��D�ͅ$�w�G+AW���{]��#i��Zq��@�yg5�a/��~u½)}�a���)	�q��^��6'��[��x(��0*K�w	���n��_�.h�m)�q�R6b&6�^�Rf�R%����Ex��o#�`�%2.`�콎�~ى�_�p��S5�����M@a��Hઑ��']���F�I7TWÂx��� �O��c��E�;I�Lh��^Z��T921+Պؓ�8��(Q�+iZ�r�6p�� ��1:�	f�5p���},�	�X�!T�XЀ��m"�D�lj}�AXg'���1��~#%��zf�82����$�㵍�-\��Z�5ʲ!7w����n��)��i|�,An����n^Qw���C���*#����ӱw��~�f���ڛʰ��@I o����F5��yn1b߫�'��{^�Vϫ����#g�l$p%�����*{E��u��*}��b6D@�\}^k ~��.��eS��I!(-q�ٞ�T��-�M���g��]T
b�V�WfX��H���-�0FȈ���L|E|�)|pב�{n��.�\�MJ�;�x�&6�dv:�� �Xq����#�B��o�l�]E::k�{3s�$������`x��-z��i�1�im�>�N������3��KJ��Cʼ����w���(9�n!�mU�+&��d�.ω�5|�m�ذ�E�w�����5K�_�@!��o"�������\�x��cMz-ן������nh���:#eU��i*��tc�o1_r�כjb1L:�Z�L�E�t=�b��9	U�7vŒh����Y����7�H��b9㯴�e;~���_+�3���������!�����ډ.��a�2� ��EG�6q�c���J�}�h�5�|J�t3�͑J.
���0ImF�Al�QS��~r�2O[��B^�Ox�<6l��S�7i�Bk�
�%�W]��-��3��R����R�k�����zhG�
?1�L�ջxE-�j����p~�hT����ԓ�]��,�y8�^������X��2����Gt٢U!Y�uz �c�h��%^kr*�x�'rқ���@y��U �tbC�40�l���Il��D�RM�,I$(��;�V�).u�$1F.5yF��d|!�T�w+!Ɋ���eD�8J|OY��0j�����T������k��帏�m�����eǞ8!pY�Rq�I����)KOt3s�v�U��� n?�vy��\ ]hN�f��9�v���g�3�|0��[����ɋ��Z�jgZ���N���V��vh8Ww@�3q{�p@E�Jͥ]��ec'�������VX$Q"����!�U�쟢[ؙ ��X��]lZTYI�9f�--{��k��#ϔk�0
�hH��Qv�����P	�=�v	����yk*Q���X��qW��)Vo�u��*�<]�(����g�3�,�>��<�5����P�#�m�t��z(	�#�)���qoֻ��I�厕vS�u%��3��\��6 ��@�U(���=�;o���O2t��im�`�M_8*�A8���+=N$������+y�ֲ���7[��,-��; ��a���jDx}�Bs�9Ec�熩썜�4�'��5x$\�䊇/ǐ_�
�rd052�y��ѣ��Y5�ԗ�!����p�$e.e���N@�v��%"G�a�D�9>ɐ���6�bv�������Y�q��{�<����](�P^-�A��\�F]�Zk�8T�(���6V�c�"�ŔR�$�H��{(M|���`,�ܘ�\0!�y4@�^��L�``����I��,����
_���2Y����R�rN"�X|%�<+[ o��K@괫ҳIXP����#�#�$cƝ�;���c'�'��vd����	�׻h{�U��!p�Bψ���]��'�s�s����ZO�����0עv:��	������_ %�N[�v�ӘV���Sd-� -��'F���X��7�Y�&QËݟ��f���Xx�.Щs�g��Zd_��>�!��A�YD
�'9j� �d6�
��a�Xm��̏���9�b~��&�i-�+Y_�=7A:�{���f����Y�F��2ϭܽ#�A����lFH !~d��[�Σ,I�z�<��HK�Ad����qN���"6C�~'[P!0zZ��4��_�v�sϖh1/��;7)�S�;A�ޮSB8�pR�:�oX6�ְ+j���D��/�-��������&����;x���2ѕ�"r0A��7�_�O݉vi��>��ͻzb�Ўt�g���(��V��jP�I���s���l�����V��BM���*$�ϴ<�X8X��	xgb|-[��"�|O$��t��B�`�T�G=8P�N��5�~�&ᐘ}Y,�QO���y5P2 $Qpg���f�䖪��p&��h��겹��1�����2dC��y�����Aʴ�xqέ�||=��}��R���cE	��;�ZKC���"���O|��]�6܊��x�0��S7�Y�	��~ٍ�)5�
(2.l��*���!��θ�����zd*��9I1G2F?�d����o��|X���8�i|o�\U�&w�,�V+7���D<�����M��;�v�@�պ��ťsީ>��I��KM|m��{4Q�Ł���B����r�*.Gi'҈}4��1�yB����nQv�~d�h����o9�s�zl�F�
�l��&>��M���BA���I4濹�	�4Ȏ�G��PCP-�Q8��e �n��pH���(b�]���g���U�zL
�OM�˖5�Zc�cۺTpW�j�BhE���2��pw`�Xl��x�k$_�f\�p�Wz�Gm����öC����Ъ��+￰�'永�h9�*�+V�j&ڬ<B��fPP�z4���"rm�����t���A��QS[	�|�g��6W���j�OG���~���u�Nt�A�����⮶,�m�X��������p��Nza��O*�.}1@[�R������L�Ϥ��o_*���G	\`>��č٧�^�VKN�t$��y�����}<��J�������mTT��Z��C������
dѦ�\��R�
2y;;V�4��p.��~v)�Ml/y��dIq��#���	Ԙ�Tx�$ZH��-�/"�}�܈;U9ݗF���M&�1j��n�Zu7n�Κw��k�|��K��;6�mO�P5qn� .w�B��6��q� !MA��뭧����R��Wԅ�i[�v��!����sf�T��ݗt�),$H�j��[�O8��Ę�c5R;Ȏ�R&�鞅�bDS��o�Y*�s�%��u�����)�'V�oA ��EU� q��qN כ����1��v6�����1ر����,X��n�עK���w��F�����{G�^>�4C(
*����7�-��{Hg�)��,���K*��q�����p�@�Q��v�Fde���`<���<����!�]�x���zfD��Oi#_�;�y�(h �c��ձ���O��$�b�Ë�s���A�Bm'��͡�xp#Z�6{.l��M�Q��t?��z�v�ob�N��͍y��;	ӄ�fQ�YͰ�c!����t4w47#�����U@R���6gkB ��Fbq2���a�3�H�q��V4��p��Z=�2S=���A�L���o$�Y o8�2�,Wc��'�Hu(�?�1���P��
 �-�v2A��7�B�~����#�9
ri�a���>�L
%
C���� �m�'��{(�K�|rJ���X�lu�"R�+G׶�=��c�4�h4I4��cvo�h��y��о��ndn��!�_�j$��s��OP��j���٠��/7�F��������[E�=I|T	x�1)V^��Ju�}?'#���F���c%,���Kgun[(s<	e��sF2��))�M�8ꐊ ��	��Xn���;c7ω4ؚZ��pB��c�1+��4�]��y���j=6|��F�Y��B�TY��\$�0�r
խn&PtΫ���[N����&mUm�	,<������� �
�f�4�	��u�:�ȠV�ꟛ�%o�;�!���=�`�*�T��._����4�,�,�M�C�1�{7^[A���I_��7�t+���ޏD ����}�IpE�sf�(kjU�^8�� �e ��#(u�v?a
�T8ڨrX~�p���2䚚ٷi���4硐�S&~[�n"�u��-$P��Ly�G`wjse�f���A�tjC��H������0�~�z�BN�e���������7��~k�!A�0�{{���LHA���q�)i�>_�R���Y)�;lZ-�k����7��;a]��)"�� T���c�8a�kFL�NT�œ�7IȼA����I�}<�ð���@�:w8�U���d���KQ2ݍ)r���Lq�������b����O�țR��R�&��a�mgt��5�>�<�`�E/�B�͔��1�-�8ɽ��+,�ْ��o�b�����e= �U�2`ޝ^����gVMqngUJ��c')�6xt*�:aG���8�v{�Ϩ]K��$`���>�V��_�����]@'ZN��A2��\w�#8`s�c' y?����(�'���Gt�
k���R�@'~����?G�B�t�����|��I���4Fg�C\a�'��8�|�\f�pvD��_�r��+�i�N��u��\yY�%S��jT�� ���z����zqߓ�2�����+l_t�SpO��]8�E���'<t~��U�f��q�2���PN���(�.�q	�C�T�ܲ��\3�32����E
W��f��3���bi��u%0i���~�Z��Bܲ�$�|�e���;i�J�
�lA�^D�����e��f�0�!�`,�K��ɋ㤫Nq�27��7���B1'?/�!;�sV�ُ�$���3�=G��|kxc�ZW��'�����С%�Z�r�OOv�q,�&�ڙ�wu&�4P�V9���j��ޏt���ޕ������K٘^8 ί��S��M�Ztc���N����{��+��;��C�(����[��!�ڿ�ā�i���I����8��:�h���u@���H��r��[�
��%鼣TBxA�vS+PV�&�Z�ٰ���NR�Kד8���T7���o5�q�_���Y���[0·�g�O�Ԏ�wح?V':9K���6�Xfb�>�[��4',3�_�������0<f��C�lQٍ�¬�A�������j���BO"4��L�����A�h��\x�1�m�b��L9�x[���Kc����3+��I ����ͬݢ�v$T��<����eW@7�d���2|$֠����׻@/J|���Y�M�$�=|�|���4;�ǝ�\�������Z��5/���I$R�1�EC�8?L�SeQu���1�`��Oh����!1��fN�Mp�4;L�������<rœ5'%�����A��l�k7�Xq�9&��-��+e|S6��=��.4|�)�k�Ȗ�Gy�pl�����|%�H��ґ6��2ؚѵ����XQ[t'`�"�\&7�O0����i�B�ڈ��� �3+i���`�P�Ώe#�z�iR�(��@ 8�G���1�٪k��%�7�̆������[� �80))�*y���t'k��M����}����F���N�"��Fأ���*�~�CfʭAU��3-�|]
�U}/3r}ܹ��Ǎ'�hL���� {N�ʇ�{Q`)�\j\?6�=�*��W�2�����!��CSSаܰ�|�:�C���sI�������!�/��%�H��~�v�&��B��+��9Z�F[O7#���mk|p���D}?bIBq^��������Mݔ���ٽ�����fO� ��O�?X4����߉���Q>��M��L}�M-�����ُU�pp<E�ޠCH
=PX�q�B�lQE.�W1/1}\��jq �L�ÿm�^
�|��Q��ߍ�5���v�%���s�sU<X7�(��>�L�r�8#��ƨRq��e�y�������)M����:�-�)�|D����Kc,�JeZ[σ�H@D�˵�c����3�}&PWu�C䋅8�{�9oT�����󶕿��m
-с^�옥�ʧ7c�<<B�qgd�>��L"��_\~�-]���V��(�KO��G_��I�o{�#{�.����)����{{����V�M8�߼�麦nT9~1����g�����Z��<��^c����#��\�~� �s�(¡7�����$M>q74K!�#������{��{D��Z)��__��܆P�ܢ��r-Z<ͮ&�Ǳ�?^�i���ތ��)��쟥f�o^������D|Q�VJ�����g|Sz��hxc1Y��=�]�M�����sx�&d{.p�.``��d@�̴:�%�8���i�#є�{QZ�����!/��~��bx��E,@�&�w�b~v����U��]VO��N�ض�
�X�o�K�`~D�����R#�=�}�@46��@۽՝
����JхQ:	X"`�"��뤋� �"��neD�}���)��"����G8���k!G[��̉�}2�����+K1
f�Kke�^�&A~��A�q4T�a�{3J��S���������3�;Sۣ~a���q�Z������� ��-���v+����9�o6�t�;l��ή�"����($�k�S�m�4�FU�~-2SVS�5�t�pS���F5F0l݂�9QND�#�	p�����RL~�Y�r����`�GK��I<x"/q��E��+|�<�'�i�
��L!r�TB)1���eoZ����l�WW��� QR��SX�'i"���Z����o�����eU#�FJFsv���q�.��g����Qp_�A���]O�b�����^�z�vؑ���LHd�������E����yY@a��_]Y�Y�3Z�Y�A�ǝ�hLir���$�P��JJ'�U�~�F��:n�Jh�笕 o������r�F6*�U<ygU�^������Y���� �=��ʌa)�Gg���L�L�l��7���ި���YO��8�4���%:�&dB�vj�q�g��l�>����N-~E��z)dd��'C#��Jv-�$�8D����vW�S��x)��vi����
#m�)�ɦisP �����5G�4T�
놎�(�S0G�藾.+������:\�v�"�K�q��ύ��r-E�ԁ��l�Β,p���g��Y��ݻ��EA*�����ץH�R���iL�= ���O���9�ݞ �$�2j��Y���f#�V����β�FQ+�
�G�b+��WtS�N�f��!'f����Grr�jo#MYv�*�.��?V2䥍�+�@�iZWh��!E��R���]����� !�N.�\�k[ez����w����y��G���	9�@!"`��p�6��<����./%P�Rv%�]q����:5o���V��M�Ŝ�M�N3�ŀ����!\v�)Iף��P�Ӗ�E��c33Cz�`C�ו�Q!�oC�/�k�oRl�b":�g��@�l�Ő}�7;���QN9����5��ፉ�u��W�g��T��=�C��ʕ����޽��pN��F���YƊ:O:>R�)��mp�v��!;=�-������PQw�d���*�������^�����@6��⌛�Xr?n<�e^`���ʑ6{���}�kr��O`��q�� @��d9j[U{�L/�k�]��B`�6���ϗsɸތ�ž��4��v�E:t��j�Ð2lH-�7��� L�X܏�x�-߹�z��<g����l��;k`�^A��{��1i�#�H�$�[|�a��V�M��lr<Mm0�2��w¿��x��|a��y�7����N�T	�'^�Eⷼ]֑��&�|�vx|�e"�[���2�?D$o���[��X��XY�5�~{puц����s���)�X6wEm�َ��=t�B��C�x��6d:l_$1�� m�Gk�{���Q�hDNRF�ߺ"��nE8��$�󌁛���Y�}��MO�s�Qk�7A�k����v�t��Q��2��^[K�yj\��'5�^�6�=3YD�K���א$�����T$�oVVX?��/j��|9(�L}!n�PW��)�U~7�Q6�J,�!w�+�����Fx4��k�8�<���*�lz�ʗ���(:�/u���%��������5�� ��ȷ��K��`F����M��{:�����4�GH�H+꩓A��7ވ�c��b:�da��Dr�ϝG��t��a�~����lX�.sk�u)�P$��^�R��Z�l�Rz��h�,�Xʵ�l3���\�55�e�gλa�����G�#Dv��ܕ̵�"u����_߿ϺК'=�2߹�ӵ8N�":��	��y��Y�h�˞M}�L&��>0^��J�.սۃ%��R����!�&IQКN5�>�z��e�� '���������d.��}9��$�֋&H�f�t���]�� �PД�X�|�Z�@��Y�F����/\�����2!�|{�(]t��Őp!�K%���<w	2�x[��9[ Ϫl!�;c����( ͑�Y�2D�U&6�$��jq�����ʐd�
LZ���u�?���?�vkM�:2�k�մ���Pxρ�޽�q�$�iWA���OQ�As^�*g�f.afގ����dA<��Y��~T���'잩�oz+��G���.�`�="5��%vc��ļb$��<�\���N���Y�b���!�@�AQIَcG.�R��˂���AH+N�e�Y�ZE3��y�,w���t�O���:ǈS[ӷ������O8���M������R�2`�����<���O�|ܽD�u�\��=��inQ[�v�S�|������I�<7E���fw�rD2�88'L貆�I���D���oF��\B�Z$���Uf�C�
�H���R/W��������a�����6���o��[��A�t�o�=�s��bA⪼��<ԕCr��$��kQS���_N�pg�㐟{�V{�hr7Ԍ�S�U�K@��E���k�Pd�u��.��?V�F���E�n�~�����.`�c�+Ld��	H���J8J�h�?n��<���g���dz�N�;���Ǎ����w��E���sw���V�����G�Z�F��On�+��5^�ʭ nH���`%��vu]n�fĺ�%袞��c/����B<Q5K�C��,��#}�b��z����M9CF\9f�%Gy�u=���0e����ob��;�A�sf�z�V0eN�I�lrɕ��mL�$#�� Ȝ �I�_�r�B�(AM��8��,	{���-I���Q-��$
j�,&��7a��e��t4V��6��Q/<�J
�Z�53�{�à�)-H�Y�$f�넜�*0V�ݩ_QV�_��]��ן�ߦ�e�������V�F�|�14�!"���?��)y~#����_�/�J���>�С�t����uӤ}=x�����̼,x�Eq��2�\`�]��E��ؾ׾a���Q2��~�A��	���ү2]��Jю����/��fΑ ;��0�2�m +z�ıH��-m��;:���[��Ȇ.y˟����܏A^)>h��ÉG鏗ə�����2z�91�рVM���B*n8y]�M�	fV��.�HE1�G�Fښq�˄�6,4��z��g_�I�E�{s|��S���х�����|e�q��'��=\����r�Qu5�q(�/?}&�*q�=M���c(�:�Z��*� !�o��35P�VR����s��\ңd��d�v���Z�/q����|khe�L�ƫ��0�i�f�h9=���sUf-�a�}�u*QbJ�9˱*r�^�����*ލ� �@�A� ��g������ ~Q����Ɣ{ru3�����5�^�P.�^z�Clk��р�8�nb/���i[���^w���m�C-gy�
�VEA+~c>��J�xs��c�5\�<��Nx	���ٱ��-����!-*8�P�ڧ�Ӌm����}$���C�����q0���wG�������^�d�e�`~�0<J���~Ie̘��;g����x���d�&RX�X�F�h����Їׂ�u]�d�J�?�/=��\B��l�q�ҙ�5�PY�t������mB�G�A��ս�ͺt���g�'�=p��o '������O7�P�-qK�n�}%��c���^à�+m���#���_�Q��"�3�I��f��Ia�%9Z"3A���ٵ����=��+K�%`
�x|�M�{��>�����}�ܣ�`��ub���E-�9�ju�{�[�.K��
N9p�-xTp�l=r9�F��C�P(u}���<!��Yp���g�~`�s��]��\,�R�Ղ��Yq�9E?n����x��3_�u�:K�d������Z�l�&�E��
e��y�k�[���m�1�o�װ����j�4��7���C�Xg�j�A��H�#`���,�,m�qm�lA6P��sdTME.��8���J������Dm���BfJ+K�i�~4G㕫�X���w��+
�S�A�O4ҏ=\��}.�R�]��@ݮ�~R���Ԟ�0֫+I3G�����/��~(A�S��~�A�0���2���]3���p�������sv��jVNo�Lt��OT�@h�G!b��������~���� �f3��b�~j���0t*��	ރ�a��@8��v�I*�m��p%*��P��*��')I*���]��rǺIV��y���(�j,��1{����
�⏠����=���Ncb�mIA5�дP	�/^��h�+g+�{x�NYb3=�D���Ꞻ�BE�~�y~Ɍ�t����|���^n�K��b������e�g�G�(�V��bK̾�+���+6����tI����)ü�)�� 9I0UƵ�}Gr�8��Plnt,H���0Y�s�%,p|4Z�3��l��<T��\Hpz��-8	�$OEa���_J:����X��zo��[6�M�=jq�UM���������g��OgG����uP������c6��Z�'���Xw����t��mՐ��S�af^��0Q�QR�[�)"�1B>\���ȭ�@AP_��s��GI}�����j���k9ǌ]% ��9r��f����e��\�t�~�����S/�.�l�P���M}��.�Z���̙�݃��l	���+��*����v?����a0�����h%�kX?�)	�������*9��TVJ��ROn]�����\�a8yD���MHu��{�&mMŐ[��O��Y�O� M<�e���zi*�-�G'B��8�l����-B������e�zک|�=�=����(jCp���]W2���	S��yp5o��=�� ��<�VC�7=r����,�vJ����4�#���3�����w5;�Q�/8��o�E��'^���������ĉf\ΰ�,�w��;��x����nš�❞���ӢI�>������лCO&��M���y4���K���=_R=���ISx�YHP�ΦV�t��s���-c�ڵ���S��P�+v2�W��%X��|$�huC)T-���|i���sq6�(�ېSp�Y�� �o���ƖX4��wC�(�7����0q�I)D;�����ŭJ��c2�Usѿ*�5ݢ�K�\S5�f&�U`ʮg#��cp:E1)/B�S[�v��Ο�E����է��1��ڤ>p���׃̬�c�� C	�P[?���G*��?L�."4�8Λ�Q�o��a������^1�9�ˉy�zDl�k�o�DW�D��I�UgQ���tk䲁�Pª�4��ꭤ� 		�в�ouU��t��<��nl���防���hr��� �9��ߩ�чbyQ���D�;M�1�h_~��F��m��M���i��07ĮA��"��v[�lSJ�J	�m��d=�*:J���G�8Y�W���0��(M����ù��8<�W�@�yEׅ��,��ϻ���"}���W%�I<H�#�S�u!m�3�9/7�8cn��\)o�}Lf�{/)� �H��p�Nrq��g����]d:�(&�������]���������B�s��z�+j���ڼ�B�������∩�l��WS�*jj%S���ͣ��/u�~�.Uo�T�������<Ӻ�eh�>7�W�§���$;3���.�?>�{�Ůw�����;z�KO�p�@���K��i�=?AĥzRn�x{��x��h�~�4�$*`Z�����f��-ց��F]#%�O)�O���Eݣ�ļ���
TG[��6hW�$ׁݾܵ(�:��y�7P��3�	z�����λw Ϥ�;��㈂�Ŋ����X� �E�DF8(`u�L	�̳B�>q��.ݟ"�Q{�� [\�]1	)T=�;�\Y"������2��1��6[��tL����U�'Tƨ��\��oGln���X�q�4v�m��^��)j���x�:���,BC�~��WI��������d���m�A�`��\f�I<&J�8��M�E��@�S�}I�*]�6�U{�Izy�je���nn��B��X�!ʖ����E-����	S��"d�0����6N���8��e��Ќ&�����]֋��E�L�y~ɝis�#��>���)����֋�ڍ�Ck��g��4m�s���NJ���U�e��m��<�WI��x�T##�6������-��Z٦��K]`�G"3�W�F����*W��&^�*�ҿ�d�(������r2�E�f	:Q�;E��Q�(I;���=��Y+�D�.p����~Z������u���#�;K�!��J;��z��/w~� �j�W;���ں�U�b��Gf�dE�,K�;�&�P=�I�?]��
H�<���Er��Œ� ��G��������*������%� ���VN��W�S�u�v���p��xK_Ј��ʳ�V���v��"���Ć�[�P�<ː�ȧ���pq�=r��Jn;�_��;�^�|f��w:S���f}St��^�b/S����ãS|ƴ��m�'�Ѷ��z�Bڙɀܻ$��qh��QU:�S�_v #&��.<Ί(��N,!���tL���وn����<6�w.YT=�QҟT�Z�g��L�5�f�R�����l�x�B!%2D��J;�5A��$@P�m©��m��K���t���.o{�y�f�i1��I8��h�`P-����!)���	�<��
�*�B!x*����6�'+�#�%�I��W������KHl���L��_9����l`�7�7芸%��Ӝ4��¿@o������)��q��۩���%��:*�84���.kk=y��h��g-���QC~��]I�N!�"��?N�ǯ]�N<�� ��� 3
�"�uA��a��� �-���P�ڱ��c�֬u����Zy0�.�r4�z[��4�*�Kɗ�O������\A��畋����[&P~�*����T���&���D�6}}*�~�p����Է�炩oy<��2?\9A��$
'�?��ᜱ��6���2F�!�?i`��1E��K@+���D©|W�2�$�lRR�B.�ьw�	�>Ϟ�����iS�vFb"=�����y���$S� W%zu�$.3��=w���Ԃ?���Y�%S~����������r��SQA�a��/�����$0���~Ɯ�Z)w���Ъ[�6[�'Ό<,�D�g2�p�&4�ng��&�t�B�Lr���2V�����~�"Q5SM^���#�@]�E���Եt>�m0]���JA�� &P��n��K�O��Km���;#�5�qXR:m$��2鈉e:���������*��$<�',8!<֠�HN���-��I=I��y�ʋ��	*�@�y�?� ~y�2��i�N]�ٓ\ZD:������O���䒟p��W粑�{+��@�WN���|L띌{����'�w���JǇF�����������]�h�$92b=Q��A��a��!Z�-B�Ȗ�Ŵc�������e��זO��sO��Mɟ;yVlMJD45LA��ksr��!�sSA���n`ف4a�.�6�/�����-���5�*��ڭ�nބ���>�5���X��>.WA9��5�O ��-�"��Y�s�ǡ�����gy��h�8>�[0FJʄi�`�mI�2�pN;Te'jo�%c���c�jD���T6���(�{����{�`�?|�Q{UF� 7~�8�n�����5�Ð-�@�+1
&�f!%�K��$�nÊ.��Wv� �����b��D�'E6�*��wJ�q��?���	�'�~>J
�3͎\4��8w�C?�ɨ�C�G�p�#�\�V.Nړ���	&?Mm� �:O4�}���N%0B*dϲۀ��/�"J.ׁ�.T'�HlD��v�h9�z8��![�x-h) N=-'�"�,�(MJ�0��}�յ>̄�:%Po�/�A
<��؟p#(�����	��Ǹ��B��o�V;I�T�����Xk��뺲�'|�~k
ר��0����zcbH�Fh�"li �r����5}��+^0�5Ƣ�_�&��n,$��M���{�qf���"B��:q�M�<v�<2V�*��25OO�p\��������y͛��p)Z7t�9�P�����Sq��<�m�D��5'�~-�F�"=�u�ѬLsӟ/T|�0�eB�����6"���i���ĩPu��{�3�(���}Op����%9=Q�[�Kk/��{7]��7���r(�J��Tw�����Ƌ��uU�Oo�[]�td�aQ���c���A��x���]���G�c��$�n�X���[T�Ѫ�1�P/_��ٚ���C� �)�J&��Z���{�����&�x<��o@s|�,�E��-��ԡ��HV�C�����OȆz�"�j���<Qӱm$�陱2h�C��y�F�ec�����=|=�������S�f�Q0�]cS��?�����X^�!�ɏB��v\�,�����r�ټ�#h�A�:в�tu��Y�Ǡ,����Tݒ��.K&u�N�ǆlNV'�f��k|��L����W�Z����N�f��Mø&2?�|~���"���-��7L�R[tI��@;k��{��ҿlt��%�dozʣT�C/�@J���E����Ub� F�'r$�e�e*P��lM��4泮@�[� ��9&ȼ�������M����6�Z)g��� ŵG1<+�4ĸ|�ȍ�G�!�@ME��r[-�XN�nC��?[�����W
���)Zf�ЍYP9�ʑ�;����ωC��Rc
.�Ԃz��PU���9��隑����ŕ����y��������M�����˒b&%�dHb�ۊd�Y%e���'AF%fϦ�˟m�Ag��~j��]YB�{S��(U�hl�\��U��������+�#��誦�-x��i�������{���Uӌ���=8�>�S���`��i9\ϼ��K�WM�y��rip H����]�[3����3�M��b�K���n�p,J3�}�:�F"�Y�F���3M�,N!�7N�>�5gƸ8Ts 3i��q�]��# p�x��]��dtN�Od��4�) q��,_g� ��g@�z�TXη���o<��xY��r��t4�a�h�W��S�,艥嶙}�oR��J	�G5��O�?T׆-��C��+���-)}�;��i���q�s�CL����ݲ�:�z����@8��3��&^���sH�4��������<d�f_�ˁ�pۚ%5���Sn�ZPDTm?����������~e_x$u�*���-!.��ףs��� �K�cf S���E+����=���1$£�i� l��n��R��a��GtNǉ�5�we�?=Ne�n;�j�"��j�s�KŠPm��\�$T��[�^���fy�� x��� �z/߉8AG�A���Du�{$�_e�Ƃ�+�Hܲ��G�T��X�_�X�#0�i[�1�{�_�� F���r��V��w�RB́�s7�Svp���A�(��
c36}�++�s�ol��-���4�T���D�~ؖ˰���dJ����9X�w[X%�p����T-L@�礽<�Eo��S�m��K�	�J��3��#$WX;XdT�mb�t)o����,l�H��R��$5i�v�@�`�?�7&\%�}:뾉���b��o:�9q��5��U��~X��L�4g�Q4ܦ$�2m���(�J�+�����?�I^���&�����\�~߲�p�N��v`:��Qƞ��Fc�#v߯dLwqI�P\�F!�ڲa������Ë-ܵ"�$�[�(��(Af�6�3�L��Ԑ�8zd�s5�5���>�V�=^�y����ڑ��5%6mb`����` �$�<v��j��&�
ꄳ��|p�z�CR�:R���(�]3Kr;�ŭ�E�8Z��`UbM�'�L��M�A��5��T����u �����/ڇ0Ȉ���
��Pp����a��x��d ��MM����]�P�Ty�wƙh�NL��=?�.Lk�g�Ax.1 }8��擹Y��~��S��t�ɹ/�:gWCEت��#xS�^�W�g�GC�/������6�.�g����d�'�=�����F$��~���ط<�D^N�a:<lzI�{(g@7��â#ϕAM��g���57Ba(���?�`��|��K��k��%�����x�T���^q�?Ȱ���ZW����Vq��/���׽�`�qW�ӥf�-�T�f#����B��J���7�VA2$h�W�gt)�[���)�9�p\ӄ=���|Sj8��r�����-O.�K������IwJl,� ���֫��fo��?ݟ�L����o~���}��%�q�Ym3M�b��BC6z�n�w��C=��m�|G����/F�3�CR��ڄ��.�������"u|��?�H��(DC��F�&
p��֙��� �/OW���&��,�P.u�����KL�ǯ��Zy+q�kq���E4�+��{��W�sM
�}��� ��WpOEc�9Ű�֞�G�:)E�+�l�j�08�?�YN�Jkޤ�'�d�3n�r��(s�x���̷sv���2���3%5l|�#ʌ��L���?���*���P�����O�*�n	nɕE:�<�mFƛ!����[=���?�M������?�B����|��h"�Y6�	���1���|�rfV��P��	�t���;��GsA��"��1�i&�ec�sB�!�s�)W6�����{Nҕ���Z�݈E�v��]}��	W�?OxZ��u߹�����۾�봈B����i��7lt!��Tu��Ix� S�6�G�5__UO�.��{��횷��D��ȹp�����	@)�b�L��v��-k�Ն�^v�
���
}%	]!ޒ�r��w��Z�IM����1��Wh�S��$��x���/S��^̔���@���4tf`>'dfC|3�3g̢����#s����Ff�CvG�"u"{WԀv���Z��� ���U�~�+�� لW��-���*��(���g��&����TamG�3}=��er?PI�a�**�� ��I���r�P��o�g�0�*����/���=Ђ�sA��9i��\$N׸�>�c����Y�+�I�,����v���i�8Vw{I;�(�lC�$�x�/��b:y��(�]�Nam��C���*)�C�7��1���j�ͷ�ǖ�n'�S]�kz;x�-��[�ϴ�G����/P�ޣ���X��b����o+(@T�H-�U�f��,vD\!��q���=iU^nǚ��
�����"qftf��e�r��~H����>�ƝtL+�󃯄��8~](oصNؕ#T�,�E�Ur���4\��[#���ƴj�M�)0�8���(1'�W��v�,i5u�kv-jr�JiJJ�\���������� ��6!(�rx�j��>�ؖ&�FGF�1�8'�QW�����~�k�T�o����5��i6D�V����o�@�ot�CP��F�}��Wrw�e>�"�����Gt~H���C�6͑$5�-���Æ��	���^&�B���gd�##CW�<r@c	��;��\4VBt��6Vm��]&xW����wv3
}���[,v�'oO�7��wp#~&�2�mM���[X��9�t���:�0S=�洱�gcX�Bſ,6/��{��H��Z2NC
� �� �<-��X=<�=E �`���^j����mg`&=%����P��5kF��p�4�N+��!���c�`�N�G�=�������pˑ�y�FY���ɸ��>�C%X����x�:x1�'
+��x�U`)�@��4l�Ty�5qg
�K��_ǜ�~����y�*=h���jj��OȬH⇹�u-�3�6O�+�I�0��V]Z��mZ?�>2�v^TcKi����mX,j��̬:k�q�޴I>�4$� ��I���o�W�C���bwU�KU�~�B��-WB[$����i��fbk˨��3��.�2/�{���B���M�8{V4�D�]߬�m&\��1+���!Ff�B_9X"@
�h�spൺә�2�~�q�L�l�u���J:k�"_����$7�w�8HCg�tb��vצ�r6s���bG��Q.ھ�bs㴛�;c��B�㮬x#��9���"��>�=]߉Vyy6� 0��|#����ј��ZW*��dՏ�^��N57���EK���M��=v4
�Vw\8=i�:擏��E%m��U�w����ny�|*�шT��(��!a�	P���tnJ_3HX��	6B�ƕǢJ�0C��K@��'����AO�yk�:���G�x秏Y�O�L>X�q�~�qQy��NU�u/�uk�nD���Z�F'�l	�	)����<>�NP	�^:ֻ�Ur��S7�n�˟����yRQ�ك�Qsp`��p9��N�`�mJ�s�L�P��o���E������b+������q_F�5?��Y�pb�-7�q����.�a�I��d�\�fɩ���y>3g�?|S�p#�H��Tg����]��w�Z��S���fl��/�#eZQ3=)U}A�n"��PL��s�
؝�'��;����FL����tBS�O3>�~ ��,�C���6t��h���9Uzf:X���?�x?;�B���tVW��D{��:�t\7������!�nR��h�1�^qv3�d!���'��J?�'X��`�)���܆`�M��`j�P%�����*�Z�rΞ����T�ŭ�
y��Q��x^��K!�����#j�Yʟ�,yُu\�$�}NX�ߦ�,���=�o
��8?�����F:��]�a�UE;�y�̽��/�C�$:5�zQ:ѹF�������ٚ�v7X�K��È(ʉId�7�j�1�759����+�^�R�V�K�N[�V���=�O��9ƚ���Z|QN[k�Q�O�$�G�r!��3�%�3���[oJ���W��� �ط�W����=��sx��$G��}��d��\`1�"}G�t�/+���Ю:�k$�7/�N�΁�bC״�@�t��РA��*l���z	�q.�j�[��cE&e�D�˘������G�1G����`i�̐�uOt����IA�a&R$�6ծ�^fM���{��)9;��q8U'���J;Զ�i�$॰��H1�}��H�hK��9%� ��{3Q�^�]�p̈P�Ϸ�v��U�E�X�'�,J��dx�Gu���+�~N��8�V*�11$.h���)u�:w8g�J<͵��ð�Pc_����h<�
�Am ����5��n��8j����e�1`����ו��;ق��)1�]�G&#s0���D�
EZ��"T���=��$�޴q0��|���:D�I�$�����X�Y/���+{��0<k\�
��rB����0�j� dw�,���j���K��~F���V��+�qk��5����w�.��|�il��*l^�lRY6i$�XY�k@'Y�w �Wx�q��2�6[�d�/��T����v�v jEG&\B���8����YW�ŝ�g���9� ����B�VO!NOt���tҁ��t�,�R��C�]Co�5��.�S�c��V	p��X���ć��iX�H�om&�3�P	U}S2���#��A�*Nqg�1_����2qӱ���oX��nG���Bvݷܐ����z{��S���JNF�
��t6��[��z](0e�+�,+bHں��pl8ȣ���:�C@�A�l�H�*<�����a|��M%���f�p}f�Vr�i	�D���F$�M��]��O�4E�Q{���P��-��M��Ϊ;�;�v����g��g�=�Ujޒ"(L���U��z���v��x_��*�B�@��Ɗ>Gh�"e1,��,�z��f"��E3�� B�C0�g���P�;���)� ot�L��s�N���ݩS_�]z�Cj��p�B�l��[��m5�L�|�1�8��ny�	�%'	��M�[f��g ����S�������Ă[3#�i9i�%���,����v/��ҳVf	�������H3�ҥ���n�E���˔�rL��,�Z~֨T��Lя~��L'v����yZ ��}�4T��ޅK�h�vf�,~�~�x�P��F�FS.?�H��3��J{k�T�u>����1d��V�Ed�X����J
1����/��]ZJ��6J�5�TW�n�G�|2�������?�k&�i�B맢1���ɧ�O�����Q�<��цciy��1��׻]e���gy�:J��7�DүG���Ɋ����I�W�Z\^=� /Dь�
k�Ts�T>@$Ec�7w��'D�Z�s������VØ��w��|�Z ����W�x�&����`��=��u���XGU�f�������w�����G��q�H�񗽷>�� �q*1&Ys�����_��>���W���1���̋"���F��X\�Tm9TN���E{�p���ܠ�<�qz��";gEC�<�c@�5幪���-��g����Y6
J��t�u��f��>�~�3jQ��;�(X�����;ݔ�߀�r]���ի7��-ju�\躬z)��nvs~�Tף�	��?�kJ�I8�E�I��~힟�T�� 60���f[��;�$3���i��c39�BIO�μ*�R�Z�>�ƸL�(Z9B�K���D0�E���r�d�����}�X�N�
� �g�RxJmG�ʶ�N|�o�Х7������������ٿ��� �ߘC�g���w�� g�n@Δ3:'.� ��[gD�=�M�b P"tɔ�OR�R��_}t��������E�R�@���*����hz���閨���%��e�7/3	�ܛ3jp:�Dlja
-������8��H�⎩I2��Ң�R�Aq����}&�DB�-H��s��u9����Z2W�eGur��A���"��SDB͐��9���Ƅ���A\�� �/%���.Ҁ7���W51"C�gj��a�k��G���E���(�}b<x�s<f8����,cź �c`�1���:�_�N��*���8���`G���bX� ��GP�ԏ�M5>��7��Ma�`��T�u��δG�t����c%��l�~n�{BW���ꔕ��7�$�p-�8S�j4�1w���4�o��tZ;/l5>�	����M�s����h�C�S��@JM�p�A�G}��{�Ġ!!L�uM2�Iu�_�)0]��Q1�Q.�7��KX��YNv ���@�^r���a14Jg�L��;!�!���]��t��)V��뮠mp4��T<ܽ�	7��+��u
<��;[�˫,>�����"���(v�k����D<,�u݌W��vG�OU�K��I�ɍ��Ӏ�X�K�n�r3��)t�)+��l��Aw�6�l���.�ض"B����@�uK������p�Q�3N��������4��� �r=���K����1���P"��Mw��gZ?X�?��/?�޻Q�u�ýϹ��䮧kp ��l'�����/�H:���o�'\�c;h��� ;h}G�����H9A��' Խ,n]$��/�����c���FΣ][���%�b4"���)�0sD�~7sz����-V�	��K�s�e��Xʛ����n8rs����w?��l�:� /2N-
2�_�t��X>�0�������)�:2%G&�)�� �`�l�o�෈a���k�ͱ2��j.�B!�S�-�2m��Rf:����-Y��
&(�+$U1?yd�8��%��%����m�|�/�W�J�L�tݡ��	(��w9�6'V�8��B���?L��&.1`ܿ� ���AmnA�c����/]�tAPj��g����#�i΀/�����������fS����ak��u���u}��N�M����~qa�YκCuW)�ʐ���k�=A�� �A���C6��e�Wa�B��N`�\��s�V�'_�9���E��6��T�/w�Ԡ� �Xb,:D߮���Ո?�«��=��[�Z�\6��I�@�15�@���v�1O��::������>�`�dN�m��|���-!w!lطm=m�F�*�Kb�rI[�F��M�{d˴�˾gNɚ!LG}�a*̦��@X�����+��P|���Ǳ՗RGE�Δ�#���7;U�kb$m�v��b�/(��F��l�%'M���1Ƭ�d_<�&J��I��G�����]�$���v�+.�q�^����&ׇ7��D����;/�%��]V�g���,gq�㠿�Zప&� �|�i�໖��2����pwcsA�cY����Hg��YI�.V	�z3�t)�cc@����l8�E$DY�z���W�è��H�>�	� ���V�9$�|���e�5GД)��4��i�r��L7VA���B�[�
�M�U}�"��� >�%,H��X�q+J�"���8��o3a����&���D(���o�#������񢓨��.M�-ȍ���P�4ǿH%���*�?�]��%"� �`�k+�鑠�Ȧz���u����Hfy�ߠt�!݇����	7(�q��T�I	��VU�f� w֕=�N��'�u���������ҥ�{�ʄ�կ�
�6�A�Ώ�*��f��#�((&�kZ11�_au��3�Y�Ȯ�<�	�k���M�'IѾ�4fN����JZkG����W}�}�X����56�r�l��?`�DA�?�=N1�M��	���·+�Z�LM��7Q�"�3�bI)�F�\Z�U%D�șʯ' A��mX����	Wf][��﫨|F���$��rh�#u&�4��l�0=gh��.,��+!�k����_��a���H����H ��q�,��]�~�"v/Z_���[�Y��{�Q�x���]<H�5�|_v�}� ,9�PX�OǓ�f��u�e$�Pd��S�Qr��G
��7����B?[9���o�T�82t4�Я3����܁��ߐ�z�g��@V~��=��c�]����]>5���f��o���C�1J�������,�C�<��GW��ĞM;1��FWk{xk��>�%�3�M��=��J���<��������t��D�p0�i�ٍ|�)��#�z�X_qZj���|��↓9j�`�$��i�/��`*�}$𞳽��WJ�f�C8�QE�*0K�����@@v,RW!t��3@2)!��0b���lo9a]� љH<U>����E�j�����~*|���ͨ3�yb0�a��ct��)��3u�i��-Ɠ9k�qJ��������om�q+,"����q���*��W��ݰ����<�:�������V���
����3*"^��9�A�8�vS'�4�J��8]���{V���"��*�C�H���̴ɋT�ڭUV�|�ͩsG�Q'W�4��-�CU���j`��G��m��Y�����W�<MJ�i�B?�՛W
N��CB�lI�������{�p���<��t��:�Z�,2 +�V��m�Ѿ�Gl<*ݹ�U��@��JA�q�j�=Z��[dב"$���7";_��4�gB�,;���y���x+��3Z�g-m�v2*F�(.����/���ꌉ���߹�Z	�j'Z��c��B�vA-��gQ4��N̯���	[c�˓��HB�I�3ud�L����&�5�xV��2�t��U�򼕯>6o��$��[�cfL���������9ӫ�����hW�R�V$�*���/�a�=��m+������r�s_@@[�n�V�9ɰ��s��i��>����v~7�[��BIٹI��{�����B�8(�$Ug)���!1ަ�k��۬�����5�j�g�_�h��7�i��
y��'�oUA5�YT3��;L����W���Qs�tx��o��k�H�2�l��fC��~��s�o9��ӽ �_�r:{�����8�H��`��I5S26�RO��ֱ�ǅh��ʹ�D��C��y{�!���0K�-�(�}@a�
��a>-j��-|шVg!��h���@��~8����y��ޥ֗s ���	r�Յ���SZ9���]�W�c��=L�Y�H��|/ȁ���[H����,%󘛆BC(I�2���m�.�|�_ОBj?�O��t�ݿ�+�i:��i1�� �2���B���/�x�L8�p��$�s��ʖ�!VS�����O�LrM,�Î��%ْо�i�d���U���y��֜~h�}�����as#����wj� ���|%*��p�Õ��T:�eT�[�uJK%�p���~q�� ݐ֢e�У��#ݴ�������&E��C�[-��J�s%4�o��/�����i�$�rR�T��M�_:D�Ț�y�;^h�zhN��L�J\�޲y�>&��Y�[X3���?�O���$5��b�ث�6ffe'?�-�in�f�U��GB�L�P���zl�]�6Je�����G�-�7�ɺ��G�	F�?�}"Ҹ�]��gNW㠤�B�Y��4�pP�iVIz7��0�������'iCV��eм�6-���OâcG.��Fya�@B9�V����e� �PE�DP.K
��:ͶC�۱5���@���QqF��- �(8G
D�(�S�<	�y�w�g8�k�E'q�&��h��AjU��5P �����
IQ[9�'�$��������g�M�P�������6����x	C��d!
3h��<�gqc��PP^6�a<,�eTJ����� ��.v.4��k	��ii���w��&��*�*h�rպ��a�{�o�3�b<���[�%�F�,����+��K�_˄��\����_�-�"�^-��C&��
�%}q�a} �J4q��Y��B2'�ak��h���¸P���&�ř��L튽��g���l�="K�̓�g��O�`G>��Z��ByA���2��I��:�v~��?�� ���Ʋ�)��q�q;wi�T��(���&M�s�>���)�Гˆ���������c�!uPc�zsi��C&2�a���Z�QP���h����ϼ�o��&ǜ��Jw�le͒c�z�*��Uv��®p�Q���ό�%4�ƻF�r��M��0�K�@gU1	��۱�Wf��h�/�࠼
�5�CaG�K�ܷ�"��� �c7%����KF����f<���L�����N\�I�������������C[L��Fٜ���������{n�ViX%pc4.٭��=���݆?�p���Z�ȵ~�����+��is��⠕Wď�B��3r��iNX�?� 4�h�cikWC�I�&p������qa~��!­w�u?�H��z�*X\Ia�_'��1�_��T�V��5�9�
�Kâ�VX�?ɼ�F$Gp��S�hO6u6,����-�w��'"G�5���?ڢ9��ڗ��t�N������T�n�r�� f�eݑ�ˏ����0�M���.�h��F20A�>�Sv�ߗ8!_�(e�(`T�a�?)Cc��q7�����M�l������ʽ0YD�	�&n�*Y])��+��������E��U�N�L��U����/M��|�N������ٌ������U��]4.�O�`a6p.č��#�g�K�ܝk��`e�ƽ-�򀈑7}l���!�����[�̯_hVo,j;ڔ�����+���ƌ=;����ew�z�;c�!�rg����!��]�[���Ʉ�Tk����*��}KK�E��n},r#Oy�Q�<���K�VމL�R0@���Ta�O�L��7F�	W*���y�+�ؠi�)�jAo�d�j$2���0�z��^�XO|B_U1���������qY�6�7R�=<�$۷���%�Zs���������DcZ�_��6 �g��w���ȴ�s�kً\e�2���}t����I!����>j���� ˸W���_>,4���DsT��e�u)�+d�Cv}�7�i�hZ�6��&듪�?��$�V��
/ L@�"B2�����4�qJD�%̨�}/�w���)0�Ͽ�b��)�%_��*�Ďa��Mp��B
(P�M $<?XQ������c\�&P8B�]��\��>C
d/%\�ݟ������^��@��4�[���7V��)ń(�G�:
/��.�z�m�~W4AoM<���RD�UyC$���0������0'f^:sj�]Qd��IZ��=獷l�M���h"���K���A�g��������@a[��-Bk��A�x-���Y.�Ѻ���3�?~��6� �	u�VҪ%z���mD�H��F�@��^���1V�n��N'�,8f0� =ԯ>�D�"�osn�~<�����da�bAF$2�O���ԉ���.�E9�q�#�;$ޑȚ0i��;R��T�:�3#���5#j�v�>Lɷ�gn�Va��Dt5���ٔ\��@!]����u�tL�6o��"+F&��i�w�7b�*A$�׾����0��u���Jq+t�f���C����k�oS�]?��C��$Ȭ���iöК��kH�cz�\��p����b˿�N�Un�<I��2�����<܆��8�:�6<���W*�� @�S�25r"9��Ȱ1�}��3�N�����n*h�sn��Y�y�$:)���U��g����%��A��{��h�O�W~.%���Fe�����c�
ۖ.fS���@ AZQ�N�}�	/�Q���B)�&ݰa�D�P�_��P��銋����$���5;]	��9���}6�ĉ2<ҝ��0��{`�F5���3q�(f�+;'���(~<��$o�W��]��I׮�ΠZ	�#I�'b���Yp��$z�pH��� gCr��N����g��OCcy���@�]��;����D4?��}f��X*"-�������{Hڤh��� �~pA��᝶m�hW��M<i�3upJ,x��C��#�Ø<�����i;P�������d��Qt��>����B8m�]q����I%�>�%�RĔf�nEM��gK����P<k�GxQ�t�)m���c�aaJ�hi�9ɁKt��+��"�H������jOF-�y���U��!$u�i�ޔWUJB�b\��]YV����j��uAi`��=��Oj����U��B�-޵]�L�J�w0,�.��,�I���j �2dr\�@�2W-I-��BiOˊ��)�)�N`d�kղ��=����68XX���?�&k����6���}(��r��h�M��A���'+��nq�p���aT'�|�l.��ڍ�v`O,eБ������B�>�(<&o�T�~3�S�!K�&vvej�$]o[��8Z��h�\/wK\ �؀jI�hKs<��;��A��R�b����~(������߻��ފ��2���g��&�>:ș�b%�q͖��Ւ�~�E�ZM�����a�u�^ec{����æ;j�!6��>���0����2�Ө��ގ2&	�;Va���ٕ�pFo!yԧ��M{Ӟ����n�N{�2�U�����\��{��<�ȚqQ���y�@]��t�q��*���^p�A�H�ٯ��rݕ-S�//��qVꢱ~G�ʷG垜���+��i�r<Uw�@���u��H�Y�ެ
�[��#Q[��P.����ϣS|&"0��!b�hNn�	�� �4�a���&+QE.�b��L��~�;LzEe)�X�8�����%��s�k��s�o�2L]��2zR�)��
��Ѥ|"Os�~�&�Ѫ,+�_�N��a1T �ʌ8������f�ݴk��'F��ɭ�R��I����7[5^�肃� ��#�'��Qy��O&�R��O�F�X��
�U&�[F����m�i��/��\UT��s)�KüQ���i*�a1����3}����r<	��-��{�n=i�������=���̞/��� �7ҎN���`Y��f��y�Mc�x'1a�fӭ�f��P+8�zZ`Γ���S�����[�(SO�(��� �Rj����R�o舷3�5$�ZM�p@���-�c{)�(��>�Zq�M�5����UC9>� 6�X�|G��'��^Ny����i���O�ħ�����OG��%����U�C����49C6+�q��C?]������H��cm��[;zLl��zKG*/��� �uN�� <Fs�yh|
[�w<�1�	47��N�����A��x_W~\qR.Ꙡ
�Z���pSQ���Ϊ��\�HI�����u��#�3?�W�^gLn�
�߂W�2\OL���=.�%k����c���ں4�a�Ǟv1�ͷ���:�B��7+%��i
2 �|L�rPV{���.)�N1p�Ȁg4��qJq�t��N�8�������?\}>�ע�?���#�4E�1��ڰ�i�\xЛ�WɈ���qZ=K~0A_���7I��:�3ν�`���1���$�u߆��ʴdJ�_)�io��	�g���S��HZ��,��`�&T�0b�_�*�?�<e�� ����Ң��xG�3h}Qv�Q�T���ޖY~�c,�9���fnuk�v2f'���Z�[��\�%�at[������9n��:�h�g������*h~u?��{҄ь�m@0�����>���>?x�+
V�U����	G��8P�m�&���8;i-�g�Wi�a�Ydt����8;�D�M��8���xu���s�L3"n%UO"�z�jBf֗��jXQ��:œ��v �Rg��_����R����� �r��T�:�N��;��Q-�9��Y�����]no��\��w��ސ�x�f?���OtY�k��/E`ne�0���BE��r�a/	����{��5����@����f肪��T��X���W%�/]�۶��Sh�]f�P��OZ˔}�`!��*�y��~і���<�_�U�cB����9�pj̹���iz�o$����E7�+����ʽ�SI�U�Fu��O�����x�^�<	�^2���ښτqV�M�Q���aT�l+D�ƍXu��	�q�QAq�[mN���t���9be�7�<��3?�c�9���\��ȅ�l��d���1��4�{؆T��'��s��>6�Ȩ�ߌ���m\�?��Z�J4G+�*|�L/�ߌ��H譤����U�T��+�'���op����E��jSzᚚMYj~a�7\�v�r��H+�}��|�2f��<�������ı�Km3���X�X(i�
T�/:nFh��l�
�H}�K�m<��	R9<��Q�=��f	��)����@Po��P��XJY�X%�3�m>x2q9�I���*.0|C1�u�X����B������ޜr�a���}�b���ik��׋�?尐��;���7�At�tl*.w8X�3~����!��h�(�����P�a��S�g�p�Ŋ��n��<d�� ܜ�c�u�w�{D�p��"��7E'��JA�Mǆ�R;G#�T��H��~�C�35���+y�q��D���>��H�Fc��M��$�2�ċ���T�Z�������a=����_i���`�VDU�獟�/�~�!�.{��p"�M* �=�2 TU�V,H����S��[P�߆�,�-r�H�(��-��P��>�{�@�������y���od"�ӘS	�	j bM�C4
M�<����ޑ��C�a��:��04���&�ۏ^��ݏ7^�jQ[��̚[Y'+޼�"��,Ĺ��3�DJ�3u3���In���f�e��P:��2F�=�'N�Py�wR.x. @ >l��Y�B�+84K߹^J{����,�M�:�`S�Ts˔�de�]^��&$�N�1���}�D�+��:�[]�������� $��+��/z��1{A67U�qK�t��gI�ds�OI�'k��nỴt����.�G>�߯X��Fνq`;ao�cSQg��V^A�2pa����f0A#H������6Z��`�4c����U�������]�i�F� ���ۓq+�|;��QI�2�Y�قI�<�?��A|k�傜��ukJH��uE�^�פ\�`�b�T�!�G��8Y^ ��!ߊF-Ԥ�ſ�� ��!��c�^�ē�}�	�^Q�[���tG���t\���'����E(�z;��2CB�ڥ��b?D�=}2oy��Vze��'S�d��]���SU֑�h|����~dӢL�7by#���g=��w$	ht����U�ń��"��0�]p@k!iQ���,���8�H0R�F*���!��_f~���5��'��g�[�S���"0ӝ�<��#Gh�G�ʃ�w>�wB�b��{d�pO���1F������q8�t dK^({�Ј���S��X�F2�'jKN���a4LdtM������U4J�%�J_��˱�<�X��yy�B`�+�8���@O`坛��˅��$b��d�\����z��tbA� 8�I.A�^p@s?����M�0
u)IE��D��F�ٰ7>�LJ�mqz:[\�q%+iw�v���Y_�j�ګ�6��)� �+��2�r�0�m|B^'lPԖ�?�Uj� ����zy�Xq�-����.�Z��HQ"3�W�F�ܾO��r-w�h��j�� �Թ�^�@
��B�\��D|��j�۔R����!{�\�����+�tA~�I/��>�P��x��%��g]�0�i2̮�a`7;݉陇L?R^A�BZ���FZ��u[��ws��z'y�i�0.,Bp�A�0���7V����d	�7@��KH�Ϋ������YKM0���CH��sN����ʣ�G-�[��<Ҵ��� 1$���t���q{<��Ћ}C�hb��0n*�(�6�u��g��\}e���R�R"�>c���c:{o�*�S|�AW�Pe��:
����z��Rg�DH[�5e7�~�u>r�/�](���w���k0�4��KÏv}����7�W5x���-���g<~�O�h|/�Xx��Kԗ���^0��Q�w��[����Y��tRh���_MZ�����`�R1��@F��C�iy�l�a���eקyȝd6ٕ��RJ���J
�`��@��z��ç5��,$l|چJt]�sD��\�3Q��n�Aeۓ]!��N��C!aY�C$��*�[���O�Ef��~����+�ɮqRڌd/�{[B����rê����!p�� ZC��d��0{>�S;��@�(h(�k&��Ь,�Ħ��v[	~��N��s���J�+�.�ݸ�v<iɈ��Ot:�'� �=�/_$�/ho�e�ϼz��2��sp/������d���,�t��|Q�;�OOD�9��m�����	c������l����^�KѪV9�Ҋ5�Î�&�X�ح|R�G؆M �w ܈��8J'��p�Rg��5�"�&|��\�t��[rJ�w��B�'�ݴ����g�}.<U,˴�nYY�eW�����UU�;��]!����wy�v��5&<��#�Ap׾�N���]=��Hzc�7O��X�N����)S�a�	��-_釲ec�?���������P��>�[�smH��/[.OX�}8�p����
���4��(@Q��x�:��4_L�9>�4-9�=�˽d�j��@`�g�{�+�G!1����R��I�
�fνu6�lV����V9����׀ �����K�߿���<!�wpl�䪝�2���o���A�NQ�|���8O�V�$�F��������%���^_@1ץ�Ԛ?�){�xA@�s8��4��a��a���N��DP���So#�����)�U�����A����F�>�-3�I��!��6�DD���=C����9w⼀������7��:챿���k64��n(L&.|�����+O���*u�ʆf�_��)6����U�a ��e��,�isy�`��0�����P��\xX3luE	�$���yV0�m=�^.�a��EJ١�e�+`'���b���"�:�	�)����O�%����� a��N֘i�����JQYz�m����3��#
[YfX��v��g|�W����K�T\�좪l�;��wxzB�?�IM�����C���߃�7��"`s�|�0%�J+v�}��I�\L�ܕh�y���_�"���3�8m�ߌ����T�]���@u��)_1:_uhy�G\2��t�09��b�9��V��F0.p+�	x�SW�S�2U^��L�������S���c ��M���oSo�f��E���"�8r��E�GDE���W��`ShU}vS�"�r�Y�ߟ�T�_s��߹�0���j�-Ar^���A#�/5
��Nid׊^m]���>\���Qj�]$�Nܿ��⊆~��/d�_?>�a�\�#�e��5�Դ	k�0�0�엸b�
 ����0������u<��c��	c��'�6�����d=�.AZ� OT�����%���I�j~{�M�<�����@�$�W�����A��[�cN��J#3��YFh�����Ȱ�Y~�nGCh/2q/�hr�lzb��X��ݒ��eC.+Q�m������>촷��m��H�GS�$�M�%b����VI�l����qN�9A��A���=�\w+5�u���Ȇx섦{-�P���`3 �%��W'��Xp�K�e���&՚:�Ч�-�l��sH��&���c`��-��3 ��J+�Hm�5�{�lqi?��X�l9bV ܓxԖ���k4���=��2Ⱦo��2���ߨ~5_����jA��®���]�~D�Ƈ�����{/�,��1lO���O�mdk�+�	���z�/k	���h�����8+Yg�΍�4*2��Gۯ8��+��)�G��Vϙ6r�m����fGq'*��Z�!���ֈ�[�Ƣ����{>�����J�
a�!S>D� �#����X"̥�S8i7e�$��Sv��_�w��s䈍��ꐞ�n��I~\����KĜ�w&��G���"2?I����t~����mԄ�
������>Ђx���C÷[����-��m��һ��|6%��g=Ht��bg�O�
��:5҉���O�7(��԰-0
Q��F��DDX��JR�
��u�Z=�{ٌ+h1����!ΟS:�h]P����.B���/%lbD���O��8�+8�by��4S�?�
s�}�>�A\�i T2�� �kc=�\�L*A���}Kr�"�{q��߹T��)��E���h�Af�]��F�P�����q���]~"an{҄-��IcԠ#k�h"�"ʇD!~,�)�����ö���Lǲ��EF���@��6:J��SU�:]��}���
�Y�VYuj]�G���wC�ly��U�"��ɜ��b�!���V�"-�v>���:�}�QA�j9���r��Yˤ)e@�|~��X+gZ0:�0hQoO�][{xf�.4���4w�$�!��g��O��I��@20q�B�҂�~^����4�|�n��&�1b"�d�$�L���GL�H�]��#�nԗ�n��$�~�Ү������s.��09b�>:f� ��;�k����$:��B��m��Ν?��7�˛0]ݲ�X4$���JJ��v��*�ꌯ��]D�A$H!�W_�v\ULJ�Z"�yS#��=<ކ��|��j]�p����@c� �mI���������$.�Bl���0`�Q��w#���e������CmK��+l�������SUcj��I�-,�W�ĵ��m����&F�5C�=G]p_*S:#����؄��`�
����YQ�)����"[V����w9��N�AO�����L��]��ɍL�)�MOU�	�x���i�_d��T]&�� f��k�~�c@�P��7
=铟��3��)ӡ�����[#�4�1X杨�x��W՝���b8�}�P=jIϹ*|J�b8�X���1:��Ik�!�� �)䂥jr���30Y��n5�� 	sr�tF�E�\G�iv2�N�S[�p�ɲ���uE�੓KQI�7R��g�ܥ6m���-�nm@�4���@t�i�_}�N�6�x����vx[&���C�s�C=�I��0��Yi[$����FE����uD��ak��P�