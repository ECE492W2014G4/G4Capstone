��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P��v�"<ߞ��&'��k%P碶�R�ӣ�sĞ������FY&i��qzJ�Y�<���f8�<FN��G�����n�|�4r{M�^D�&�p3��'=?�B-ƍb�n� �*CU���p��n�\�P��s��;�W�6a�a!A��	!�k[��{=I��F�#|��1̩�5W���"����TG+�aㇼ�&��j�5�P������'b�^��S�;f����2x��/�t�Pl�qZE"��Q �b=�޵K�;�ƌR}�<x�t3�W'xl�]�*u��6��氭��|�>O�o�[v\Wq���;��P4��#���ʿ����徻ySD�cSD�p�r�R�ج�:���Xc�M��YF��VCa����c
E�x"�مtݕ ���prݯ�3P�)����X%����v�t?
'7���O�H��;��Q)n���U�9���ү0-��K��H{��՛TC=���g���6֧k�u�3�/Q��訞��:��ϴ�e6���\/��4�r�n������tH1v���7�����Sw�T�p�����7���!��.�8�n77|���2�j�Gf��~Kj2���r��E�*�P$�ݩ��|��N\ �O��钽�VXϸ�3��Մ�ORlE����#O�蕪�oG�0ߦ ��_kPS�	C�|M�Jn���E%椱�C��S�Q��ƀ�b�d�>�� �u�S2�� �ӏ�C�S�� ��.�%BmG|6�j���.7���k��R:��O��ה�,���x�����6iHR�c��
�F@o1�p^h�P��/p����2�Ţ��~冶!��X�"�$b~ePA�Fxݗ���M��i�$��3�X��%��&�4o��T4-H��}�QNǘ	����%�6��wW7�\S�/\�O����1��/�H$��K��&T�9.ف�Yh�sok��H��.��%�E=\L�\��T-*�w�RΡ��������7��e<�>F�����M�����/p6Q�"Ry���"�µ}n�'��]2�DX��7ٖ�	��:qpx!����YDa^�\"&���K���.������/�vH�I�e�A�ÔOrݫ#g���<��v�y��fRB�RR��Zmb$X����\2����V���Cy>���C�iD=i3�p�'�t|�&�y���R궿��wN+G��w���lz��ݽ|
N�֢�A��l/6G)����>�#ߋ)���&��g��,˞�%T�_�ؑ4w�7ˋmWJFB�� ;.�����d}z.Rv��^Ɇ�*$�
��T��k��F�����N�!���V$� ���������qSW���o�.�����Rĉ���U��U���u��;}�`C��M���I�VÛ�j��S��/[2��7��s��]t;��[$4t!�Or�M��9����NGy�/�}�5�|YT�wz��1���ݗ����A��u�b�7�Ԟ�v𣏕��j��Rl�>�p���nX�v(u��wN���㭙�׊���v���?
)��;0��o�0��)g4�b�9[`�����]Yv�ai�Z�q�wU�r�����[D	P��󋨪�1�����r6L߻n__/�Ǆ�J.dkR��'J*��M�2��UhU����Ց��l���{���3�G˛�`�B����X�+2�)F_X=��۠�̨��ġ�Y�-&Y�@9c�lTT�zb�¬MъJ�|(��O�P�=���rSX|�0�8xA��5��X��>�IbܪE0��x�N�D�(����~�~�\j��yfbz��R�ӹ�kʘ��G8v�G�3�V�8��7�zs��J&��ˣ���^��(�("a��'@�qz�J��?E�U���!Pa��o ���H��,��8Qz�/z+zF�|�w�UV3H�<A�5��ճ�Q�!w5��$Z�D㝺��1,��
3���J�0�+a�;�����[��a\d=t2Ix!�� ��V��S]�
��:�k�(!:�\�@����`g�
93DC�A����t�=�tA:6�U�}Y�����ǜ=�;\vG�e�@|9���Zy��Q񙡦��@iV�=]�խt&�,��ц�\��6���J���Xâ�ݧR�B�\K�xusB���\�ӗ\���c��9���Z�j��L�m�K��	]�_`G%�w����X����p��02�.�(���~%Z�K{u�x����~QH�d#\A�I�	��݆i�9¢D�������i��hG�X��+��_u�]�[-1�B��wC��>S6
Uu�}
��9n�İ0��2;b��{ b�(���6�_�¿QG��<u�rj����`1�Ns�j�8(�@�n��[�n���6q�ˣ�(<Hi���:ej漍��������17e�9%�}�	���}!�h����T@�JBƑ'RU����I:8�S���u���k��V�dPp�!�ǰh�Ğ�)��������Y��������Da���H֕���w��o���Ƞ����EY���X��rn����Pa�b�@��r�os��:q2��#��MM�X�m.�[Հو EC��]����
""�DR�����C=��R��{�DE\ A�����H|
�,�,�p���@|d�cɱe�֎y����\��p�>i�7�y����boP
���a�g�U�<��� �^������n����f����%���K<̷	`�Y�'�%���U�ƿ�	8�	Kć9�O���FK��~R5��������<I�����Vs{�ȱ	Bϖ=�������Ҡ������6w
#f ��B� C��e&h�ő���m�]��T���	�FL.���w�a*��pwJAOF�D"�K� �"�������<}�"`;��WA���	^�ӿ���6�s�,���&S���-$tʊa��Ek	܀�< Q�k�sg�� آ �ҥ�:p�#�ؑq�'X������5�ƦcrK�sn�T.�;|���Ҹ_��,�$`۵5����x����/%���}6V��c�=�et����C^|&��x�j���1οRڒ%��?�
1�����wyQ�ĝ�+�&���"��{�N����s��D�cJB��P� w��4�
'��vԟ�z�m��8��N�൭�J	k�/j��+�Y��.V=j���.S�$Fe�G�VC~Bv�C!�>���Hd�0_7u;(j�9�k��f�!9�����4l�聕��x�=ꁂ`] �w��.WQw�3��y,@]��I'�����,l�/��Y#N���cd�8��^��^.�+�9+�Ŭ-e�SЎR��	M�+	�3�Y�0L]PP%5�x�,)˝;�����������z��_NC{���ט~Xz�VZ(�v秼v&������e�aJ�_��ٵܝTeWf_��8�Fp�tw�A��a�i
�@�W�@�y���A����9/М��Y
u�(��x��S�[��`�?ߥX�=����x��f��ZqZ���C��/��<��gm;w�\��i��z~�:=hh5����Ƒ]��Ӈ��5���sZ��t��i	�ۧY�h��C/z�|�+�1[c���0��iӽp)�޳0�,�H�������d�P�z�;(@oڲ搭����[Zz*�C�u=�$B�{�D�dCo���%��Q M�!6舂���)�"b��!�,���x<�D˧���L�+t7꟝��ӥ�ߏ��T�+��ON�}�Ķ�2��j��URܟ��F-��lp�"� Ίɦ������*�ѡ�,�G�@��p�J �E��oi�y��:��e>�I���TE-���g1�F�0��]^tJ8����hz�)M��j��|4t��mV���<�hoo=k��M�K�R؝Y���s��	��G£}FU�O�L)v�'��>ܮ�9
.�_���T�7�����)d���*�I��u���T����/�ۺ��"�{�ٮKX�(_��I�vu`tx��ᵂ^!�7�� �&be�1����?��܊�1^PU���CȌѳ@��v����h�a���A]q�ip<�Lk�m����������p)k�tv/����[�����`?��ۋ���;d�9���5IUN>�?���`����Ñ���m}�>ym�cQ���9�?S�	
d,�?�k,�I՘8��m�G�=�M ���.��j�����34�,����Y־�=������;��攊�g���I���
$��l�/��`�clHe�vA����^�hASM�?�ŝ�G��߻�5�8��Y�*����w�,�Y2���o�eS2�(�T����E >�UI��}�kH\
" g,M�J��+b|�s�,�x=L�aiQ���.X9�8�fVf�҃X��{������d5l~�֟�b�YB�x�7lr��AE��9�r< ��"^�U���<�8��Y!�K�������ה�҄�()��Wջ�yN��� @��x�屶��w:��1ןǱ뒙�X��y�%.!���_�f���/Z1���J:1�6��5���ۚb��]o���]�!{N��*��\�]��cՙ�����b���a=2� dax�M�CW;{��Q�0k�����oD:�X��>]L���ѷ����p�{��aSyQ� ��M����ۘ�l$&��B��������%�j�* L�<�*��b*Ȇ�<�� �s@�0~t$� ���N���#=F6\�]e�Q�������yڼ��8-E��^��{��M�tծ~#Y#i�X�S��@��̄'�u��=��|���6-�}Ԁ�3/M��̪�"B2�i�J�,zW�rK8��o@�n@���J���
�K�?�j���`m�4I�n- ��ٚ���C�V��03�A�O�[����Ե��,��R �>�T�8H��+�	Z�����%��͂W���~�����
F��K݊��U+��Ӓ6��prU��6c���U��ʢc����J�Ō0�T�%�,F�l��|PK�)^l^��h\�(l<��堢��Xer�6�hZ���rej���A�F9S�^(�����io�_mrVz"С�i�M�< =��P6��x��a�!m��8ƻ$[Ұ�
��`3�b��@��lN��Ũ��V۩4t[��g�AAʈM.!�%�a��u]d�s3�qF�kpǢ�J"Q%����Qs�mK3�`!�ZX��H�&o���州V�蓮��^�!����xM�=�K��s|
�&���g�t�C>�.���y��DG�=q[T�VI��2Cy�O�{�D6�3HC���Иޚ��VBD��	�H�yH�����q����7%S��f6pA�2��:��/ˉ����1��>~�M�4�����vƚ�c�߅;���x�[8Ujo����0����m�����i|8nZ��ùFx�y@�	txWq���\;u�i�J�r�av�C~��/4��HB�{�LR�ut2�_C��ng�)�f~Z
�Gz<��O/_P���t���K�.V$ tn����faV�R�ճ�ٴL
\�U HK�PÀ=���^�r]�W�mJ�gn)?/)'�J�]C�Q�����I�*�|WM�Ɩ:��6�mIT��<����> 
1��^��A���1uK t`�ݧ��Xh֩@�3������^gzRrk������Ŋ����^���������?���+^�<V6eۺj��E+PN�'�	��6��Z�q�n�ք���LL[��Y���D�{�k�j�K3��kRSN-B��C�K��j ���.�X�5�=��sPOv4�,<	Jt�FZI�R��!�h���MpFS��d4��w*����5��>���ʇ�ҷU��.P���������C�iTf �����顴��G��n��/Acj���Upv1��,�y��?