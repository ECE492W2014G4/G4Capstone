��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�"��F9s�`&���a�oq���F�g�O�]�<ݲ����eCL��D���{�5��8̝DFI��Zp\m|Q��
�}�6C���UnF:<�jΈ�2�����<����sf�k��,jڙ�����2��X��Ss�HL��	�������+g?���N�Ż�����|�v7�{M��VNB
��Rs�゙�Ld\��X�'��R :�J���^�����kMkx�Q���3!P}�e���Z�Y?.�U{�RP	�)��lI{tI(S
7ZF�W+h���ګ�jc>O�(�d���2��M�J��`��Θ�£@���~�2Q5�Ҁ�?F"�������m3*�D�dD%���Q��OEB��rn���G��w�3�4���L�ఆ�_�X<�cgrEf2f�2+�цO�dyǘ.�,��OKF�^����q� ����IQŲs��U�&��!�  ���?G�=��Y�BX�	���2�̀��\	c�Jk�F/̐N�����ҧA	da|��`����\TQO,^4�n�^.QP��0*b�� 7>FZH���~��,�^:�����Y�S j�|��ƻa�\�iA�~�i1�@����,E�7��^)!'���<7a�o����V��;��2�'5pV��3R^`�Z�Ë��ӆ3�h�� h ����kr���iHi<V5R.�X���9��՛�FHI�`ԐD���Wpm�c���Mo�'C>:*�dU]��,Y��L�܋�8��-~��1빮ߕN���qݺ��;��?�f��N_�`Ψ�L�T־�b��ؕd|Q�'�tGI���c6�Y�4�������[Ɯcp��,�2����+1�+ё
�y�Ƀ7����?��#m]q��_� ��X�+x�XO He��8ؔ�F~�b�GljTX�>��t��؞�E�hB�&�l}9Uڰ�e�������T��⭘П� +R�S��+�t��~��0�L�aXϢ�N-H��,��Ty4���S�J���2bh���/"QOi	���16��y	��d~۵�*bw&0�/�����1�5�aa��6\ɑNt=��{��E�f��7kx�������kJV����-��	�@�Ә�UU̶�j|%�џ�:�'�D�M'k���7ReeH�Pt����D�lW�Ҋv�SR_���� #B:D��7�`s읈�J���Uę����,e�/Klo�Ii��tW���U�����n���G����?�w�޼��`������G!�R�L�1ϒ���`'��:�xNˋ�nV�ڔS.|�Ve�H��J�K��6����_Ҩ�����%�I$����hF�t�!�l܊S� %!S�Y؜e.c���'�Knnв�r����kA@��,��o�d�i�`�V��ӊ�U��9�߈�&b*UJ�R_M�r���(Gg�E����J��z�25!��a��d��:9������2'��`Н��5*[eQNl���N��+4Ϙ��Ǉ��ߝ�W�]^^~�."F�8��j�:d�����V"!.�|��Gگ��y���\n�5R9���o�52�U����K��@�Nr*c�Wy��+��>��ozQl�$a���Г��S���#T�)ӹ������e��}A`���� ��0�G��h9(Ҿ�Z}�E��$R5�z>�8����Z��0�U�sv��_����B�j��F3�@r�I���ϱ�3�P5��v�'��"}���&n]tZǲ'8ʫ�W��*Tћb`Ayyo�?je�a�����sg@=ɠ-��P��%^�Ǫ���ט�P��b=ᷲ��r������1��@�xWH���L"�q�E�#0^~#Z�T0�Yc���,�jK�R^���PH�[l�#,�o%�U�|�q��岾)"� Y�;�>���)U��v8��Ɩ2�p��8r6i�����G�i��6����,{N��*�5�E%IU+�<�h�w�"�t���\J�n�)�����uн��Y���_m��V>�v�ȓGP�����؋�A�5�#�O^<-��i�}X�gb�d	cIV�F�g��m�*Ka�/~�@��q%߲��B���ŧ����Au��
7���ic]hq��E$#��Gx)�˟�8�ܗÂ ~D<��6L�����R|-� ��s<y�k�VHXT�%y.ϣ@�GB.6 ΗJ����:H��'�2N)p�Guš�_����Z@��
�ZRu{��
0jʊP���̑��Ϙ�Hϯ_̣�K.�M։T�C �I�d1���	�?�s��{<�g.q�q��?D
�4Yp�%6��#7��2s��1ɳ���\�č�mn�aF,E��Nڵ<����gi	@	���R���Xح���w�v~�4��KIy�xW��g�{����*r	��1ql?6X�g�s��c%擾G��~��� .� >M��b�IHc��.`c�gɩ-�`�	AK��p'R�ʭu�
o��K<O+�H�)J�mT�9�.��B��I��ce�e'���8�����l8w�0"r�?J�/'
o�2����=�P�u�Q�}���R���C�H<崓�����:�����>5��9,��n�����R|��A�G@C0w�}�r��c%兢gl�Z�F��v�S�9\���~�
:lB[�������pEx_e�H�D^��IO;����OU�|=6�h��%���D��%����$��L���Q�5� ��V1D�*�r<>�?oO��p)��&C��&�����ga^��uá�.�[�D =�0L+�١{o����)��W�j]W���<��M���C���i?�i��� �����]N�0�����Zvv��/����:)�4٢��O{��H=�oFp/������k�{.s��V�w������P�8�#;e�)X���u�Yӧ �w�C\��0�L^u>)-��.!F������Jn���dן�\�$�n���P�)c�=�2hM������U�N������rxSM!�j�R� � �N�@e%U9�4g��מ-0���&�u�����3�O�o�1%�Uĸ{�$��?��Tb�(�ؿ�K���J^�n�g��ϗ�Vv�m��)�%�ԡ�sF`�@�
g��Bb���G �>��������߼��Ȋ��t��u�F8�c��Ls�ך�w�u��l��$]�$ꫀj�$�I�[��X;;[��5S�9���JtLvO�0�T��.`���T=�E~�U������X���=�6l3N4P�T�L�I�e=W<�VJێT�Q��+�f�v��f�@�-*6N�L>
���v[�MP��W��R���:��i)Ci3m��3л	s
?뛠�(�f~ƌx��3 m��,�%]@����c@\|�`��j�������13�&������6��'�)�8w+G7�@����y��o���p)F��`�U�@n`��{�l9����~��! l��`��QD�1x'��*O;�A|����CnR�i"#� u��fZ�}hA�I��aEN,업�F�s%
��Eo���2)zM�.�����N�-I�������yNH��˾qf�m�E�������a�=�M���� �*I&�R��Ŋm{�~>��E-�ۓ�� ܝc<�uM���+Q��{��3A��Fz����@	��QՂ�GݴM^�qw������eƇ�u��o���|���^���C�S@������\'�}�g'��\��$K��;��J��9���v���(dLJD�)�IG��>ʶ�yĈdyq��
q\d�{𐐸�Q���D�>�ܦܠ�u�l��e����(�*(*�����uc"r���\Q��&Ӗ��w��Z|d�f#�B��j!��I���;�WD��s�c������f��)Ϲn3i>u�$2���̵�?ݿT0����4[D��q�����q��!��r�Tn�����+/��$Գ�@�q%�\),ڑ�)��7�d���L8vb�듌�xx8=#aS�����mU��&#Cή��;-�$�p&j��]otl)pNI�;���w��}�fi�6�Q'����Y�H�-����>�fX��k�@�'W���[�����q������>�$9D\^��x_@�1q_U���pt�b���Ǖ&��U��挑{i�f`ԍ[��)�pa����u}�^ �)����6�qJ8�lc�M��*�3��-?/��c܃@z��ƹ,�_��<��n��\&7�7t�?�ە�A��Z��I6�IG���zq(/�Nn���l\d��M~aD��N�]�nX��yq+�#�v^v񣦩/���kM��F�+,} �DuX=��U�n(�Vk���M��Eq����������˟��w�N�� ��&D���W~���|����)����R4v���ת����?��9-n>q��r��W�fm������\��	��GA��,lْ�,J\��rd����@ytqj {[����b7�s��\a%D���Ѕ� �������L��j��C�bq��8l6�2&��A��`rI]�ԕ�F���_nL2^��I|(��]�-����v�(8�2<�!Cҕ�<��ގ���d���ZH�KFK�X��28O�Y�p����eϲ��^U�?d�>�ė�2
��Z�P�BM�A�M4+�{�N� ('24U��ȱ��MP������Ah{���ty������M�O��W}Ü{���%�j�lR���wq3<�|N����>z�E�T���e��`?�.�=��5`��^�I�m=D�Q,��ܨ����	���0��̫5�v�*7~�U�p�����Qa%�:���Fz��ELh���;��d=������@�����)N���������GSa�˚�dߒ�݉���O�B�T�R��LYbA@6:����)کݘk�Z�r�0e�CR���3ظ��*�;@��-S�h ^}7�*hc.<��q�"�>#����ua�r���#AqB@G��;��cU=�+����{utXn �L��^���g�g�PiQ�����;�n2��Ob���ً8N���:����漤���{������ ʌ����d�c�{1~��z�P<QN���N�
�;�����K�w����M�BtvMl#�1$m=��r�j�*'��Og�&٤,�j�*C�#�I[W��=BQ���%ڀ���v�^D�\�=VN)�D�xq�����)]]��f�B�Bި�J��q��V�I?�{-�[�0y_��oҶ�Ѿ��=�{t��1Q�+���@<Iu��63�B�lm�����jYD�3���݃z4����ǣi�.fAզ]%i�������kq3�!nę�����3kd�Js�����C�֣�Q���+b�ޓ��'�u�Ax\�]b <�(�50���]%9��B�Q��$[;��ή�$ɽ�h�ۖ}`���%!���A`���t�W��j���_O�|��I��S)�L%���-n�C f�`��b���#J�sL5���?�7���r��f�)*?�)~3��כ�Ӌ���/c��������ve�W�EqD`m��³W�w����Md#4q	��ܑ�v<e5u]ћ�Y=R3��21� ��
�)@��4;���#��v��(�\-C�-\��H��v�>u�UŃ���p�3��`=]7h��k��� P��f2���%|,��CW��!A'	L��l�~gL,^�����+��Wf�636J �P���_1��;���X#b�N�͝�c�}�`��9i�BS�;?
�@�5j=*�n\;��������&a�y>���ٹ�I���S�j�c2	��X���W'�\$�.���Va�2��9N>ͮ"��ğ?�so<��%>�`E�S��.����A��[	�*����.��=>��@�4�p������v��u��w��S����@�/�#�s�$�53͊�4����"��l�n���uw
����;�="��l�~��T��ȃ�,�E��0�1�k{�j�&����S*�����	�:f�D�L���(��D����uU�G�.��jV�IX�o�&����v�l���^X 3y�Ez����Jf���V">�J�xPŕ�k�x��5�����Y�Վ	�v"�sβzMGD6ւE,�j���2�B`ؼ�#���(hj�����1��Y�m���%1���l	Nq���s���K;���3���g�i�,��!�Gu����E�u�Ȩ�͌N88dd4�T��Cv�ʸ�H2#)�=qp�C���0+�c)�p͛Gթm$�jR�",|UŌ�Ř�睐�[1����7f��5ǝs�>Y|�Sˠ�ZC,���Q��Ɏ�xT�U�|s"( �5!�:�LB˖��j���l�V#X� �9-�ݾ�
6�8/ ��s8�!��mծ�s��֕�N�fӺ����U�k7�(���Sߡ�����n�9k1, ����3 �ˆ�߄c}H	���Md��58�I|�����xW�R݃5���_\}3�yێMx���2�XDF9�Di���\�:�ƦY��Piw�$Dh�a_�H_O��i�)�׀fĐ��#�F�fY�!����{��hG�AC	)W5D-���=|#1�Uo��8]�@�ų��EH���,^^�5N��4-�?��{���t[`n�XV�k���u����	\F5��4>�~$�orM��@gl����\�H��je���P5J��b�Ϲ��J��!��I�D�v � 8*�����^,%�
�װQ�D���&6�	n����r"��l+�t�]���Sfct���~��ŘݻL�:SBh����������! � ���\����_���;I�7��4i�]�߮aeE�Z��F�<P�^�a��P�c�2���h�o-�wH�����ѝ�������]�ҷ,ciΰU��t���%J�?@WLXe�m��{��q����H��,�E��PkC��/{A�bh�l�g�_��&1���K��I��K��5��w�xG4�Q����(�K��`5��=L����緒�#Ȩ���ڤ���߰�0��ݮI���~Y)��.*~
X���"����!�'����%��d �uL�%��W
��pI[:l&vN�Ƚ�m'7�L����G|�/@��m�g Ӑ�@��L?�R./����;?m�.�r�4�%�ٷ��!Qk0&Mс�x��b�~����*�<i��Z�r���V��2i�	y]�#�k1�k�O�8��&�������+[׵�ԭ���@ y�y.~�Zz��ã$��۪�K0Y�s$�i-��d6n���M���1r~8�6�<7�*
������Kl̊�:�?���#�n�L�-�ۗ�e����Ρ�\��tl;�����MȬf����ޢ*o]���j���ui� z�)⋌$���1��T��J�[����9w��<��;<����ڗͻ!ls�Zo����ՋmnX�sb'��y���lB��;+�2QJ�����s}�6���Җ���Wuq��"��:�����Yf/�%|(�� %=��Ӟ=�ĂvLɸ�=w��@+�e3��D�R��Zږ�'_܈M���OӃd��]tə=���qh�̈)�F��d<;��})��"WϞ��n �s����Ρ���	`�H5U�!q�{W�p��L�F'Coe���b#�2���Í_,$\�Jؘ'\ؔ�P6͓V׺lĈ�J�ѽ�.2�ɽ�`>�0�u�g0 �;8ru���t��
�H�.U��3�J��W���"����[*,9�gFq>(ք'������}Wn��sfSn�P�??`��%�ֲ��6]��A[�-w�3� �� �6m��u�Q�{�S�j�-[m�j9hNt ���CMrC~6t�$b|�X�1<���<�o�8�C�C�"�zڟ(-������wF�:�)�{bx�1e\�,]+�� �!߮���a�zۄk2Ė�C� 2a�#	C����'���uO��"`�L��?�	ۃ >D@L4���@���(��G�95���t5p�������@�J�n�r��ײO�Q_uk�+�(F��{L��oX��� gNcE�+�c��&�I�@��T�=r�9%Ɉ����)��GY�$V$�%�d����0F�u�����
2�o���;�z�����K�)@ˤ�#K�g.��9�1J	�J��;Q�O� 62x/jK����������2��8\3��,o�Z#B(���.�֙�-�q9�^w-5�h�25M�]�E�D9��(����9�P��6�0e$u:&o����Ô��*��������9>������<<�ZDUH�Ҟ��� ��!�B�M�mPB�����dX��&U/K�7�g$���� �Z�?$AF݊�qh�v*'�A~�G���}b�e�]�e�	�6/]d���-�|���<���aF����i�~^����a��-�	�<��:B�P��1�v2�i#��N��������z@��u�N/N��z���`vH)�ZҴU�+��8e6�*�lč5����A��P��p��g2��	�α%��%�(���
P�0�V6�*]8��Z�vW��^Z���c= �\ms<P,ѼU����_���(a�:�6���I�hB_)��4&`�"��R�����n�?��pqc���Ȟ�&%|�Y����u�f͞��.�Y�M)�Y߄�V7̑X��Јe��^�e�j�8M��F�2]�1�kk��兩���%)=��Z�6G"�r̉+�U��MuQ��%�SmZ�3r�}. 4�/o�ŸH��U9��Ĉ�&	���/��"�����7_��C�f��ʳ���I��r�؉@_6�c{�͋H��Rq�4u����e��2<��yf=!rL���R12��A�7m��7��y�)����(r�^���������[�z��J��qh]��\�����J/�L�:/�Wvs��4�u��e�E�u
\��(g�A�A�[a2��5la���פ��h�?v�梳�2����I��f�>ݺ�^��d��{�g�V�<�^�U���NZ���\�H�|^YB��̏��?ΐ�"zO�*��F�r��x�e�$Qv,>���aIGU���ײ'xs���b������9�u��X>�Z���o���5_싶f�����R�`��ӶTH�͠� ���A�/�M�|�!�'u���9jɩ_����c!�Jͺ �6��.^=� �]�-�׎�Y����X{�.�WB�X_�-G_�uqic������	��ʛ˃큃]��
U�bp���5���7�+���ղ�=a�o�����>(��#�e(�'�@:r�`ȟ?�[�9���a`Dt1���n�=��F��7�f�ˋr;p�[��Rū�E��'f(ee9;և�ʛz~�h��Bp��٫r��p$ݨ$H�ߩB����O�iT=٧����
�"�~�`F#�\N���_R���&A�Q����V�Z�;]fW���,����&!��Kԁ��"��mI�P�\��3vOg��'�|h4fq�&z��>���.�_��fe�̍P�<���7QR�fF	zε�+8�oo!
��LY�2���郢��r\I���X��Ժ-P[ȓ� ���o�k.-��k�μ�,���]�c�����OFW�7�X{@�n��;�}z'����2�X�G-u^!�fRAL���2���>�Qi_�T������-�v"'N.;s�Q��!�<�P���S�vt�o�)�Nx�I9.���W:;b�i�&���`�k ek���Z%�!d�8\u��ȳ������3�?�-+���Z��E6j�D�^�Du��~�Ɯ�����4�p&���c{3�sZe�PgD�
��(�;�;p͂�5tٹ�Em�f��ݺ!D_H�']7�#�7���䰘T_[�-�+q����k4|:z�n���k�S]��LPq����W�����Q�f_���x�~�* Rښ��w�_�r7Z�쇑��M����~�1�Û-G����g?�=%�w����4�$$ݨ��rP]�?:�ݪk�9%a�ؕ0��o9��L��٣Q~�,��U���k|4GA���a�����?�5���IwwZ܉,�͈avq�����3c䊚�����Ϊ�v�v���ʣn+H�8[�7vp&t�x24qp�#��T�a�vR���.�&����T���?�����d��w�@��d�P�E�'r%�{ �59���H�T��/Q!�ȍ�-:��7ؒ�/c�ﷳ���|�� �O�}�R=Q)<e���1����iPP�C|�5p+ڹI�uvM�6`Z	��k��Y��n����6FO�H�"]#�z����L�*�}�F���d8+/��z�܈_�2<ݪ�Ә���B񌎩�:C`��?�Z��\.�u0^�׬$d�It�v�e�$t���0����r�@DiU�W���R�rZ�u��E��|�;K�<9�:f�<�Hx��~Щ;+LZ�����*(�oO���2�F{f����Ƞ��\�A׼�s�^<$��>�vq�= ��������&8�T����css��T��9�/'�|�Y3[U,[����ސe},��9�3����� �f���I���L-@�^���T� ���_�4��pnszڤ���K78�a��O���k�7��J/	~!��ue����خL�����H��+��	�E23Z�Y�*d �#����Ό�aBi�v�*E��l���zD��Q���?�O%�^ Y�"u�"i�P������at.���-�_�h�8������F6(~w
bH�ݸ�<�A`��j�7���Ct�A/5����*���sϐ���=�Vx�������(03
-�xI̴Q��d�w)*P�R,c��T���{������V'����:�]�J ��b�;F-Q�����2H=��%�"-�-��v��P���+�y1����㬣�gl��+�>� <� �ܑ) SG�RW5��h�o�	��<U�"���2���_.�B�E�&�����LFԅg\e% 8"�	|�q\��S&3�2�sD��w��i�ؠ��G\��Z]f��Sn!���;�xn��KAl���ﵼ�A���y1��I�}u5s��F����� O��^3J,.�G����!S�҂q��;���u_C&��M	t���~����?�T����`�c�?⌒�"b�@�«��q����6���e�I��v��U�~е��>���ǈmTz��UvD�}�>����uBq:a��C�-�M5�g�)��5�*��r�fg�,캫�Z-5o4�P�|e�b����X_��Y�V����=߾:�/cX��G�H�`�	ֈ&�����(7�`z�,��+��ÊL&�W^1���MH%�$<�WBA��@ &UZ�+-�	����a#��NEA���A��95e��Y� �z���!ʻ�,��/���͸�D��`�@}������ �>�B�9`���N4�����U�J�����o��_��Уg�M$�������ޔ�"N�� ����؎�f���q1@
����q��{=N��j߼Y?Ȣ.����J.�������L��7��rL���z�Q,t
�F���»���姏1_��� C[ʑU3@��Y�k%�����VG��²��ޑQkF��c?Q���A����%�&TѾE�\TM(��z�bV�
��YqQTQQJ���!$.L�NOʕ��)G�J�<�"��*��>�S j�������c4�:�FZ�;�c�M�5�5���_r=�j�����S��3�(K5�y��y�+�=�{~��_Pj?R����є1��|,����8�|��P-�L�J�/�}b*�W����$Ƥ,u�x��m����@�c��<(Ɩ���C��Y>������G�ѿ�d3֚4�x��6������9�I��՟�!�������}f�!r��AT���-$��V뭸�DT��$����"F#�9�׵+�g��߁�O���ȒKA��R�#���r�������J����d����(ɻv�At�)�5����5�Zr=	�ԓ�!Z�QП��G�H:�Y�/�Cx���u�����	��~����_He�	|��^A�y%n�����`� �
��>�f�2uw�+Wd4]��OS��Gf���4�{<W�qJ��@lNRW<[�ra�BϞp��t�Vi؆S<bx��#����ӹ��v���u�m�G�����V(�������Fb܌�T�ݲ�{4E����w8�����K�&�.��K$0�×���Jp�$:��/�u�z���~Q���@�����#�wTr=����/�	��(�x��Z�.iO�q�YxA�!�����`ޤ4(�T����¥ ��J��y��Y�S�H���@]�{�L;uS;��W�~�R#X���o|��K���oёx�.�B*�Y/1��Q�
4c�����y���h��uCǤ���ώ?�C�(�'�U��om}M�N <�\��r������S�/n�*=��ݖc P�|�[ИK�d:�f�D2������{�Gߣ�7tͻ�$��[�E0F��`���7�6�)֟ꪺ�
j_4_C����}H�b��[4O+M�����\�:>n)~>юO�RQzE��c�BS���|���0��/M�Ԧ{N��x�M�ڀ|2�K�y��輛	��h�O)m�Hx�׃I����{Nf����)�aa"xjg��R���Ix����	��Q�9[ea����s@�^�7F1b�ē�{C5>������I���켖y듋�2��˦	�	9ݻ]��ʞ��.-k���_WN�2l ����+���8��,G��Y��<�s"�U@�=��=��8/�˱Ƥ~��ץ�u@�D����xy�0D�.c{例�0Sc4K�h[%9-"��	�"�O[�="^L����֠G�]@����q�U�f
��$�B�O��B>]��U��ߘ&��U� `�r運n��;(ҫ��!Pq�ğ�F#�ުk�3��~@�$�����NI�+�[w�A.8ś�<��҃k�c*%'麓��|<*�Qj'����c��3�%��E���*��{&\��'����I�=VVn�����a�8�S���Tģ���w&GR7�M|�0�'3�t��b>��()
����VSE�1߉�˖���/�΋Pj)��˂LXk��r+o�{E.�g�=�`�Tr!�����lq���\�/y+C��K��-ذ+�)b��������d�R��M;R�ž�W5�e�a^��:jq]ps��wO�R'�,ǍX�Š����n�*���AS��b_��~p]s�߅�3Es�P�q�%�x����@;;�C������]a�cL�����ρ��҆��iNpj�ړ�uI*��������ɦ�׶��2�o(�`\��r"q+��;!��-�&��jϴ)�?����-���S"D�K��hTc��?��x!��0�Ш.�z�\�&,'�A S#�m1��Ix+�����
�OS��>bv#�`n�5˓D�����,�mب�~�% W���������hV� �PW�� ������$���b�L�Q�)��)- ��?E�pn���XB69��b��.�u�㗿�}�=��������#e��/*�������s���T�%�7�N�ӛw��y���a�G7៊��� �%UMn|?���ؓ�_D�q���N�Y"���=F�7�Ԏ)ޓ�G�Z�+1��uVj�>"x 
<^��p���������ʩZ�������Gʮ���ͮ�`���/R��[$�E�Pz�5t�Q����gm�s�Qݞ9�'WJbo^�E��A/���\t,���,�j�^2;��@���XNɒ ���$���*���6�r͇���}S�6J��~܇�i�����T/�c��[�����6�mz�U�J!�fy�i�- u�ڏ�M�q���WN�!D�G��<���C��� ����Bd�C���'�F�\�yH%E�d�,���L�$�����5a�c��i!g~?`��~�ȸ�'B[�<g���<j7�� tY�`���O�4�n��E��,J���}� 8��ܯ��D{�Σj!l�br�9P�
˜ǾP%����U�S��� �Sɵ�h���K/4C�@�_lL#BN�b?G�n<M�
Y�O�ʃ�\�?!�$��Q(�%;(����$^K��F@ń`3o`��xR�-��21���i��pm/�`*u�b�_(g�F�e�M&���;P��ID�B#1�q���tz�HU��{�E>�i��}2[w�d�#��q���Q��7��R73����j���~y1��rѝ��H��c�P,aW����<��_+�L�|<Uz�%-M<��i���]�p���F�Ŭ�L$�uv�>^7��j������FO�❲#u��b$���r���Hݜ�_A
�P��)[>��ëHmo��k�������@�f Ys*���8+:�r5w~�Wy ���&�Y�քIb��w$�����
�e O�wOt���QOn�[F5�h>|I��Mj�DԶ�k�K8��Q5W@�dD�¢$��A�9������NG����i�	!!/��'�+�&��7�Y���Ej�V�'�ī����Y�	��A$��)##���"�fkEa��o�I�E������4��rC�vujC���`T�'�	�%fu~) �7�}H]4���*���>U8���ɘ�/\��2�����d~�7�E4 � �p���hļj\�	R�=?֒�"�h]9V0-�̐H�;�	å��B�X��G�b��;��ǂ/ya'}Y��l���FN����!��ӀẂ�QG=��+��z�����U��6��x� �|
��΃P��j�Y�$��C}v�Z��=�bo��ל��=eZٻ�O��h���E#9�I��b�	uڶ�S����Fm��]i���=a�*�?cvZ�t�.�قwL���1&Ŕ����&�Ww�W�l�PjO�����YKDU�2���?��"	�~����t��+z4�ٟ��1�R�"�QN�dSW�4�A����4�k�[�`�!� �O����1���gp��Ҫe+w���Bh�)����'	����ᩆ�-��M�67����U�(!��E7�鵋�3{�2%����$��p�sM��(�-���j�A�i�+�m��=:����7���H�G��~i��W�qް���t�J��GvI1a�{�x�B���$����վaὍ9��.�l�O�{]�ؒh����!d�Oٳm��˩�0j�W��z^�Ou�!�(�_��;�< ��� X���UY���u[��8W՗��7r8;qʁw����$�e�o�F�ϱq03�=/�6���닧4�����f��Gޮ��r�^ۀ�@zbv�{�F��`lK��R���ٛ����V��G�����X������2�^lAR���f>��7�����*����T>�?��)�v�1��Ӷ���2+_�B3^���^�a��-i�����U�8Hf�����d�mH��Ϸl�gު2�n;7��[�\|D�ʪ%J�+2��c�yvf�*��"|yX����\�a{�hu�s��9��߰�¤�L��/D��b��ң�����ft�k���p#:ָ�o0�#L.�3=����c��8V��'�&�V[N͊l(���	ы���sN �宺����U{��7?A��w���7�xz�	`�r�&�i��O���Qj*>dC.�6ߩ������>Մ����Y�&HNa�1��r�N�X�f��jT�"���Ax;�5@�fp6՞ޱ�J�ʮ}_GG�o��=�C�O�4m~v���jB��Yi����%u����}�ܡs'_qUV��l�R܅5���̻���7,�f{D%Y>P|�M���k7�F��P	�G����"��?D�I�~/���Z�a񙟸��z��G*�3T`Iޙ5BW7��W�K���Ǥ7�)8��UH^��<�0R��YK{���`7l�8F��'8���A|��;HW�Gg$$DƛY���IM�ʢC/�yo1Qh�P�]�Uϐ���d�]o�M�`����\�� ����PDڴq����b�y	��8]YB,H���<��G��������R�"B�*W����!���>Vf
��,:N�H�nto���i&�CQ!�YS�����4�g�4L|��pGX֮��!�w�xo��*��e��)\A%���/;���s�j(19䃲�Z����XB"��+�(%r��[Ү��Æ�&!��//|&��@J��T�8��˨i�Y=��6Ã�:m��JZ�L������#�^P��C�\ ���(��wt���3�\J��W�u�(2������[�-�� mF٧&��ʻb}B�d�'U�C���p��U��Ť@�z˒ 	 n"��n������?b�������˧�����&�CI�=����b?�R���kn�Խu����4
�@X��1����������[�>���p��[4��E9������ѣ��S���q�X�%�P��y��?���v���a��\)^��ը�X���"N\/O� Q��cXM�D�mN�Ћz���k���'�lw���ppQ1L㞰�u�X9���D���ɕ�+q&�Be���h�?Uo���y�ܞ�ᄬ�� �)ن��np��Y��ˎtî&6L *���h�;�1��uלHrG8��������Ãe@.i�k���y��la���<??���ڀ-���PbH#(1��k=�,�k;���Dc_�7���)������_G��U-<���gU�tX���ʉH�Kk�69X��d�YTͫ>�� ��M�7�ty���II�'��v��� Uq¯l]�<��(x�+�ՂH(gN�Z�,��wb@��
�ާ�.�m��m'%FNg(K��9���1��J��LЋ�wŴn�=�'��G�ZD�=ort�첤=����i]tOcD����Ծ�]��T��z��0��vMA"R�$j��Υ�v��BO�T�PhN���7I#G0�Z��uB5v��6��tj�� ����������� Vl�i0����0��ڨ��1��%Ż/1]_��(O����8�h����s":���@G�.�P���� �&�li{> t��g�<	���$����[fYo>��l3��t�����x�U}�IS�����uej��OM�v��밬2G����j3�����FY��0�����^�:�j�P(�#��!_/y�p�_��ܝ�!5W/.4��$�f�$'}�:��4�a~�HQ"����T� ����|a�gr���u`մ�Y|�~�<a~����}b�#�F[J�IXj���4/UʅѦ��f����/.4��,�F�_�F��Üۢ�<�������l���W��,+�E��2(*2E�l�^oV����y����\��_���AEA����4�5P3j]I$y7Q���6�@s�Ն�,����oҌ�_4q`�V�%�����_HT�#r�nE��z�A�r���xC�+�v���3^V}�**�-������%��x��$�Z�N�ǩqK�V9��U���r�%8ٶ�f$V2����!,�m(��g��?�a>L�	3��<�f0I�u:xg��V�u�@s�B�f�]$�vYL�D��O���G�vb�fDt!"�ߡmJ����?�� �5�김�� ��.2�)�Ȟ*�_�������&L��F��ݮV���{ :"�]�O�����z�^Y�֦�
����G���yƻώj~��B�n��soV�}\XC�\�/!$ٍ-@��P����.��!��w�tT����E��C�L�JZ�ba��/n�v�q\k��e�2�a�Q?�4.V��X`�j@dQ:�ѯ�j;b�_��r�]F����͞�rx��3s �uŲ"���q;;j����z�8%O��)D��@���\�/�Ii�6���wn��(˘�L�&n��+���+.M�X�4`Ôfo���h�<�=��|�L�������/�F�	���ci���T|T�"��`bt�V9vC���v=�g$��EZ�U�6�Jh��?9={iIe��a�o�^����ʠ�����<:��(k'1�ǍL:�|����X	"ln���C�3�b�\j�:%4)�x�P�r���U,�^'��S�����dG(��G�$Fb������jSA�Vu~�#�p�f�KJq�O�[�s�ζo�G��Q���!wXg�!--������;K�3�T>�%�ޫ�:���]&ՖT�Q�><�5��cG�����s"P��k˨,W�����pʑG#|\r��3hp�.F}�Ҹ�]��o쯓����t�:'�ڶ����3;�s�F?!����fzr��]� +uc�J�C@Y��)�㣐}�nzT�!���Ɠ�4m����aw!ܬX|g1 0�jO����L�;9�1�b�i!ޔ�D�os"���J��(-�T�q1��\�Cީw���3�jG��v�x�wÓ@�O(>$�&�N�3rx�E�ރM���\�$��i�Yv����#G�[VD��CS�Y'|���T[G���	�}���d	�WPD�=����G���z�{���f�i�_}�����d�q ���/@$���
�N�o?�X:��45��SߌA�t�נU�q0���Q��K�Q��gSy�o� ��>��E̎���EV��>3��`���L<$�D�լ�G����D�S���j���70;9Ѷ��3f��G>�5����K�?DR�4�56k�WN�ڣ�|%��k��on��}�	��{⭁L[X^��2�S�J��h([7@R�4�AT�r�`̥�PQ���TWfs][4�-��L\/>��:V?n��� �Ă����Q�&�-�5�G�`xS����0��.g[�d�r��͡⼘Ǟ+,%��\m�[O�����8�dlM��ME��s3J@<D�}Z�6�$GNv<�<�}�/��w�� �RG�.򡬏b2�_�rJ�?� i�p ��p�J\fv4��u�`j� �D�']�M�R{r�S�7x^�ン�V��h�M���
�D��C�g�2��y�O��F������g~��n�s5��2�"��J�g�ʴ'��2��Ğ�Qh��쑂~��X�?� O����Ǡ-!J�a���!��^��W!��`���7�C˧��S̎�~�Cf�JP�wbTaC҇��8����֥��<3J�����A�^���A�TL�x`ŏ�{�n$D��o�9��P�y$yNa��螴�	:�4@	����Pk��l�Z:�L�(o#)���O�2���)�?|�M(�����g���-�?A�O�����o�5��%�%�Jf?��Ӏ���@ܗ�:��1�,aO��t��$j�>��u(��TOZ]7X�g�|����$����-Q��5=S|�ړe�t�ȦÿR6'b{֬\]��'b";b���G�k�e��Q]�������[�~5�S�h@ٚ#�B��H����E��G�hR|z�n2B�-ńS�����dh���Є�*�����?\9wr��ت��MV!�*,^:�>\�Z��S����S�n� ��y.����ɁG�!2�D��ܡd���1���<W�w��}t-�n���X~	8�Ғ���3�r����З�Ⱥ�x�6����k�$1~�x���^�{P��>5�'`�?��T��Á���L0oN^߆W�=�p	�n!-�}��f�Q��kL}���C�l��f+YΆ������8L4V��U������Ih�/�Zern:2�~���$�bBvO�^�z���_'�n��:���w�|V�U���z��n70W�qΚǫ��=���Zтt`U;�.x�[��iy�� �8�=jz%|����@^|���*ӑ�0��>��>V1:�>���Je��1�8c6�<��hed�TH�za���0bl��Ͼ���o4t�XL��g쪞���]�h}ٜ!���t�����eX>��D��j���Y`�N2L���܋&0�d��22(����#T�K�i	Н_B�e��� ��)E�p̅�Pg� k�5N��Z�92�ì�/@3���<&����[���Sz�1�6q o�㔫����Y$���ՐS���u����a���/*��̬/^v�`���rwI�����l���
Ѻ���۵jd�W=�o������-�)�� �N�c��_s#�Mzٞ��Y��E�&�N$'~q����{X�YN��s����(��F��7����>q��_���\�Z����_�nX*ȗ��,�3��n�e,�x4,ǤC�� ��{M�w�U�-1�V��:�)���x(K��R���ӐC̀���9�0�v�-)H/���V*^��1�$3d����7AW�k�pD�
U"uC�d��V	u�@O����l��^�{=oS �xv����b+�G^��Ɔڞ�i�N?+�:��S4�u�NS�w�f��0W�^Gd�� r�!���0�yu������㾒���N������� ��h(s?���O�5>�ӝi���e�y���	��Uy�~�6�ÿ[U3�X���$#�b����~LB,�pɽu���4��خȄ�`w�Wٻl�ٵhN�q�*�Y�|���,��:�*d�v��f]���O�F�qV�)i'�z��'�3u��u�7P�p�T�Y2��0�
NL��
�4�l�*�o`�����s$].��ܢ��#^��7�-���D�����a�n9�M�!���jm,w����v�.=�����5��l��z'ӓ��7�phP�}�j�'���,�rJ��z�g�Ǌ@�,=�鵆��Ld �:/��ݺ���"VPx=J%���ǳ��	��{O\�8��<�������E[2���`	 �>�<s�4�q.�;��_�p^i����D�J�\���)/��.���F��N�� �?��%m|���
)*��N�3G��I�|�?���RD��ԋ��`��-�˓L7��P��~u~�u��3�H&�R̰r�{/EX�%(K���b�q�w�K�a<�~�����N�_��������h3��_�L'�&����k3$-y�*�ˆ�'���C< �G����DZ����b�ڻ�H]!�{o�K�Q�ܩ����P8�����s�J"��������R�6	��,�~c��,�a/��V�s��l�Z��8��4�T�f��W-��{.�{}C�7\��g}ty�l�,��o��! E�/�I�dt�Ʒ<Ƅ͝�98=Z"^E�K�������[�{鑘e�f��w������RcZ����ӦW#�����F�����s�i��Gbݪ�䟤<��^�6rJ��ZT���3V-B�V��nH4숵y�ïCiNƙ���ہ�9\j[7���?��y,1�Y�"J��|D��>�Vm��
����R*Њ_��Gw���ɣ� �Sx|��n�O���\�e��DGd���g���HOhw�$A���M��l.G��H"|�/�������0�?4ˏq�A��xC�UJ�	�^�_�b��ƌP�rQ��/���N���:�ALr5�+�`���(=m2��(��B���7fS����.k�:M��N�MӜ��z���<+���{�b��-��K��ū�W:\:�l���L�xMӖm�k�ʤ�#;_U4��s�Йi�߱$�U�$�៮�#�"l��M��}v�r�_,te��J�ꘜ�GJ�rB�;�l
�SS(`mf�� ��������P�Ժ>�0~�Jm[��
^�9�1��a�_�8�<Q��EJ�����
)������2�e3��K��!n�|�}��Z�ZYu ����mKP��̳jA�y���Dۨ��2����&i���yl�=�s*/��G(������1L��0�"���Ǆڕ��hԡ���`��[*��R�#�B��B7���_�Ԑx�|�=��`��Ü�`�G���q2�=��]���j�/���\�e�}��ק�zy��)�7�]��>��P6d��(#��6�~��u$mI2�?*O�����E�h��S�i�yŰ�S-���Y�Ɣ���?��4�2��e\$Aӌ�gvI�j�ɆQ^ξ?�u5^{S��n@� �Q�V��@W@��#��t��c�xK���G*�O�Ue��'ߡ~?���wE��i��i�%�b��OT�k=�yT�8N��$ �t���I�>�N�oUg�t~�=������Qc����d�V��D#y��	$뙐}}$)(o��j����+"�ԊKo��l���ji�xB�r������p�`����"b�(�a�hX)�C�e�����c��^����{Z `)&�Ų)���6�E�s��b[�V���T:T\��n����(Å��폮�F��2S�`���){��鷀�!�B$Q{-<��t�?l�zax��A�l�OOMp�B�r���]�@�Ә�$��X�n�B̟��P�k����JD��$�O �0�<J����.��MQ.b��Q�𴣨�5"u�W���_ qɼAL>g�R��X4X��Z+,Hǁ��Q�F2��r ���Fi�Բ;]꿤�����R�b(�LnS�0A���M3rֱ�S1m�3�D�@��]�肙)��\"
����:�2*��\�\�O�08��ü�ۈ��?��&j)pƺ��q���~_>N��t�8��77Q�AJ+�im��ڪ�y�*Wm��1�X|Q�#�Tx�k���1�0qz{�����)"6�~.�N��uZ��#�vb=� 3`Q��!� ���o^L�ӄ�l���.�a`�=��hV�7�,"3'&�_��5��_N��cF��v2NySP���#'����ҰL�$�'`Lދ�N�x\X�>��<B��~��k7��N�E���1�aNa{���
8Ι���pB�31�j9����x�y�a��L\�4�L@�'�3>�BSB:X!Ґ�"�4s���o�K0���&s�$T���7����e5�{&L�z�`;��y!��6��Yfoܴ\k �w�"�e�F���};�����\��qe�N�%��8��ò�6h�'��'�^aG�i�� ~��S$���H<l�6�ty��-pW�\0�ә����j�g���K��ʩ���[�v3	�ar����c���	 b}T�wrhD�%J#/Ϯ���B
����gpLS`K�L�}4[B�!�6��bg��{����P��;�����x'��_/��EpL,�֭�`�9�|���&�oE�[�nZ�XG����4��k�'�OLЩ��b\� x 5@{7���tU���&��׿z����BOb-�Qh ζs �w��(@�yR��}���{�Na���yӆ��4��' #�Do���Qط�}E+�)�H�E)�;��ĥq��༕�t�h�G��h->f{���;R�����{.z��w�V�� V[��0�c�(1 ��{�j�XB��v`0�(f�A/�vzٍ:�xr��@�O04A�>�y��^�a(���RaI����/�=xӸ4�_���([`�s�w��4�1
t�y�l�M�6���+?G��,��xշb��,��=�s$��YQ��S���a呋ҋ\�W�$�눟�q�7�o/�˪��e7%���� *����Aѧ$~���@M��A�~;Е��K��5{C⸄v5j=so3R��,�K4������;4~*��[����H��C�f?���WSpMT�/V�}�P�T*���$=�w@���U�<T��8��봌2�<��ȴyS=�Ke��ˤ�Z?Ϙ4IJ
*v@r��8k�!5�%���ݶɣh�)@Q�I,�g?�4N4(�II/{��wR�cQ$ I|����Z�9�CJ�ȴq�iXQ�9��@EW�g%dP�W�M�:x�ZlلJ �\--��#�]���2 �4t1����A�2\���?��'i�8�h��2��8����W&8	Ev�nL�6OC� �0�lT�}|8�X��W^x�G]2�4�%�y���D�L��"�����a����g;�P}�`|T۞hw�}¡$-� e��wb���@� Q�!R��D�ΰڊ�ʔ͐tM�X�}������UeA-7�V�T��QNTZ�:АG결�����_zcit���~�t�5���#���qjX8e���t�"o(W8�%%0�v`-''�#�2��\�lg�������z�n�t�$�jBa��W�(ӷ��(�g�{&�\(&���34�d����$%tY���k.�����,6�?�	�M��T7~.�a�S���Zʤ �Qc|��R��y���= �"�� �ÌTT粮�� �l?�b�djo-R���n����w��AAڜ$BG|�)�Y�v�Q��Z�h[�v^�+Ia���u��C�$���ٍ����|1	�J��'Y���x�#]�2��ܽ,�{k5�"���0��rz���P�b���o���M���h\K�O��3dX����/N|�iX�/��H��q�hqm�oj��P���^�LL 4�3�F{�PUMt_�E�ʷ��f�_�³��F=`k��
fx�����L���q�?����2�=���c���{���ey���De��!�����U�Q3'�%� ��˕�%����6o��n����_�#j�,�"i�7�WX�3.�E�å@)!�NH�,!�p�����-���Ҿ��:'ҐrF����*�˴'�|��z��AkIE��h	WF$�<؃���Z�M��_��=�_���<�/Bp�<����r�%Φo��La�����Ş5�_FՋ��KòM�����d��bӸf���{�ٛV
�&��sBo���T)��z�k��.�s串����`x
��e��N'�?���n�&w��p"P�ʞA!0GU A@s�]�8Qz�S��?�$���b3`�0�c��i]�h{��3��5t%���9{�X�	D��ƨ�X�a�rNT|�<�,#n�O�����t��l�9uW�� �.��*\:	vNy��mPЪT�����bU���S[O���W��H#J���*�Z�.�' 	g]�/ rQJCD�_�	��o:�7�%�Y��3V���G�:��F��60Fq3��*~.G���`Rf0����Ph�X�)�����'����#�� ��'��I�d�Х1}R�=$m1�x8��H'�z��#�^�Q��Dg�Z�" 2�0�ie�MO*��UK'�6	���0VO��G�� ^}�I(�fw����F;��Ӈ���j*�3E�(��>3��Z;v�LD��&^Q}��X<p���s�pI��&)����3LG���]=�A�~,d4朌���Ά�
���kP�YV���Pj'M8�B��ֱ�?�ꮜ��*5�d���C�"|Xn�%j�:��Ɣ���C��!f�}�b	����%��v?��'ݭ<��\�����7C��Q���LfHo��v�ɲ�4�Ώ7R!0fh�$����b!��k�J��b*J�ɘ�Nn��F.��0�ԮY��Y�K��\����v���H5q�x�L4�C�44T��9��Sq�o�B*"%�d����醼ݙ~�B����un�BpO���?�w��i�3	�4YI"�6�ޖ}������y�n��S�-��枊n�1�Q���=��$�����fȓz�1����)$����S����`�c��J����׋�h��4&�����i�?���! �=� g����Aʾtd�w⋶r?�yK��:�E�1���Wu��Cj{��\8]ĝӈ	�alq,�ZQ���
��|�U�2�����*�I����]�ٔekL�N�Uy�
~�t�-�Fތ}�d�䈊C�ؘ�S@ #����緶���.�����:�8iČ�	"1
��%�ϯ&����YPS�F�qs5Z��5T�x������>!��>ֶ��xy�Q��$|��}�"�0`��,^���dd��"�+�S�O+}�����*�v㗱�c,�dhY�4�O�j�Oſ��~Ǘ�����]ӡ�I���Q���{1�MB5I9:$l���X�j;���ҽ� (�KE)D�L���L���g���ξ�]ľ�Y��	�:|��nmӬ�H�����@Y��ʞ,G���H�`�&DH|Ҏ��/���V����R����<�*~�fm |c�7O��&Л�A�΄/�N
uR�;�qփ�ب���Ѝ�6������N�����n���aj��У ��� �{��	��Fk<>��a�,�?��2��<Uc���ш��j��l�G��N뽊��w�.��_��=�X��}�(+�~�z5cN��0��_X����k�.%�e����.�����Z%�B�pyќ�q,�����*���UVm��v�ڵ���W\���C��B����N�L.���R�+�=�E,Z}�U��"��Z�#-z+�N8}��P�{�+� ԧ>qH;!�Bt��]"�w��vY�v���mNn�#�s�p�������>����u�d�� ������R��.�kFBI�$B�AsM#l�,��%\Cn�:�.�G<S啲 cIV���qLb��}|}�\H��P��prb�4�5�m#���_�1�H�c��Ƒ/s*3�uZ��0�P��x��������S�eƴ�V|�����v��(i�~ѭ얢�z����hp�\��7`���ݐ!��TM��@u���I�Ъݰ�$H
�-h�=j�7g=�w!�c��;�-ߚ>��`��%�F�s9(��=4�3�ܡ}4t`�����j 
�ݔ����������!򻖥��]?k�.r<�k�l0�2���&��#��W�+���?v^`��@6�HC���9[˭��-���!H�5G���L���mؤ+jݶ�(?���ܚ�� ;��6ǞΤ���"�B���,�&�"�V��M��=�h�HIC�V��OM��uȶkVv��XS����(~���|,w����|��A�.n�X��Y�����q$���A!Y֩�t�q0�z\���A� 2�ҹ�G�L����!$m��ՙY�d:�c����hI��hq���Y�3�}hnB`��S�e�*��90�)�1!�5���������B<�N�!Dn�s\�$r�� �*�.(����'�צ��#�k@�� KT]W;,.��-���#0��K�a�+l��].Ѫ#0��(MI�М��������ĢGVlS�7��[B`��Nѐ*�t�jpS��rR~܃��D�]%�����$���}j�q��)���Ii��g��6��w~�B$���pA�N瑵@89\՞|���]�d���������hnK~Blm�3���	O���w)E���yP��O�����o�/8�4;�ZN?���.��;\p+"��a!�Cb1��ǚ�ϴ���8ɟ�����A�t�ҽ�I�\�#�Rծ�A�@Kj�걑U��P�1+���V҇�`��gu��\K���!0h�R�lG-o=�n�-�)��>���c�b{�>Q��8ȟm�JK;.���>�<{������ךtv�|7���x�
�a 2��kE��ہ��d������x�2�4��[��Ís���V���TQx3°a:��<�^�`����xݧ��Q��a��Iص"Z�^Ғ��9��݌�m͈��?�Q�Fe�^4>�p<`�M��5����9'�h��5�'��]Ml7ZS/�H1�ڎwT��a���y���yr�B0�b8����ɫ���T�0a�+�Q����q�a�.�o֐�⏖����1�t����r9Rq�"
�x������O��7�e<-=J�ģ��m���h����Ś:�x��v�k0+����*ҟVA� �`yY�B`�W`�Rk4ƹ�\����Z%�	�����-����d�bK����R�χ��r�}�8���Q���w�H7���q���u:��n���m���G��n0����_b^R���H�1V��
%}4���~����ˁ�����'W��#Ip@q�Q�q�\�'6���٫�e�9׶9u�����Y'&RM
c~�y���H:e�X���8ij6����r�g���\p�Z�.�p4e�� 8�&1�;�TyR��lIѸ�������R�H�QX�}�Kd+ȥ1.�88��c�I��@n���}�k�+	�����b�����%K��Օ��y��ۍ����e��6�(R`D_�(n�j��%\�
}`PsU�I����.�sp�H��&H�?(�F=N���*J�i�C(�(���J�0RO�=�p	@<�S��̿�W�1��;���q��3E�(��
TX6��X��PiAyc�è(��o[V{��v�B7�Q�v�A_�ɲ3S�cf��'��Ā���󆍈t���B��
�����As.71xnҭ��֋z�#%x0�Zs>_����t�67Vim�D��.�7i%³� �*��������a�I����<�?m������Lo�KW�W�ک7��M}.�I�kk ����Z�q�?~}�V{\Tݐ�דvbH�XS�x��U!�w^�#�yg�.~���dX���@����=����/�1�z�߀��ֻ�����g���j�u���
T�3Rn6��?$=�L8N�3+ѱ�h�$ϵL�DB��[���0{�yH*yb��pM`P) ��L��޺4��B�7Uޑ��(ڣ�6������y��&���e�d_I�w�Cle�}v��O�>z�!�.ޞ5;�C�U?��/�n=eS�$��n7X3�s>��
��K��Z1+���$l�S�S^hk�ˎ�B�b��g� �n6U�Ѐ�v]���h�ذ�Q�� � ���zu����Oe���/���+1>a?W|C���V�c�[C�Ꜹ�i�(�j(����cT2e��KNd������HEvO���5�^e0Jx_v�i${^��+2ĻU-�2�w��T��$R�O����/K0Ve��x4�Z�n�ץ3l�L�:�"<���^hη�@�g���1Wސ�
�4.ޥ�|V;��Rb&�!���NTp��L�@����扲��
$R�t.�\�u_;�ȓD��ݚ%����l�d�>��u��^_,ɞ�Y�����A��^tWB}����ĩ��f��EY��LBtnӱ8�Nx��RXw�@c����`���B�dv��YQ1(� ���{��q����e�J��v��{n���u�����Nŏ	G���J���9_�I��U��9��Y޿l�pF�DmwoDnl���y�.T�V���b��7����}Cn�TI#-�n�ċ5�*��� ���;-�HG�u��Y�8C�%�J�u�������׋�8 co�5�5��_M� ?��v�������T�ւ>�l3E�|�o�,�ON;�}g���ͦ��#�����g�I��BY�ծ���E��W�N���\3E��=�B�ו+���0��cQ���AR���~LKp�X���LE�緃x�O���i[�f��y���L"fJ���"2���,��֏yM�_�V��][�N$���[ԩ��A?C����� ��( �X\� ���)�t��{L&X�>ʾ��y�zBI��7r�_!��[����\�I�����H��$���Q_[�31����g�*�6G�$�E�7Mv�B�W�iX��y�f�u�Lpk�8ʙ=m>�~ ��q�=��]��j�"7p��
zx��eм�k��]ڧN�y&��2ګ�����s�N����h�/l�S���oh��9Vv�͵䄊�Ơ��|�������狌�N����d���Y?��L��_�x�^ �R���l���`NP�s�R�t�T�5����bد�D�ǆ�K��9s���"W�#�#΍�ν^��ÿ�h���$�8Uԃ�!���*�����S���"�瑰*f�_����Ra�AX͜�L'�}�(����U"�Bkݺ���)9���j�C�rcZԚ�z��{�2�#����k�x?Hㄢ[��Á}�-R�����47�δ&���e�ҲZXY��7+�����T l�E&�
��"*�o�Z�g�����.���U��@pཱུ��?vyfHu�Q #5����	��؜���^Gл�R܍�~F��c7:���o��&rk_b���)��Bz�O2�v՜�q�5���W1b�?C��Zݖn�mg�v�:r��Lj��kO^íw$K�� ��{y}_a���9�p��;����P�~��%Q�Ġ6r����p��7����n$b]�Db>U�2m��4��I�p4����X���e쨳n��j��w��ًv��(�Jx�����yt/S���Ȇ��io4V��eF��[��)�
���8���-ت�E�E������PcN0@���io"�`�Ai��T
�����AP�;�Pʐ Z��Ǐ�z �rL��8(��?D�!�dqͣw%�����+q�X�Y9���� 4������O�f~&�����M��i����O]vu�=��	{�W�j~��~��H�����M�<Z*���Ё2>d�\{h3�
���'�$�m�ѹ�)���߭~S�'��3��DG��o��nL�(N���^�-9땸����W���`�ω����B��c2�e�B���O�j�}?��CF���i��e�ugv�S��!}�v����,\��U�'��� /��(���Zo�d�Dg�e��};m����!+�s��V���|~��qqMڭ:��n�7e;�+:�u{���M�$��wp��h���ٓDo� s=Sq�ԡ$;�O�ڍHYAR�DwI��Otv~�����b�V'�gR��Ê%<����[Qu=@�������i5D\�<c����v�1����4���|X�F?��=�j`
��/�mhx���\!Cx3m.�����1a7��"�u."�_i2B�E
��1N'�L�.�4����H��z&p��U1یa2����:��%��J��i��J�܎���{*�@��Mb�}�i��BpЩt�gԗ���iR?�čF�����i������dc3��y�s���=�I��1�.)&�C�i(��ŏ0Ҋ�`ͮ��E��u�O�Z�f
�^{�n�t8�g���s���%1��+vR�o���=,�#V,��+�o���b�b+��3�L����a��QNq���\S�{%���ϦQWQTN:�R~������Ͽ���\�m�����^����k�>��#�_z���v�3������ J����Oj�S��V����893E��&yb4�o�j�v��Q��� ���w�䝫,ֶw�3��^�
��|��F�JP�k��:q,[��,�!�B
��l-�x\Z� �A���Â���ې3xn���	p�Y�(�ÀdL��e���ۡ�P���?�f����^A]�&$�>��W}#ΠW�)H�m#䂹5϶G�� 30��C�58����Sg_U�
5��]Ʊ����~��·��Ȍ�/L�N>$᦬QGM�,*��=u���!3�,�!�b�C�fQ��6)� q�0�:Q��no����V?�F�_�]*|n�QJ�C�?^�1�uo��5�y{�1O�"���~�]�����4DG�B����#�X0�7�S/�I�3[RDZ���Aɧ\�8���Y��<d�v�T���C�U��YP�����e8v��rӎ�t��D�:�sVq����Ȯ�9�.��3/5^�Yт&��:���7��['��Xi�j��CΣ����!!�����X�vI^O�|Z�3Cu��G;����A��,A�f,J0lm}�����\�Q9�O�ւ����D�F@���k_/~z������nо�
�a��� ��s����Oo<as� 8x��wXz�F�hG�b%�/���]��̓Ƕv!��|a8��A �jj���=5�ٙT4l�����/VN=f����`Wq���ixz9�|�vϯ]P�B�Il!'M�C\&�h�U8��a('�}rH��e v���������b���+P��𶦃�\c�_^XC�=�lZ�f�����"X฿�r�F��Ҫl�~�l3�CI�M�r��'VTĴֽO�r8k����s�2i�:Z�7�� ��̎�g��70�����z���^�gy�䀔3���3�Nt!�
�<�ل��h������ytڛ+b��.gkgt�7�E"aI>�iʫ��`�˹Jy���]�ޗ�@��~h�T4�������>�j���'&� D�x0iu�)�͑!�L�j�m?�غa̮�����{����ɶ?&��&�B*���q��X� ��c�b
�^�#'F��QȘVȎ�[ �����M:C��������%����;��ڨ�xv
|;95��J�D{�Vh��ǁ�P��e:KsE�੭�譳	u��� �]L?߀��ؒՂ �[�-��KL�P��
��Ȱ]�SC�C�]̦hf���b4�P��R�{�0P2��t(�9;q��A���$9�^D���V>��f��j�γ�$�d�����Z��,7�Uަ^��/�z��Jj��,�yr�A�"d��=��4�������ߊ�,�4w��p������x3OC��J!r�L��YJ�(�	 m�ƞ�\~߈�CbY�X���9�Bz��/`V�F�DOWы�9J���>L���t�9DǼ�l��\�z�7��6Ֆ�*�}ST�[�/&I��!8׈� �ؕ��ڂ5M8a�ՆAc<}�6��w-���>��E`�H�M?�����nu#p �����\o���7b^�TE���a�=/�Y˻j�4ߟh:�{4�F~
C%���WH��*L��n�����g��̫shi��N{�ԶrC�M�j��4�s��F,f,N���C&��H��
r�g�Ne-���E�h�l!0z��t�b9(j�w�Ȩ�1��	��$�F��\����*;��f�nQ�	m$UJ �G"��^����՛<�I�֬��$�s�����dl(�,"��a��D�͌܊�HX�WG����L���ĪD��	_ׅI;u#/���G�F��B�P���\�L��۾�մ�1��pW�~���.P[���n4E�"?O]8�p��Mhҹ;�?��R)�R��_�g�1��Nk� �8Y���[�9ô��`��S�4|���K��U~�$lON�K� Ʀ����G�o���ؤ/����-/gO�Wgʨ�a��ȪԚ�a�[MΙ�4�R/��-�3-ќ�oI�@���x�E�����,a(����D����ڜ�$���<,��+������v6�S"U������qe~�j�a�#g~qN��a�˦ӻ�c�XE�
k�Mףg:�`�B�k��7K�Ni8ޟ
���W���n���8L��.
���L��b�_i�`/s��l���r��H"|_���k)���z� 5�`ztHs��嘤����1��{#�%����Xt�I���p$���v���$��1ӌ���T�s��Z|����!}S���Jp��6,�������u|쇧���5��px+{��&���]C�0L�Ɩ���S�d�,��0���:��M�4���|S�Ã�O3mLC��v���d
Ĭ!�|�28z�J�3:����v��>��l��HHN��R(�A�b�ܫ_27��9��6\�B�퓭SQ�~��Ub��O3��9f}9�\_���s��"�pЊ��G�<�ҷ��$�*���sL����x�m�y��m�����>9�+,*��FW��a�i��W*r��<̬�& �W��YY�P4+������xqk)�Q�&/d��1~OG�.y�${!|�T痄�av��N���ƹ��ls*�R.H�`��N�����y��t!WS�� [O!��� �
�͠���G%�5����?x]��H7Nτ�8�}d7�&ק�Ǆ%Í\�NKa̕TO.���r���:��Y���r�'����}���e Z�R��*y�g{�S1Ps4@!4�Sa�x;}u)^�=�Ϸ�Ψ�N���"&|Dv��7@`��s��6*Hx�2�!������A��Q���4�g$��Z��w�h�XQ:��:F!��E�cQ�F6��p������h�$ɘ��A(3)-#�W�f��JE�T��HR���� w������[�T`��$���0�*�&�������rGՐ	���� 0��v�(��`�bT�$��UA�L�p/���	\U��N.C����� ߰(��*�t~�&����.�ݳM ��u�m�2ý��Z1�l�R�N��k���Z�)�^�M�?{�w	3��C;=��ik��kx~��q���G��O8����v6S���������'�4$%����Wbi
��a��崒U8.3�@b���Xh�L��V`��h>�6&�}�0�}R[�ȇ�a�Ϟ�\��Z�XK�  ���_+�G��tѶ��IS�d������+l��u��T$�� Oփ�m;`c�i�����p�|R�+��X��@{�����v�Z9���g�j~�Ծ�#h7��=�\̓����٣��m(c�jQ,�u��rW�{l<�h��P���Q�eǂ ���>�`A�M{j�ƍ�������p5�� �g_�d�/�<ږ�����M�8�V�! ��4��DA�_�סH!�`YM#/��wB`��6��4���v8�$r�Q^0��++��=j��1�|'!_�����x&|�8�օ����,�1!0t��	�'($�M%���f� �!�
�"C�B���6�?
`�A56?0����W�hz���h��>-�AKxE���
k�dF�������˺��{p.�r�=�T~�i� 1���N	G9��ok����;����K�D��i30t�:�"V�' +�ql��r�����v�����j*N�ο;�������ꒆ���xz>p�?���ݍ�@����g�g�-���P��R=�xO�-��I��0K,'�%�a������?B�Nb�$ѿ�@�=�������G�>``�>����4u#����OA8۔���?��\��3"�*U>s���D�3��^9�$8�S��*�r�p&�ݎVP s�@q�`�5�]RMi�:��k#�}1V�cyE�S�9����3���.rځ�ĈTJ� �lBy�/���^t5��ۡ:t��U� 9�a�� ͌�%S���7��=����	�<`>]�o����*h"IK�&	�(�oF��@�z{�s�I]�x����E�L���m��y���3<q��$Q���%���l}�W��'Y	��u��HҬ(��'��/<��]��f��l1���73?�,����.v9�,x�Z��q�(�-�.J��I��rȳڛZ=Ƅ"����h� t'����+�a�s2���n<2�=�wl*f�q�:U�T6m�u��\2������˦;SWύ|V<��f��;8�>�W�,�-��F�B�u,�E�<�G��_��,���cݧ˯p^T�k�����M3�DC�Fg���л��<t~�I��`f��f%l^�1�-�*):��\md��~�&�i��ﲧu3*2;/dN�)�h��#���f�H-�5�4F���1�ꤕ�n�賅7���na�{͌�a�\?��,��b@�ϸ�1u��d�~�3�U��c+Db�yw=.�/��[}]�����&RB�m�"��XO���V?��������m��m>�TwK4��Yh���ɛ�5�'�+�qh,�;�x���$���K�hp��#��5�����tw�m��0�O�5�Vќ�GC���%	���]6�	�N�R��I�j���5��bR�� h��~�Q�8������:�b��4_<%n��j�s8�[���'>}/ġ��fW��{Xp��#Z� ����u���e0�~L9Х�?����oLYj
6��X
BQ�p?�ۜ� E�^�:p�i��?l���8�&qT�y��9�j�~O��C]��u<��y�rcaC�F����5��Z(���,��0de�/1��� 3�)�Z{B67�k��oE�u�e��p2[��ZO+��qX�I4���p(�^ڵ @E�Rۖ���c� c�A-+4m�f��<�y��W��v��?�a��=������W�W� 9��\J��Rzڜ_+y���FNٖ��(�{@@Ȝ��^/��j��s��[ra�Ǔ��Xv�ע�HK�����h�+@�ݞu�;��.�%\2�v⵱��*�ݧ6��2�O��2���b��2X�Z��=�4;�S��i�Q�\�S��YBWtȫ��=i4u�b��k�`J&}xp3I4t�g½�l��UEmu�>45���((�|�6�N7j��}�ag+�e�&$��l�a[�b�֘�Ǝ1����:u�VN�5E��@3�q��ݾ�;"m<�yu�D������f��L%Z�L�-�h@�F��ցK*A���B����)LԪ�A��/ו6��=��,SsֱW��w#������EBu�Ju�2��[�YG��%#\�Bk7&2̍����9��J�I��������SKb�2j�+��2���;nk��T���n�fD2-rR�2g���U�ߪ�cp~�y��`ᥱ���i�=pvhI����B$�p�ֽ�$K��M�g ���O���%=��e�����������Bq����s[ыSЫ�x��[2$�!< �D#7u�iL�Sé q�������S���űS�>8��K.�3�|:&t�5��VfM��:��Z�P 7��Vr��Z������)��OhiF2 O&�,�!�gJm���m<�`P4���Pڰ��_�t�����Z���zAF��Dߔ%���޾�1bGXgx��@��xzQ�1v��H��J#^��tS�������_�I�ג��d�����8s��hu������j)OƩ�rט(8>���ߜ��0I2"��a������=!gg��JJЂe����[ޘV,KC��hy{F�
�Iϧ"�I������K{�/#��W�ߙ��X��M�=�q�٭����޴�6b˩y?�?^S߯l�䘀�,��D��p�	�k���[v��LfD縭��X���Ya&�p��:ģ�����=�V��U��A�;XY_*�l�5�)"�S@,Ӡ7 9	��j��[��0a���ǩ��閣rN��%e�q��J_Am~�0�qlTl���/��Q={��>��/ռ��6�N&�E��ok!A���_�Q�q��z&I�D��*�d�G���`8W�W�f�qRp(qƣ��o�n��yj3׍S7�m��?��B/�)^�]�C�p��q%�|G�~���p_S�Ȼ��ª�_�p��M��)9E�%~��tQ��2_������+�}���ԕ�7��I�mbDڍ��g��g�k�y�$!��_$?�v@�~L�}�$������ɮD�Q��u��sM�3�6yrxz;ˇ<�,��Ѫd#�~�g�w�U8���0m��@wϐ�ۺ� �ؕ���<P���:�����g�gS�0tg�cl�gw�/>I+�(�o�>�]�8n�<����|�R$�Xl��BUz�$>:��Ic`�#�� `z�/c ��3�[�!���;�"."��Ag�
[�51�@]�X��`Iy�����QmjTap��e�,{&~7��*��U�k�dJ(Mdm|0t��`8�(g�R�]G\��̾�%F�����/~j��D�HϞ�!,�<���ߎR3�|��w��5��=���q&��v�V�>�q8(N��ొA���*���������o� ����-�d��2s��	��'�Z��zv_9',m|7�dS)�Y��v^���$ޑa:t�㱯K�
%L����A�Y��zC<�b�';o�^y�̆�!�r�� �~j'`H�N�¯8�L���ސW�}�}K�m����	S�C:�2B�`������<��@C�~���3S�5tMc���~&��z��R8��'C�XF^�3J!�O�F1������/q%�h�2fYO�?��L��)�]`��d���[�J��>5#�}#�2I9��uR�^2���2���Nݤ� �����e�&[�n����u��	��)-J�辌O*�A��L�:0��o�CnnV�K�l���[�R��U�{��������|���r8���2���]�q�����,��%�4�s,Q6����~3	%�-\e�JT�f�X[�A9�������g��d��AVigt�1���USKa�K�I�.���3Sj��[�V�9o����$�X�WXSw����u�4*>�eU��a�}]�����ӿ5̆*I�A�ו?���&T�J'�doC�5w(Z���;HB�Zʂ)�A�A.�e��{y@M[s�Z_�0���=��Q<�-����������Ç-�Dt}�Z���tbt�	�����=�����@pOz�����fgܔ5����Jh%��Z��&Sv*�N{/�b|q0D�jC<�c1��E��#0q��/f.�{1�:�[*7ƈ�ET�Uy=W���8#KyT3l�y�r�{��z�c���^�����n���kg����g���RuR���H��I	����r~����Դ� �r�T[���5Q,�a(���Q�N���Fq��NGy��Qwo�j�o7��3��\i"T	k~(�u1�Kσ-�=�
h�|6ڴRuR��i7
i��u���mǾ�1��r�a;�()h ���@0���[)WG���u�L&˒"E���ۧ�P�������#e���Vއ��oiS&���j����1���	Q_Y>)Β������Dnt:0�`u&��8}�����Q��W;T��u��u~���z���2�C�޴�ۼ倗f���é����u�b��h��1�[�0���%���H��ɡ�e�j�x^N��Ëy����NZ2ɫ�<��Ie�{��Ҁ���r��yYӷZ�4���M������1O�)����\҇E��g����<�I���&P
	�ho����%&��?�L����
�K�t��S��+�C.s������[��ek�����%\��m.6�T���_̼��6ǔ���0�t��R����Zs+6$��d�jq��J�=�y�&���H�:�u�; ��u���O��?��|�����7N�*=�v�! ��Z����vć�:;K���p��>uV"�C"$ȸ���#h�	�^��Ȓ�N��gW���	�F�Q��bҬlY��/o2�����1�k�^�:�BPG�/ +�Dj7U�Ų@]��ª)���P�L���}���ʠ�&Hv��	���S����}cy�v����gT���F�R�}��鮙&	E��`J�ECI}�������x�~V���[gh�7I?�����<�����ya'^����(�[��dV x�Y�Ν�ۿq��z��SN�̖�^�M�$���!��9�\�����q�k����(vۮ�~���dj���q��x`��m����LO�p�Gz��.�B�`.˟�L�'��ky��U��L��g	���I��Lc;#W��@M��K99���Ѐ>� ��pۏ���={�n�]SF��D�������.dj�6I2^����/@~Ԓ�.��,�C�m[x��8�]�FݰĄ	;�����uo���%��y�X���\���-�=�gОQP��NQM�{9�Z�]9(�V�{�	~��Z��U�i��d��r�Ňk=(y9RW�¦��"�-ԃg��7��w<a��o�F��l�ښ�Ż4\]����q7�y��g��l>K����w4�����k��=?�v�0�[����j��.owa�p�K9� �~{�K��pj�:M$�ZK'�<#�Th�ٗyr���^�ȩ�{��Ĭ�r���m����Z���{I&�X��xW�Mw�ڲAmzʤ;�r;�f4��cGr6�d�5�'(��A>]h�n�;���v%p�1��4�ܜf�=�
x/B�����¨����u�! +<K���ӻ���0���J��N�<+���3L�Ȩ��4���%�G��K$��Ѹ �iဥŞ��XPƄ ���5��<�۝[�1�Dn�J��I����週���O]�n$�[��GDVB G�i'ԗ�`����`J�7��u��u�����%A��Ms��9�g��d��u�ز�պ�۰�Y��rɜr�L�><�<h��?`�É؍��ˉ�AǶձ��]���'q��A�D?��U��mUp�t��%��W�Ek��4jqM��hԌtw��(a*C1.�؀F$%2�7�:o\Ϣb��'(�5*���O��rt�mQ,Wq�g�Ze��� .�����SQ���/���#P)�@!G�g�Gcf�����v�˸T_�-7I�~�J#�zP}��� ���pZ7�pc���������:�5)�{ꬤul�(_>�8|��4�#c�������Q��w�EXe\0����W"9g�Ô�رI`"���JCI��W�ۿ�������vğ��Ț�̓�E~{��tr�΀V�ҁ~��(}$1�b�OF�c�?�&KMfd,8}X�ᣀS�����>�w��-�"�9'�TH�*�,x~��Si4���
�xZ�H,����Х+�a���z>w�x/��{��4c]�w���.%n���p*,R͡��U��I�Ґ�ͱ��*zK:^�Lw�3�2#�w@����y=I���L��n��b����J_�O�1f����nh@�$Y�oh��nB���~�O��OY�#���b�`���0/�[T�ɠJKXnT�:�����[o�s:�>U�H�i�+8!gÐx���$q��S�:a:����\Yu�<bW�rR�3���~�{��m���̒�qx?k���d���UA�5, �Dg��j�S�a�1$�[<�A�˩����8�
R�	l��	 �KFs(�x���4aB+1��\�������#������G��v!�bܛ�*�|�VȳanV9$�U�?w6�]���"\�`�,f%5&᫖�Y�2&b1~8�Wk��0ᡂM�9�l:��8^��@>,��e@rG�M��(�.�`��J�3O0/����2�v-��B������7�aP1G[4Y�`!c�(���u��a����o��ڝ�4<	�}���ar��Pg���FQ�����ۚ���2Q�r(0x{^�l��0&���o�p
��ͻ/���oL��X���.�$�]�gCC��-覟�����C�'������ki;�A��E����0ISm��Uܛ��|넷K��Q�:��5KR�/�e� Z.�"�oPw���!XR��LC�Yw�V�7Vs���_��/��r����A�+8g�IoȀ�X��Z���Ĝs��-s��螯0���ኀD0뉦��3?��6`E�^�����[�~Gww���*$t͇�Lè��;L�ãΜ�댍�Š&��>�T�(5�HG�����X��5[��ؕ�LH=��+���J�ȳϔ��De��&v�M�	FJ�I�oX��Z����\���Ԇ:�.(s�N��<H��ce��`�������FF91=*O�v=f>x�K�LфM70�
��j�K�]O|��z��;��)ޯ&�IP�5��J�ԯ(չ�^����'�}��l]M�E�R��4�q��=B��e���^%K����W+�����������-����xk
�?S�B�E��M�?i��'�����ϱu�T)����
{��f5[�MV�֔u9�m/x�u,�";ő�%4=䥝�/�Q[}a��`^y�Y�m��l��M��Z��"�ZO��=})u�w���y�%�h�wB����w�+XV�q�!AE?����GO��K�V� ]V�ȴ��u=eH�u���#�ؚ=��]j�NIBFz둫N�;cL�V�L�*��}���-��	wR�G�A�'jllQ}����~�j����S��T�����^%C/^w�C6�%��@�͝h��r�m�������ᝩ�/ת��:���͑�����
���i�0h_Z[�m;e)ekq�%��ʵ>��#�1�u�Q��ڨ?�[�lԛ|]�}|�[m}&�92J���W0"׷j'j+w�ӝ�K��B���V���yp�n��	�f��,��ϻ�D��(����2ە\H��=��uE��0b����dI���;鸣��&�:_R��.T�mPSG���^�$E��WPZ���~�L��'eE����jo�bߩf�<U�~���5Ơ8C�Z�L)�q28�[�	�������n�٤���s�vG���-}�N�V�D�@ˎ��[x�%���ў3{�2w��Ǜ���s�4��?�;4&	�oA�]z��1����g�-qԚ��
�ο�K�_{N�+4�M.G��CN�RB�d��'� ��\5/�����=��P y�纖���!厍�17��nܙ�3���7Լ�V���3��7<�	&(�r28�ujo�6{���P�Wk�L�T%�x���A�-GX(��|nb�V:Ib�0���e�j�C[�[��;��j\��K�_�h>�LNdf�n%�v��d2��$��c`(���܄�n���Y���G���F<�L��(���gm,kO�T�����.(���;ؾL��n���tI��E��H(��@�6�-�9�̌_cT��	6�I>:!�ܛa��@=%��2�'�k���������c��@�7�r�d`2��8������M)�@�$��Κ2��8����V
����GWez��f͠�$������y{o����叶�� ��!OyV���V}a8��4����1�m�;'%��ChO����~�h�_A ̓��/�5\�x
��Pu�bg��d�F�� 癹O���d�2���Y��:�����W��RԜa�Ogr3P^��}WE�ɽv�S�%*5����7oǾ.:�Pߓ8d&ݘ�O/��^{�?�XNF�ގ��us�] �<��33���Y�%�(O<�'�Uύ͈���c���j�Y�[gTc�1쯼�=�K�(N��m�-K�7�C]�($Q76��,M�CN�d�G����Kp�y9hv^�������;��U��WP�Rz����
)__C$/���g3HFp>����kD!F��"�$��t���}uǫ]J��q>Z�"N�&�9������:��=�d�gK��Q��⯡�Hz�\�Y�� �B"�N3�(�{_m_D�izN�|fH=��x��Ie�.�����π�3ui��5��]hW�^��-q��	���Q_H��i4Y��o���,5E�E��	@^ٿ�vE��R�r�{�Y�Y�Hu ��~H�aRB��k�ښ�">�����%��d���Pp��vF���j��`�`����QP���t�� �r'����E��ǥĉ�����F�0{��7��r�y���y���K��vM�9I(��ZeܥL���I�������<�6��#s��({\e���QΠ�8By��#��Dc�����	��۷vH _l��kDY��_��l̉�����(��!�|C�W���c\:H+76�t����H���'`�S&��D��~&�t���c��*�9 ����������[6U��P��Nq��g��d44#����Mh#�T��P��>|l��oڃ.i\�7C���&S��	��3;��u������nb��,�������-D�Y��B�2���Jl�	�р�v��e
:SH����|ߝ*�v��76�C�YLP�%2U]��ȅ*�.z��z}����iSGϭ7�M�"z��W�Oe�p=e�`�]����0G_�)����pm��=.�>�_:�9����1��`?���%Oq��b<�]f۱ě�f�j �"��NT ��^�ae!d ��6��7��0^�,v�k�~�'��|��;C5�4�\����MX��+�%�{o�*�_��ۑ�A��><d6�9m] %*:�C@~���E1g�����:�X�e�qL��F�T�^�IO��ОZt��ogn��qg��^���;b-4};	H&ȯy���ȥ�E���+9;���ɣQ����3^ED�_��H�[�����#Ht�o�&oK���pҙ_7���~mjx��Rw)l_�`k�%������ �h������iZ�0tޗ}�y�M��ll�S�=J3O��i~�i����Ch��xi�԰���ʳ�k��$���c�@��an`Ox���}��|�W��w��ܫ�8��y�
�.�h*l��0���ڠ��<�Ǘp ��i�^ѳ�$��OE�~{��<��@now�/ �/����{��oB< %P���Awq�`1�$�tU��F3;�����Y���*�Z�#1���\���:�ǣ�=�������,�OkX�yN��R�܃�=�G��iFr=6ĥ6~u��O̞�p)�W�x�2����H?SOx�
,s�m�����]�o_�y@�vGP�c�ٍrC+^	���P� 	����X���B�ʹz%cc���Y��1�Q��g�����y��;�魱�*�1�L�a0���V��K�$U\�ہK?�t9�:�^�}�_�'3S�6�q;%\�q��}������C��/+]���rw�f��G�p�Hu�����
�����W�Nq��H�Fb[�M�x�_?�ҕ1g��{'�;I��ӿ��j����?~,��Vǖ�%z>�J}��_�����Z��Q�:j7_gH)�����į6���e��D�tgQ��(}ØR;Z�V�^g<�+b5�ΉSB�ְ�V�w��!��٥������Y����3���o+��O��~�4�=��+X���&Z�VM�Q"��Lp%bD0j���I®"����ك�6J ��}7���7�䢂���+����Ng�<g�D(i�=�b �ě1^��lI"�@cj��-�7#^��'M4T�s���.Cd�#X�Z�k�h
�Ъz\�qȳ6��CM�S�Rt����ݩ{��Is��bʍ�W�Z032Y��G�D;�jv�]�����=�_X\}cQ�y��ױ˕f���82�����L9�1�&��xC��0�ߛˌj|��F���
�5,�g�.vC���8���������Eş7�����nZ�c^�&�q�k��B��,�D��)�A�W^��6�͉x���sW�4=̇��&����@h���7jQVb_�܆�ǌ�����X�Rs�#,BB@3�FF��*��-�ƥ�}mZF�tk��a������p��a����z�q�蕩�
F���,al|�a1����ai?q7G�(o�~2%q;(�
Hx| \���L�t8�[�6j�~����9n%v��nv��J��'��Q�`0ƽK�W�U\
�* �?桼�(s��bҮ���֐�s��`��}����(��~T�9����Ή�ǧ��9�U/H�	;�զ���8Y$�h�+��Ը���<p�P�4����Q�z0�y�ɰ T܏���A�	��Wr�R�  ��+j7I4A�� G����� l�qozQ{JN0�����3-,+|Q��#&�i~�]EH�A�z����m�)�u�f�c_�A-8-#������u�������H�6��9<JY�]H[br2P������!����p��K�J���i��(�E`���޸��ޟ*���hJ'm���^'�pnZ�����e�T����ŬI�A8󙪒�g�L<��]!�������Ya�� �����E�����-�u)��ʡ��u�P0���ϱ��)�	���_c�
ش ��ҝSKڼ=b�3*=��k�����-en4û�K�]Z4~�	:�B���O5H�|�՘��(�0�u)�2��Q��m��8n��Ӑ~��ٓ���9Z�zȘ38�)���rHb�tXwq��/��g�m��j�v�[���k�p����U���dM�S�������Y�c�j�'#�
�_:�8N�WM��J��y�gѸ�yb����Ԃ�G�b5[W\�`X���������F�5�t;�W8�:�����K�_4=�O���Xi�����o4���wSn%0�������͋����1�F�7�k��X�&;����p~a�Zj�*�S���o��#���F}�E�e��~�FS��D�����}����~_9�T?��.a��ŘK|�����e�vVu�=�����Ut�槺*
P�B7�a�xi���}�sN��x�8L���j7��B��x��SmoG������a�Z�&�Gr��d|��3y�];P��I�ڡ�eb)�<1)CUu���?s�;��{�F7 ��-u��Y��}x�|��d��i�!�3뜐�K�϶g��9� &��9a��!�KE��mW��ٴ�75����v{�m�M\��A�C#�}��L�z�*4N��B�57h��v>�0�:H~�phᩧ�nĺ|�|������8~<����l�[�E��%À�nX5<�E��uF:{.��GM����Uip6dr�kZSq�0FXq}�-I@(+�4�vb�ٶ��V��MY�����"
T��m��x���-7V
 QG[���f����?$�0��F��y��{g_Ry�̯o�c�s�n�9cW��&��I��l����k��܂K��qn�q��������o��O�J��Ħ��(]5�]�Y�.����W�v�ʤ2�j/V�	���!8l�)O]"�,V~���P�k��(� S��r�_��?.K2��i�ZL���	D!����af��.p!@�],w�>��jVeb.��^�L_P�f��⫩�Z���c-����tkz���V��Ԭ�a��OD"̲%鉣�V��\Ó�Q`�t����4e��MC�ԝ�/�}в���J��|1�TW��O+�A��;wP��fu�!5_�\T��T}'T#wQ�H�����d�m�ڇt��p����z�Og��r�q��ume��� ��t�#�k�1
��K�I)Ď/6=P$2w���a����2ٹy	I҉��: et�Ka�`��b�.6�ZY�iy�� �=YQ�WΘ���UT��-]1�r�����t�DB�(vGj[<+����r�w`��*	<v^�-��>*��ط�Q��E;z�x��~@7�n_��EǸ���͐�ێW1H'yJjn����u���Ue3;$��7V�d��.!��d�c�厱���ʱ<^o���Jf_v���>+l�"*�`��~�M}/k�I�Z������s�nuY�����]�\�Ȑ*�2G��������0޾�8��fg���K���X�a�g���i�cM ����T���s�ͻ�0k��*�D�I�Em�8u��o��}x�'us2[q��@Y��E�����h�)�tר��j܊�[��o�j�B�lv2-�d0��&<����)�vF�#k�W�0��)jP;/jf���?O�ف
�1[#�P՜�ZZ�Όӷ���@V^l���	
I�LW��;TȊ-=�IL&w�)n|�Cf���w���`"�&.���R2͎�A7������)�G��TJ�+�:��xT����������%Y
�~�* ��h��9*dKQ���p�ͷ�>��?��V�-ُ�c,�J#�٤���8��U���fq:Y�.�e����x���Z/�)L���:sY���v!���QY�������g�ʶ�����v�95ˌ�t��=LG�H��%�𿗛�8ڬ��YX?�&���ώ�^MX-Ք`v^Yz{Z�����p�$t�b�V����CHV��hV T�y9����4�?�b0�&��Pn)?<����J�,�_����!�8JM�R���l���"�����E�8]�,��7���#w@؇FF�O�Y�ADV��G���އ�u�]^�o�xn�A:��9!�3u25t�ll�!<Т�ܚԂ���G,�����\1��Fd5;9P���Q���?�����h"	?`��6>:8���$ �
o@�1F�N\:@�����8vĬJ�w$7�E�yN�QYP�>Y��`33�r��4�F���a��	i�@�[݂>tLx��d�8�ުj��.�gQ}3
L�7��V� ��r�|��]��#}�G�h���#Ei@0�M9V>���ˊLy�B�2�LA�k��Uqn�6���ٓ˯d+s��su�����"%gyd��|(�wJ�++�OR �5�_�ŕ����Z��?o�̜�K���ˈ������Q�s�UN�Z��U*����\�3�&3��&�>ĸ����>.j&0��)��c����0����KL+���#���q�-��=S�:��.����o���x*�����ܚ��I���~=	d�8t����`�n� ��n�g����Ew?��j���鸪&��K��\_���/8���H��fU�7�Y�� �+��Cޥ��L\XS�l�6�{��I7�+�1�beJ�t���Q�E�[��Ŕ�:�޿��g��w�0��|�$}�Z}��"�h<R�E�
kg�4a�#�.4+��ȼxA�B�9j|P�/=��m�5��M����?h ر&i&�H�QTz.��*`w]%�=m��B�%x��)=Dz@=�������5'>�ơ�����!�XPt�Uʲ� �������史�P���}�k4�m�3�	�����~�8bs�pw��� P��󡕮3FN�Gg!˒X�U��=@iމ|���C:``Hz��z�!���~vOQ�w��ˤ�u�5t#k�raӉn���{�{�)�؂�� C�4n:�ϣ�+ؿ.`�N]�8��H����z���T5�� ��T������E[<˹�h�.Luּ�P��7�ke��_N>5��&�칚���n$�w��iLdC���+�7$`-i��	��/G�#��M�����\��F<�s�r=�+�̘�z����K{w���X���o��,M��p<�|�!@��W��:%�wR�gb�b{���l����T!�	���	�۾���  Q·���r��9(����rh��՟�%�����Q��Q��O���z�CQ����2ƃ3���ᄪ��#�t�l*9a�V���b$�\pp������؉ T�g�Q��	���0ÓBq�v���	9����Q� 
f�? �4��t;Gr����mv}�+u����>��4����7���5pP+d�=y�f�����n���:O�F��E;ĳ� ��Zǻr���9�o�� :ܡ���R
��`y�Bx�*� X�:f�i	�p�X����^`��#���2f�Ys���&�b66�=6$K��>%������Y�O��ۜ僊%����i�<�2>	VYUM;M�l5���F ��~|^��%+,�Up�p����@x�<J�`x�U�� ���SJa/	��?Uu��T��͗�')?�v����)��n��XRG���	;�C�/�?�#�~d�K-�I4r��+�	�A�_����ǹ�{�l)�kס�de0^&9;���s�Dz��~�YfM\4uq̪+W���N��-p/M��~<�a��*�[ Q��]f�����D�D��`0/�%�<#�P�|�(�R�2�^e�a��%��C�o-�+cPg�F�C��bVt�U��\�g����� ���ɖ�2�%t���`,�[w"���֓ �Q��l�VFJ�B���s�e.�f4�Aj?8�i%m��
�M�#J
Cn���:�xJ\]t�a�\$�����<ϋ��j��%��佝��� �M��瑳	��<�F��HW/f)}�K%�K�I�Kη��b��Av���X�#M�_-��ԤunuhN�&�^�lJ�G��d�����gk�c� ������6!Bf9�N���7Gu�ަ��v8W����Ĭ�PxB����f6urt�T6����YV���:Ѿ/��nY�4Cۍ�$��ֿm��FS}nb��0 P���o�՚9=�����/���g�1��UX������1��:D���0i�j�po&BJ�pp٘0�q��lc��x䊱,���c�tj}�zaIpi5��o6Drc#�W�t5[(�B�����ͅ�NU'��@�@ɡ�B�&��Yh���H�2�xM���i�$�cl{X����G*��; �g�p�8@�N,�-�L�m0�z<����b��Y��N�?w�V�P//%���c	:;;������H�˦(���1!�_4��ևg�Ʌj�����Yo�2�D:,L��=�z��ם�5I���W&�*�Y=���/����2q����%�^L�[��@3�+���Q�}����}擅��!�t�;�;v����a�Q)J��ʌ7?iSŐ���a�Q~�1n���nx�\IwU:N��L��On�`Ͻ�Z)V��4jlH=�I޻^ED�
��nt��n$�x���T2�+k|��}�71Ņj��Ț};�#k\Z�w��;P�e�1��^���o���>��H�J�q�!�姾�}��W��Y8_𼟈D���g�I80q��F;��|���Aְ�b�\�P��G�1�ҫ�_?).UU�8��K����o8-���Iw|����0��{�C�+��=�v^[ZC,o���(�u:��WI��2�74f��ǁ>�z��J�f�����U�U~	�$594�+�մ�B6:�c�h.�QJ?脯�0~e-��
��|0��@�}{�`B��y�"#]�Q�>\ �@�\��R,�a���f�:�*�+�����O9Y3����Ow�-/�\i�q�p=(���5Xu��.g����A����ȸ���g� �<ũ�ݻ���R�12A�Wε��k"&p���".nrܰ��1]f�*3�P��!���r�c#�!���f���n����]�ᚤ��ka�H�N�������&�6�K�3��K�4
t��1n�k	��$������t��x2��6��҅�˛��&��g��8�|Ȅ���һ�P�k��y$.��6���+���RSL��|k��Q���k�� =�RIKdɘ�6�1��a��Zщ�K�������<^�	�H)k��wG����B@�ZE����ıeHL� �Ύ�`Ϟ�|�=��~�V�VG���A�.!
6No��_a?�쭱Rb��bW��J��!�ӎ��\[ܿ~�jXIҫHP��Nh�"��Q&��E�6@D$F]S��/�ȷ��6�j�,��9�\��C�m!_�TG�}kF�a܍��-��U�c�_ f���B?���W����5�S*�qex�M�31��b[�gHs�7F�߰fts�K�f��:��������tu��$;�x\�u����DI�=����)I!�I�J
&~癋���i�󦟑@X��
QI6��┪.����O6+�w_�f��n$��ʲ�=io$"Pj클?�����2a�j�3RHt�b=�4��L��i��9���A82���M��!~���7r�4�2�0"���H���,A�\�h��h��G$ưu���B�!S��γ3�������0˸$��&7ך�]�G��A��mN��̿���.F��{ӰCH�.�._sː3t�^]y�:��O��0��q�ǧkr�M��rY:��$��0�o.(ky&�[$�4{*�#�"�cu#z<0Yj]�Pث�[|P��oH�⼨�2y��qI�����H�������]�$�	%���8�iD'�����]ZIyl6��wx�~�I?�����OzI}pj�/Y�.����5��^G�zC�<.��-����� �*"cu��I��~hL�p�܁��5=l�'&>~���k&��B��� ����m�"_�E�a�:`/�K��`薇Xgԗ
��U�M�]˚a�!�L�@�J׳MeJv��nߗ�G/�9k���j�Ol{x*�G��a*��5Z��c]n!Zf\c���A�����n�@��h�/E��Y�m���/x,n{0C��tg�s� �xGא���2�G��{���̪+�<����Z��p<o(򑝠?=�;į0��$��:���1�G�+I���|K�\�z8��^�
+�36T��V���������I$Q��[��_V;�j��X{�њ?��7��<r����&l,�D&�y��mএ]<SB�
>τ��Y�9�����｝G����L?&�w�\��ȹ�/�����n��dF�#i?uw��IZ�Ł�Mqҍ�_wh>����ފ�b[)�3@+e���]�qm��Xh��=�%XJ\k�F�J�a��f�(,ERk��Cc��v�����T����(=�����d���S�m_.G�[h�Ĵű��s�Nbmb��[�T�ջ���X.��������z��?��e����ZuC�F�A����B��Kh����;�_��
N�>�>���?A�n�!��m���B�0�'%%��J�k7���-x��Y�9��WIy:0H��ٲ���)Q	�<!���$��V��Y-�My摐c�XR۾�	��S�afq�݅�%4VfG1ѕ��V`�Ɩ���"�]Pr-5�W�}��S�b���7O¹�}���K�c`��8���Z�X ���*�J^�$Ÿ��E��ݛYh�¯�pҟ�T=\a-9�X�e3N����]��� 9�b�YB L�<�4&k$�����������/���j�C-1:����s�f�
�j�|��.y����:)�%xlJ�� �ruO��Gϻ���\��Z!�n�r�d��R�Q����Q@��h��Ęd�I�0	6]JX�QR-�S�QA����Q=�'�A�̑U�W�	 Ls�A���~��g �C�A�8�a�غ?j�i$
#�ruW~�3� �#�A�@���#^B�k���릺6^h#n%��P�F�M�2�&g��ONz&�Rܻy`*&1ũ /�ũ}ӦFMf�#�����a/�ju����5�X"��)���c���`xo��`���EG�XI��E��1p �S�~���|��m��]�{UL������PpBm[cf�M��Z}�~{��t���ޣ�UVK��D��+��v��3Rm7Ｏ<_v��>�RRV�|v��w ]�텆�Ŋ�<"l����r��"��{����z����&�?!�%Dd�d�J���ԩjA�fƙ�z���i蕇+n��Q��OB���;��*��xL�f�YXI���[!n���#[9V-�	<�" �f�Ǭ�q�	��f��&V�I�1����b9l[/W �V���W�C9�~<����Z�����h���S�-gw�%�D����h�H�?��1|��ø�"ͬ,��w���!C���k`�NJ}�$+P�C�%OC��Ym:�W(sm츥)�!|��=<-Sp��wb�nG���B:��h��]x���eާN���o[��Q�*Ehd�7��}>)π����`�1/�%��V><��Z��+ix�w���j��Hl)�Y*U�紲?���6sEXy� kh,Ɍ�R���"-*8 	z!����[֐�&�z�{��{���N��A}�pࢎ�ܨ�/EN�_7H�S�>.M^Mk�I�7q���*28RpB��Au	����SN����n��E�̀EN�,6�8`�V��U��ʾb��������SС���gYh2u]�Nd`����|��VJ*�&�H��s/l��U��nez�"���;���Z�8Iatue��Ā�e%9��B�w�a��u�B��?�*Q���yDܨ�xB�k�Q� g�+`�$�$�2�'��V	K�9%�ѹ}�C��S��X�K� �Y.�h�%��?[��_P`�����⁇��Φ_���	���djբn]K藸�5~sƢpM������P �NT��8:���#Gm���ze��R�Y������$lZ	���#����y���9`Ap�(�a�� ��9��O�.LxF*20�-7N�N�x{&cw^�T�����d<5e(��B+;<��3��Zs#�2�&	����)�/xu�*m���&`	5Za�D��u�Dz
��䟳,�a�ܒ�6��>r:h�h&��^�������L=N��bm����� �jb{GHe^>G8'�|���u�� ��0aot�&_üT����j.���X�m�JK��	�ZN��;O������6;���-�}�$��Ƥ����y.�1�Sxa�c5 �v�Ǫ+[�~���>!!�^���rr Y6C�tNd\�ZE����V�-�(K�����σ�~��n�ۻ�+������
�W�_����^���<�/��N?���N�g�r}�&���&�
�N.D�zĉQ���]Ro��]��R��E:.{�~MW�Lk�5ͧo6��[�?��&�������m�T�p+g��D�/�5�H����Ni����}�>����Jjl!��QA�>�l�A�g��m�7f\F���Ǭ�[e��x��U_��f	�J:K�f zOg݈��o�]#|{�ROS]�� ����nA��f��آ���#b�ԟ(թ�/����h�yc�{l �o ����?���:0��&Y5�\ɘ�\K=T�������=���V�N��+;��he�F�1�W��}�����7���u9Z���M_S�����&dV��K���4����$�?`.X���e��jاR�vzn�b�qF(������Йݬ.�[����]$�H�v�^!���L]�5x��tES"� 4S	��Ht�M'�L����\��w��p�a�]���Wbs��;�'lc9J�*Y�&��t�DKh�h���p�3���w�J�� ��.��tt��)��eٮz�x�vt��2zhU����F��2G4���S}w���7�#���T�L���磌����n�����!��DsЙ18�Ă�����3C
<� a�ɲN����th�c͜.5(���y�F���Y�3^����=�O�o6�"�=3(���>���1�Ж��}|)v�/�<�ܳx�����!���@Trn�ax�;:�`�N�ip��m@כ�r���U݈�ܑl��h���L�������c��:=5�}�y���%����=@q�|))c�>�x['#9w���Uf3۟'iK(�0�� N��c�c�I�Y������ڦj�C���#��f)��3L �g��N�]xǛ�-��)����+V�S�r���SxmKk��n���o ��NΣ�I�M�bH	ߺ�^C:��kM]t�&t��=�|U�\�X��j��	��A��d�/�H��,���a g����,�P��?�/!K��g �s�L!� ?r�`[�D��f9_�#HR ���l�Ŵ?anE!�,��8��>Y�+h�W(�,�8�����+p�
�b���:`����ei����>һ����>+�x��%�l�-͕�B�I��u� �%@��Q�H��K���x���>Kke�����
Rp��Z%�N�{��Y]��X�"���bY�	{�砤E�G#�;	�҃{=�ܟk]���7�͉�7Zy�\m�l��r������l\����M�of�m����f��xb�C�+�G�܀�Ab+���-ϕ�G���	���B�#^�[kn��Wd���lD�׆r*B� sZ��f�r��B�~.��B���tϮ��UM[~J�d�*6=!��g)f��䪃�Gk9���4&��;���_;���nw���j=��d4��J? ,��j ����p���xw���&�d<�U¯��� �<?��5k�v�t~c�D�<�%��Ey�'~�,� S���=\�,��M:�Z����$߽<(���Sv'�Ǚ%�X�a�R��U3����Cր��c�����D�c7x�`X�iX�I��5�CHP���׾�;7�٤)6T�߇7�Y����/���V�U���>�SF��YL���K"5�՞�JKk��o޲2�Q�X�J�?S�w ������d֚eD��k��~V�E���mCF�^�FC��'��[մ�}=��i�eIXͷ�Ը'ߟ�^ ݻZ��rl���_խ�4��+�[���W�g���7��P�]��[M�����/�����T��'�^t�,y��+��#<ۧ�t�j8u�1;��ctæ�T�,V���n�U�)�f m�{:�o��V����7�Bbz���	�N�;%wz�M���#]1`n�4* ��I�K�".-+�6�pF��g��]_���=r@���E6��*'�qۗ� �X_��<�?�S��WYu�X�{��j�d����/�C��tTF��{��1�D��r�:4�Myp�
���^����'�����W�؃{i��s9�W�7���t���{\M&&���j�?�p�%��ᑑ��������]�z��)$����O���C�E{���o����[s'�0��Ͷ��m��l9�ϖЁ�(},�,k&��ϥ�wZ�;��s�XL� Ӫ�.ׅ4#:�6���k�of�}H*rGϼKm��M�5bM���Yvx��k�Z]���F�%��M�x�Ė:_*�~���_�I�W�/����ݓP����h|�-�B
��~)uT�b��b)g-+�*-��EQ�����O�"i��-N��[��o�K��k��"���s9��:�ef���,ڎ7Q,L.���17ռ	?NTc�l]�y���T6�������+���e���x��GSދ��wE4�xQ,�x[��|oI<����h"(i�_g�W��%�LB*0;�9BO|P��d�m�V��c7�����<������\�OY?���ub��n�����%.vl�����2�49 2fĊV�$	�
�V �.(�m6T�:��7�����%����A��106Z��{C�P0��8G�{��D���������a�s1h�����Pr$]|T���3_-����p�W���1�M��4,�hEIq�����7uKj��EЈ
o�?�O#}���4�j��q�RZ����\~&���9��9�].�>�մøF����֮`2_�N�*S����7��y�6�Ț6C�C���x�����H��4�MR���\_@�Y/�K�M4ė�c�X
���/l6��FsO�Ì�:{��Y�F}���N�#����&��	-q6ˀ��t��9l���q�u������{��yGi�^.�u�����3Н�[�/7F�8[�(a�t�@8�@ۣ�FV݆z3�C���XL�������T�JQ���dw`�l����|i��6 t��~���|E�-�����:�iE�@2����Ҷ�3ۋfz�s����o�R�#�l�t�y�#���jV+{�wCh*h�0��0n#�M���h�"P�Э���� z��D��� ��?�dGn��Aa�$3�=��ѓ4Ibgdc�
y��P�!��V�x��{�b�%y]g~���@4��{=A7FDZKn�_<��2�P��[�KYۤAI�9)�B���s����t(�'�{�?��z����[!�4�?�1���Uۿw!���ʣ|�	; ���]~�cz[+�$��/U��Qaپ8x'�t��_2���-m(䕟�����́��e�]&�&������7�g���� _)�^R4[������E�L���� ]��?z��)e �qD˧&�M�3E�v�.d����C˻�Z RT��)1!h��FkOS�[�N}���
���;�&؄O䛉&�V
 =E��4���"$��L//uq}�J�cE��9q.fB��Ll�Ujǌrn�"Y��%��K�`�����<!m��ϊº"h�Q�7C�~k�Pj�?���Ŕ�X���)�>��B{Pg�R����ЍV���J{�$pa|��(�1m�����z�7!h��y�w�~D� v�T��Mɯ���(z̚pb�z}����h����#k9�&��bʙ�w�:��� ����5i
��(%[�����Q��*w*b^CX{?/n�k_��[��K�dR�����[J�:@�
�8��<�7�����I��qK�����t����L\�U���_m��[^W���
p�$c�	���Q��v��Z�݊�i�K���p��ƶ��UU�iZ����.�VZ�=�p>6У�;x����ד��S�{���W��JWN:�L<�<��7o����R���>�ɪ��OE��ĺ0l�ً��*W���f+�zW�H��dL �Z؄���D�ڛ��!���rL9r�)�dy�y�g��Z�mf7}:a�.�+Y/�0��ǓT��Pl,T��,K+8[�� ���2y�.,	�����0<���TՐ"���!���fd���nA���>�e�/�^F6�@�aD!��W��z��D'�֢F���4}���s�F`���JA�c�\��?�rt��rX�GV���i<[��ǫ^��V���&.3���>�9ܲ�<�k\݂JAF&	�\�쮒��cg��/X<�Ԩ�N������(1KM0�%�:�tL��z�z��`�����S��L�O�خ�����Zm��#;o>�,	�K
G��}0`R�hf��"�4Q4���̱��w�i�JQΎ��Rv+x�a�lf����_݃�%c�P��O�l�<�k�1H[[n~���:��������o݃�r��N�����KQW�B��p�����ΰNSʃ�Th����!�v��˘��+~�DPM��g��z��� 7��t�6'{�G�&�{	8��>�	��f�C)���U�i^���[�!�0HJh��o��ܥe���|�VY��:斌�<Rk��rM��g��P���.��!���}���>9�TL� 5!�z���넚�����#�A9�� ��ipE�:p�A��6\n�\�|�;�}����U!�px4���,4�[��MO���/�R�
0MH�S�~��� 5�s<��(�݅�Jy:�@�N����&�L+*��7�C�͸97w�L�ez-�8�1V6��6����f��z��5��Ƹ�������'� ��ACsY�a��]�aͯa�L�\-^(�FNI4?D�_���(s#W8���2t��e��K��0��@^tZ�>���=l���s0��ħ=��cNu��-xO��E�S�SM߷��^7a#�@�h;�z�L)��F�%��B5DG]��k��V+6���ߟ�(��i-w�[4<{W�B>���f�Ȯ>ݿ��I�� Q�#�?fCԯ]�=����ǟ��Q(��3�m�cJ�x�+G���2f����ծ��&�Ĕ~r��d>��Wp�1;9�gO<%�͈&7�}]"a��ݴ*�S������\#�Y�+R�ϟ���UMW��An�c2U�/aLvݼ��RGoL���:���\c�zq3t=7�`��iN��rِ��s��JKT[���r1���3�M�m��cYJ�AU��,{�aW��iթ���w�"H�O�Ȍ�
:兇B�|`�U��K1/K	�,~0$m/α1lv��T�PۍA���;����;�u�������_�9��)�B)C�n 	���%![��k��1��s��Q�@�DR�����]7��Kp����(L<�m���۴]D�X���	�E���c5��1E�&u֚������	���˦����zӺ�z]H�ͭ�����V����ds��������]RX����fr���"<�i�%F���yz��5$)�q�4����|e.��<��WVB��ͣ��$iHz�B=!�O'�B ���{J�t�c���\iO{��ě˗���]�	q�ټ�����8�`�;�t�5��W5S�e⶟��\����R�H�ݾ������N2t�_e��e>I������ck_��Dcj4������.R;����A2�_3�-�W��a��&��ԇ
�O.t�*`#����0��Y	��+�R���ms\p�T���}�������]s ���Оc^b8�Q{�i��>{��>Xp�U˥ht)��GHʗAs8�����PM���	���蕠�a��hG�)A��,y�{�q��w@��S �𞒗N���"�w
(���%gJ��V)P�;i�\g�"xC��.C����[�6������K��\���q@մ�%9�2�k�y���i���8XW�Zl�Rm��9ё;.:�|�I��>��W}��=��_�
�~���Iٯʰg}�u�`ۖ����3�̫&d��N%¶gF:��`���׿�K�B�ݿx�'B����/%���Fz���A��vY�ۆ.��:	��J�n�	�;�ˣ�rZ~�j"8�O�*`	;g���X$��s�����wS���c�O�W��J��N_�KK�CK��Ds�TS�!��^DxL�螌�z�Ty����s�!}R��������f��լQ:tc�S|��)e�45�e�\�^�i_#y�n� ��e(\�y��,�.R~�(�H�-���˲D�K�Lm.�!iP���B�׭�O�ڱ�Z�h������ה1���軅����������[v�U�BX�, 1��y��<sl�Y���v�I�ʟ¤�7e_�&~7�Vb��bF�ش6���������Ĵ�qO��j�@$��:B"28�c��NϖoJ�>)�u���o9.�8�q? ��������o�Hg�E���f�bŨp��oY��֓GT��dCƱ��Id����V�4�+����Az
9�ZMz�$f��laLY� ��犉��bnO*�F�:wA�"I�gF�$��g�!M*��'���mOL��j�BM��	V��Ǘ�.�y3��-��o�R)k���,��2��m�s�3���+ݑ�uj\�v��	I�{Y��L��� W�f�AL �"���CWf���gk���♾
<�G�i¯�i�G�ԧ~5+�^���\KKqa
�Z��^C��z���5M#=~q�8���Р3f+��Of;��t����(OZv�ܥ��(���5d?��-���VP얘�eF�N[���n���"�t�vY��߉�W!������eH�o"0H���.����XMR�(A�iC��Y,��ؐ��p�;�$��a�!c�.�#!t�&� O�lר�C� �]��:k�D�aR�Z��.��-�\FI�l�_�!I묨z�Y�~�˖R������Fʈ��(�=���pRaz��I�n�]���oG�n�9/��D��@�E~~C�cc�"�ѣ����;��^tSǆ���p��"}Ξ�B&-Ht�_������c'��=�m({�n�Qk�S��iٲ��}	J����7;�ꃄ!�	�taUh5a^1/��s��X�4�����i�Sz׼��~���U��_���)��E�$"),�����&(��S+�1Nq�Z�	fR]�>	o�	�,��
��m���p����Ge-�xD��ʖ�z.�ɱ%c��و��~�v�g0�d�0�`=�4S$�����LtT�N{��\��vk!���>�vOϣ�1��M����z��s��+u����en�Mn����sb���A��SX�MZPȏ��.�|*�����݆��q+�wa��M��}b͚	m��y��`I�]Z�/V�p��*�Y�i����V1�m��Fu2uѝ����yP٭Fn�>r��W�a�e��G���e2��
�^���2���Gc�kb��z�5/�o�¦i�~y�	���@�#4@�T)"Ԋz2i[FS#�؇��3���*��V�v�`��M�7Ԉ��)ڟ�6��W~eݢ��O��BY/;nCt��Xր����(�3���tb��^d����+-X��8��e5��e؏#ݸ7��m�c��S�����ŵ�5g�'&ģ���lV�%V����H�?>T���4�P�phoz )�)_eɕ���*_q�U���[<1W^_'U�tc+��=�GK�8E�-����ɆF��$W��%3_X�k��=����t~�����J���k�,؁N%��h~�.T^��A�e#ڳvu�i̔rz��-.p��X�-Y�㸿;3����X�\^��9Rз3��۽y��$�]�<�����K��@� [�&g��d��-`����O�x�}e=����i�YI'N�� �Ш])6��E^0=��� �M���+��C?�Y��ڕ�9�N��Ő�2�^V^4�����F�b�_?J$�3[���NYW�z���Ts,$?A���Y���{iy"�v/V^e�J
q��B��^�9M��lf*�סj�W�6�)��B���bN5,�)3��_�s�G��%n����/;�����U�s����`9��XAh}��H'�[_aTr�)o�b7��Bc����,R��5֚
�})�{�з+6k	�w���� 	A�!%z$T6�V� �eh�T��Ă	K���W�,�~��h�Qj}���l#�<�X�Z�oz �U\)�}k`��k�Eߊ�x���<5l��^���w����݂�5\1 ��d��"��P��Z��.ZM!)Zu�3�/��� ����=�H�e;p�pA݊�6�I�and�ۘb�l��0�|���uQ���>�><i���jl�p#GOjŴx%�.�|i2��Fa$	Φ��~���͚J�(�Dc2@*k���T�J&���i�7�=9�l����)q�<�˒&���~�W�JL�g��-��0s�5�I����Ū��t~ GI�qg/��GOR�}�~�������4r�GA�P���@�M�L�C�3]{���ov�!�r��X0�RYͫWӟ��:|��fC�9�<���]�sO����&:�,㏂�j�V�r^}F`1O| �N���_}'ӈ�oo�K�j�+#�Qvu��m2�PA$CSo;X��C��\j9�b��2��-�$�р�7��[z𭖂\�m��	��r:Wu"��/����T��ͷ���2�Q�A��5�y� ��!f�Z����_N��<m�?۬�k�h*��*~q.�ߐ�r�4��i�����H?�<�?%��".��B+�v��(==ȁFͥ۶�57*�9������F�Q䏀���>�U#͓��	�����ˇ
ZL�*u\|_QǛ$�}[I�;�^��u����I���	,Ѧv��U��= ^dzy������j\�{�;[���BQ�bGf��-jMr��#�ɩ9�X0�\���CҎ�1&1�{su�w~Sڝn�"�K^��P�.BBi�Z����0�΢ر?o�wc!�.��˹�H�Z���As ����qN��c1�o�<z��eql�y�H��`�΀q��+$D'��Ox���c޿jb!2��Y7�űA~����w��$a��T�蜹��~��_��ܦ�H!3?M�XB3&'�ЉkR��ӂ�޸�/l���~�Ӊ�}��.�sG�;�����Rh>n<�ٽ�ɩ��aJ}Ido��B� ��W��������[��g����3T�����@���(Í��# j+�����a9�S��6��հ	�msu��ίiV����A�c�}؞8��-:v�ǍiК�yNǂ��9x��`l�$l�`Y"�1��*Sڠ����,rb8%�YXv3=)�� "�P������ ��<����y:�5�w6C�!;F���7��̖�F{��CML�������ȽLTNIc'����`��D)d�]�Q�C����#�.2�*�"�����6�B����d%�(|�XiFU9��8���|��u�a�:��>AM�:�xI<���ZNc��!@����6�c������-Mg�k1�ⵊћRFP2���mD��F&Ɵ:�9#$��1#p'�m�啦��ޮO(���贆�*�Dj��\z̨p�<�v�^%�4�9D>hE�5c:�5�
��2�K����c��W�p�.���-�Y	\1G���7o��aid��[�J{�OǓ]u�d[,il���IW��Vc�ؕ�H��]�ܵ���ї�d3�d<j��j!�:���}�޻}ʂ*8՛�v�B�0#M��c�����v�� �c��W*�W-,CVȍ��?��8�ZX�N�����5�-�o��6��uG�Y�Ek�lC�`��:��qF\��_�����#���e}_Gy�6K��
g�]�I{�ڂN���`;�-�?�>��8�G�@KqQ9[Z�Q)ۈ��� ,7o��Sԙ�8)*G�;b=E+�c�?�G/=���0����f0fl�)��HT6q�z�-���g�mh�	��||�� (�6ra�K�������Y�u�`"Jx:�� '��Y�jU2�w���{Ov��i~FRƈ���_���~u;7ڧ�,ѫM�4�+��
�'�F9��1��O��H�᠐k��(��8y>�I�뤆|�FW�%� �{�8u��1�k�V�ۢ�c�IV8��	v3�����0�c2�����E���x�D ��{�p��z��uJ��3�_�ߨ��-*�A)LUv����_|���]�n
��~��DXXͲ��ᚃ�s	�
���%[����i<C��e��jI�>���቎ZPdq���(�֠�[��=C��i�2�����w�����3�v+
���S.jp���j�$�d�k�3K�(���-�A��-�����+��C*N�/9|;#)�.�hm����"��>u�c��2�p��T��Ӳ����Up7Yb���_�|��{�(e%�H�F�ڌl��Ɗ�I���B��ʿ���텺�H�7��^�뿭&�o�g>ݰP��dS(m�s��)ুtţ��4�gU3ݸ�82�z��j�v���i��U?I΁�dl��if#��=f�$8�ͽ.EO$�.e�'��H�N���潫*����6�6q��:q"���٭r)6\FG�
{}<�S��~Į��LÆ�/q��~�j�}�q'���H�FK���3�%T��2q�f7ƒ���I����ע�hbl�:1�X�l��J�ҚrEx�S�̿�gv99'�?7=�"�4�\"9��|&���;��t��`�\�8�t�\'S����?ݯ��$N���{�uЖ��
�ܪG�?�]�%�p��>�l5�1����AoUW���R�U��IN������ 7�mN<��]�b�iƀ���y�����]4^�c,��`z��N�>^� �;���.5w��z�M`?C�G)e�[y��Tե�u]�y�k�3�`��s��u8��X��<z��\���WU����a�O�l�YH_gD��3�$q@S��a�p(oO��MԚ\�$�9%��|�Y��;�W��sh��	}1%?�j+2-��5Z�n3��E#,c:���DW�4��o�XI ^m���ك�ѫ�#�3x��Kas�%i����Y�9NR�b����"ũ�1Fe�	6xv���O�+��7�j�$Ԙk3x�W�0��{|�p���M�4FFi�o�R��'R��}�ɍf
�w�����:,
�p�ψHO=E�?�����F�`n�>�Y�i㩒"�Ȱ� 3�Zgvk��Iì�0Ցi�HA�~��rȨT!�"5���00��V�^��d\��}�R�zMe�U��F>5'�����)�a���!�p>?�|��T��Zz�uS8�K����N�W�3B�Og]h��y@� �R`���_�ք5<�����C�eT�Kx+=��S�11>0h���M�B2!��mT�s�B�B�"1��p\��G���9���S%?:�8�x��+<>�P�,�ѪJz\�"6�aQ�t[��Ä���t��Vd,��{	�5�!=M���D�9�}A�<��B�L�s��" ��DXb�>��X�^�F�����fʱ�.y��O��A��u3t�r��
4�3G������_�u'����Y���P|A8�#}A��&947�o�|��DFN��j���	�������:�,�4!��L='=�]s�7Mֲ�u��OU��P}�tu�>�z����*}g�s���ޔ��(���^�+d� �a�o��,�Kl���>��p���W�! ��]C)�IL#�/�1s�>񆈲y[�3�K���61��i���<���hݡ����"���@tz�Df��N���F&o�w��dw2 $�Y��uf�w�����ZO�:3������@p:�x�� ���_��:��6���_'�� �NR�t:�$C�P�M�G��8@.J��'�fg��x��2臅h�����)���!R� P���-���t�xb��~օ�+W�PԢYR��Ɖ���ݱ��n����ڲ�żH=��N�5�6�Aj�2L��� S�;ua��N ��)�����Q�i+օN׈�o�Vme}��Ca>$w[Z�����1Q�wF	W����/���h�.J�˪X^��1�}?n����r�f�B�v�|�m}Hڄm�j4X���,T��wS$������CE�ol��4�`��bX����v��_�V�0o9(�����L��ҽ�U����P��e�wx�tK��7bꟶ�B
�Ų�9�fН���E�2�����s��`|��j� �DF�)'$.KI���-k�)c�S����b �F��Qp¤��ln�4i�m�da�ƨ/j�<���鍈�k���2���~h���\}�S��*��W�T������+i��B	�V�6BiMJ��R|�9b�$�Yx�'J�� �V4 �:���HL�z\J޶Q�miX��*�ю�&m�I?�:��3�ї U�Fj~�4%&�fvxvv�jɜLV���5z�*.�%���_
�
�Z�p�~�0
x�nϸ��cg}�A��Y��c�F��ew�tD���VZHw:��������;:��	!n$l��jA��i�h�i ����Н<��a����<J@Ź>�3T6H4��1e�J�{~���D��U���0X|Iw`�U
�ޝ��<]���w%�R�U1-^�?��Q����̚zЉ�lؤU�#��]��%��8�!�X��s�ꑉ������Z�lLu�1�?���?U �CW�����=y��>����Lo�S�⸿�iMW�g�t�QH| �F,�d@���'cBt�p��,nj�X�������w�k����|�O�a.�[Ⱥ��������y7�s�Ϩ������z&��f�&����NO
-���k����QG���0w���j�)��~�H�������I=�ާ��Ϛ������O��f�Z2K�CE7l�-�M��4���
�ˑ��T$�!_LJWJҡߚ�=���:��������߁p�p�Ax�+�\P����41�����X_�P�R��f��G����u�kYY���a�;�eR24{���� 0�{�i��֏.Sk�coD�RE2@rx(N�3�\Gvyi����/�sg,�y	�.P�����S��ts�6S n��ck�=���: \V�o1�u�ec(��P�����m�[[sK��h�n[�j	�H��Z��~&UZe���'�y�Lo�����͡����Eˬp�F&�F�|�mo�,�~�٢�+�Dy�c�Y��q5�o+�����^#�(���\'t�X���a�N��"F3��ҶBڒ�|7��j[O���Z��l�@5�!��k���l$?RD�&�N%	�$�|��J0�0�/^�~�[���ִ9��x	�?l��X-�]��M����:�:#̰�E]O)Ѭ,���s�G�͂�r�lyn��=���U�-}�4�Bn���m�;�zU	��g�L��l�c5����*����k̮��zwz:��9*&�D8��\T,��	y�dc(l��I�E"�j?��P��2���ڙk��~��i�хt
�Rq>�L�RG��M����3�V2��S���~�X��Hsn"|�hW�T�(�T���5�C�+?)NT���ū�x�Lv�#��U����I�l�l��Nv�ޗl��{���w����%,����0�	)X�t�f�Vac<*��
�$*L'ϰ�G$���	.�Jc�װ����^I�ϴ'7�'5B/��3ǽ4X��/�t����'�/x�oJ�L��U��Ϊ> ���i�ٙ����=-�P^2*��Cu��|��	�O@��&R�ܐb�+V�i��e���Y�(5�?�m_w�*#�״���>���tI��&����$eRV���m����)"6��B�sO��>����Θ��sEL$����ŝ�pb*�g(m'�r�w�,���FѼ���9���?�I������<�������~Z�@ew9VS�� �6�J�Q����39X��'�a*�ֵ�:�ρ^伅�7��~_��W�CM�	��i���Ӡ�ji��F���&�)��7чo6���nw���+��tm��٨���!]�+��qT�	���ؓ�v�w�*�Ec�`u���^|0�TP�DkeRnԳBA�<�+0qM���@b�_ ��n9$���lfm:�7��:(�8�·t������h.�d<:U��i�6K~�G�p� ��&N��'.n�L/DU�W%�~c*�w���c�^��{��lIy�UgI�����D+��}�^���:�Cn4^]u�����ϯ�e�7h��CK��\���LdV����
{�y}�vnD���>�)!��L��!���/'_� ����f0�����l�<NUT�Fk/��I�>�3ȯ3�%�R�����v�|�g[��cY�H��zKC�Gգ���[����RGR*�|$�['4N\z;U�ƳU�.|	�t7�2���bly4���Ò�ƻ{�2��Ɠ%k<cC�I`�JU��?��	�tg�A��@�Ʌ�Y/�RX�'' 4d�̺���z�V��;�+
�ݪE�4 �k{_Et��Z����(9u.4q�,�#H2bi�o_i���d�g(޴�F�ܣ�p43�X%ča�Q^wP�ck��Ī�R|����02�ޔ�,[�C�֫U���{r����o�V5�8���K�j@l�m�5���V�Cv��E9K�Y�1"��f/'Ĺy¤ �v�m�c�I����6�*�5�DH�^�$�DR�M6]6�����B����M">�@a7�n��^_�b��JU ��cY<,��o���'��ǁ�__P�$ԙ��n��SV��-�`S�3NqY����|�e1`���~2La<Z�3!o�{��u�0B��o�ͽ�Y�y0�/�Q��8�{w�m0>b�b	���P����ؒo�T��di��;-k��K���M�j���v=���r�;k��	o#�d*���+ܸ�G���~��@�o}����(�B�k�o�,����nz�Z�/{\S֙T
I����Nhx�,��R�H�h���u�{bF�^r�����Z��>Ro@7��b�k��T��T8B�����2�[���F|?�S�eꤠ��㽡�TP�E�i��&�2EͰK"G�'�\�ІЩX�Jz�n����D��y��)�(9*�(�>{%T�*�<���i4���ZC=[�\"�׆�����M{�įG��Ξ�� A�"�\����dt��l����<pF�7d������O_.��.˨��m��|n��}�Zɐ��3��"�/��n�B��P]e�tN@�Ԉ�:y%G�/~��:��}��(�p��l{|` i.ēןQðd;����H����fE/�z �S�M�n���O�h;4�N������둌GX����vא��	����,�BY2��ݘ+�ú��?�_K���.i���U��#��6c�5�R���3�{A�|���|���+�b���m�A���*p1dE��jn��|l 7���-�-�5�x�:��v�wƔ�+�e�`��i>�/+����&m�4cѠ��4d֍�0�6"�Qv����S�%����%T�MM��mW�Q��(���7�Y�Q$�B~�B#�� �l�W����Oc���{�l?�R����j���~�8��[%qKW��VG�0̽Šr�E_�����@7Z9�я�����@����}�S��T��چ �܉>gvU��i�})�DҌ��f˾J��N�H��N7�������հ�Ϲy�����)����XYE�~Q���"a���(d!]�GfQ���.���,Ty�e7����B�η�[�d�Q�(3�T K�9]�{ն֯77�0���Kj��/�dj�$`{AGzc�®�Rn���YN."/��R.5G]�ŉ��-l�i`�]����:Ր��#$O���*�\`5�tm�^d��lv#���}�9���\���n��M�_DS�x^ �L�����G��=��t�f�0���Jk�y����+�d���)�W^�H�l ��`$���hY|��p���k�c���o�h�oO��P��ܸ�WZ���f�?P�vo�7c�Ŗ$E�l�u�7�'Z���KEy��i��l�çc��g�����ul�T�l�:_���b�>�0!�4x��GbU�0,��l"�_�w�	�3`V��C
�ܗÏ򑻋u���E�됰2WF盏Ϝ`ݘ[�W�������bD�kR�Q?�N�xU���g.�Ӆ#��g��gJ�]e&�
)ν�a2�8�	~�������>�;p��d)f�$���Ik�ǵAER�J�[0�T�D��Y��R�b=5�c h�5w*�vs�d�tǹ�9"W���;:M��V��/�H�p�v.��8�1C��2����%��f ��$;�6]x�<4LI�t�q���p�-�.݅�(>�����7��]��m#�_ي��=�k��|�96�_��@�xS�fП� � v`Ǥ@3!���s�vi.7=�����>_���Ϛ���",����~,�;~V|���X�	���ʟ����yYM��1�r�&Fu���\1o�E�v��
w�|�D:��
`������Z׫C[��篳�������q~���Db��Ɋ�������7YB�H@�����������w���������m��e�I-62H��r�
�yq�Ied�$ȩ0=��A�v�.�67�d3!z���ZX������|�e��.[t�V0�⳻L��1��w��x3�ȡ�oT(��6�p�`�G�FV��C����>�i7w���f���G������M�?�83�.�'T�h]�n�������O���#Iw"'Ȳ�"Ty=⥑3��r���R;��M�zƇn	�/ذ��!�u׊��I>;�~Y�3��کH�5u���b�Y�;c��|�m���w�Wþ_�hJRY冞Iuy��?!�Y�Z
B>z�ّ\.�@��zq���%�f͈vrr�e�1�[L���J�+��;��"
��y�H#f���!k����SDY�|�9��h�e�������Tdڨ'1.�$<=)a5�:
g�pl�b�eLY�Y��w���r����Э���>ȃ�IC��&f,�ۨ�C���K:
������t���/���q"�r�3,�Pq�C��ˍ�b{�+��g%MO2�#m�S� �����7ܝB
�j�L�����ˎ�������ف���H�&b~���x'��tw���ͧGk�h�.8�]6U�)�!	\������kg�6�l�0���周��3@���3f����n��7G��U���?�p���t[x��Dhp�S;�2頞Ɂ���'��0#�"�"�����Sj揆�>N:��J��w=�,]&����[倈c�4/&�\��o�|z��Ì�f�{�{��$	�k6r3��4��&�PG�h����)���(`�46�O�ѵ���A_x<�1E�2���x�BP3��v����#d0Px8��,A�<��
4�|l�ig��Z_�R��7�K���
N�-��ר���g�z�!F)zĄp&=E`uA�0���z�=�^�O�O���%���ۚ�\�{F����Q����.m~�O?"n���*t6/�"ȥ�8�bl��K��
�~2��EP:�Z���+��������Z�_Df�@���Ԏ�Z1�g����:�xƧ�m��!�֫>Q��@Ϲ�?T~��U\H��h�C��ЋWU�"�� *�(Nn �>��L�#A\�)e�3�pI�k�]�3TLꐈ�����1=�'�q����� .߁iuZ7h*��#<�\_�|$��ݟr�C����;\������#[��f�Ҹ[L[����Y%l$zW����Qlb`��:|9�L���$����h�o,=�㪊:%[���v��}���M��lŜ����aB�\hJ{��f���s�A���~#��b	S��x�J~zմ-$y��2�� ���!�C�
��Ze���_T0��5�H��+��ٙ�A�PuC5�t�����vR�Y󔠻.u��6=��+��.K�)s�C��U�TE4����@^g�U�xU~l ���zw��憤o'��2��ݾ��w�?����֖�0��@m��~(۷<'����Z��_Z������[� ���_'�&�������v�G\�
�4�u �?'�N�q1}L�BQ�C�lV�X�a3<�y�Jx�������/�T�j1�zB���K
�K��}e�.A���."���N�����,+8-�����\��Htg����yف ���-ɹxÐ�%Nv����uC�,�񪦬N(�I���c�u�:;6��HuE�Y�Y,&����kCt�w�p������ Nc+~��C]�P�#�bԭ�#K���xue*)b �yo����1�Y�	v��6
���59��>�?�le�BЩ,�{Һ%:�CT�%U��E#��3h����}�PoV�R�� �}�kO����h��3�~X,/Ӂ"7�T�B��@Boo��D�-��	�2���7~J&ڀ�.����(r@��$�@��!�D�QeyL�T�;�P�X��9���x�e'C�Ңh�!�>��e^a���|O�7��X��[?��]����3}[��a	{]�`��Ny?/���DIg��zr�8���YEm��x�s��.�~J�:ɗ���#Z����L��>���j��4WQ���]M��5!j�b2#�3�!���� ��.g�C�LEb�$ �����8�ag���s��K��F�=OiwJ\A�苒�� ��>>�^���D�\zMH9�*w�������ޫbϵ-a�5����Y%��,��f<��D\�?�ܙF:�	w�j�����`���3�>`bv��XGe��؈`�Xv��f[elӘ�N�jv���������]�>65Y�L�+p�0�p�`1v?ƗPԓ��]d��}'PdO�`W鮢�J$�)]��Vʱg�m�5A3gk�K&g;P��]\Jw�ó�#��	��Cg{M�a���O=�ʟc`6x.[/V���$7�<P�����.�v@Q��vw'W�S� <��IZdꇼ��Tj@	��)�)�̄R�R0��A��{dS�!�x�xP��Į�󕫜H�� Q����^�D� v��eB���M��?Gx�ɨ1��8S&�X�n��y��p0%�q����ߛ�52i�AK��I��&�sJ������ęO��'�p� ��S�2 ��m��g���<�=�$�
|V��/ػ�jӦ=6�����.��0ߌ���:��p��U0b�6ar{�#�dYb���Ы��0˟}��.!D���1�s��������$�A�������ls9�w*z�L������<��9l"��M�*��O�������d������Dn�f%�:;~��ť?��S�����ԋ�i���'�\K
�(���@�#1���A�s#-�.9����$��\���^��@'^y�ukdV��l=����FEMs#��6���шd���"�{�BQ3oEd<h��85X% c���d80�hNE4v�u_5� Yp�������k��:U�aɂ�|�)��ȏ���O���:�_b�s�H��LR"�:.�x�bbH��L��P�[s0Zq�ɸ�Ɓ� b�a&�*�Uo��e�F��q����ӝ.�W�*��Z.h��77Y��Ҳ�C�ڞm�ქ=�_集�W��֣8 �6�]��X��%� x���\�#�%��ۯ�@L0;q��+�$�숿�8UCn��[�r�av�B�ۏ�؏J@	�O�TSw.�� �h��1��!g�@yV
x��6����v�$�r�rE)=���,F �<
`aتWu���o�s��QQ�ҥo��D?�%b��+���m��޿.��}HPl��,��p0�؞�$�6���6%
�%BU9ז��=+95��P���0V/�𐈤U��|N��(�&�!ѽzl�ތb�/!:�0���,jx�hI��>xFP���1���f�Sm�ݠ��i6w�6�}Sτm*���7�Ə��m��'�p���������+�6i�z>;n&3��=&��ϕ�9�-�,�r	��E���3�ČM������z��]����Jr�wM��|z�����(~4	L�?�wt�Z���&�~ <9��-`;H���B�B��i��0���]�6\r<,��&�izuv��[�����|ԓM��*[�;��J�ӆ'�ȡ��k�,W>%b
��kf�*r�`m�2u���)�1��h�t���O\�>�2CX-��t<N�-�j(�����ԾADUx�����-��J��P��[;���aL5�#�����YA~{q̢��4�Q=��"��1+r��l��N�V�����0�3_�(`��(*��@�ds�T�	�6��+a��yO5�v��<ϕ.�hX�۷�B-�b;��6��,���_��SEXѥ���ٽ�\���o�4�nޯ��]�Oۮ�h4��8癑���ǰ�H$`W6���	 �V�'r+���];_�J�,�V��%\m�v;��C�}g��V��|3Ɲ�O���&sv�=G�	��4�������*�b�jtI�'zC�鏑X��CnP��>fy��-]�^��Jauq����r��Fp�3�(Kjв�0����(�,��;?���?�&��.)Ev7nA�RQ2	�1��ZS�Ԧ� ?�T{o�@D~�:����KPw?3$]�n�����<�T��ш��	�\�v�C�u}〇jJ�`U|qo�x;%�D�X��OXaXY���7)O ��[��o���d��gr�X��:/<ך�A$�����ݑ�p���a��N�4_�ъs6�.�m��:�g�������V���*߷M1!("-�s��\�������ԬV�έ���1�UF=3`���+��i�+�X���Z����z{�ʵ=��L[d� 	8��BT�I���%?,��kibppiȠ6���3eR���"V��|Nmt�����M:����p���
�w+48xC�ְA�	¸F���}�,��)~g��:�����4��7k�U��+�]C�s��-`�L��@������tGЙ����\�.2��\^hpS�~d�1���x3��K����;-�2[<��id+l���=�F\=+ct|>���h��#�
���Z}x��j~�R�Ԫ��Y���[t	���e2= e ��  $�e���B>�w�iNa�����T�{IU�5��s	;�����$*`^�. �3O8͇E�WY�k4^j�;�|)�V�w�'2
�ؒ�f��O��Ja�����v�A������v^S�@'�3x�Z�wҶ��{���T4�x�B�3�I?������grˮ����5������ws��8*��͹y�[r%6JYj��� �+b�c��q��{.��.�-U4�r�������҆�-��" ��mKؿ?�-�V)h5����v^�����q�\W��c��|\�8ʞ�O��r�T�q��LOөl<�>��"3MX�̽�}�&����5{�� z}e�P@1蓼|Y4�Q�9<eļJ�aYP���%}	���n�)
(�~ӻ����JlY��z��w�i�(=L��~ij0T���;)�����1
@�(;��bAP#p�֙ơ�:~)ݧ_�o��;����BW�$��c�B���W�n��wͼJ웿�����x��А>4��`������О*���/?�쉅���ݠ���M�Y� ;JXlǒ囼�����ì	PiM7�5��b���?��fd��堘.F�87ee[0�N�~�Dȫ�B��1��\�oc4�Q��I��J����2r�~
�E5ǂqfV��5��l��+�$2�i5�¡���$Zн���`ΉA-�LJ[=Q���)�G��:�M�1өG5�hEG��|��	��ҍ��b1�t8��g������ML�UZ�Zu6C�>�5�9��G�a� ����-�A�mo�������=�z�����%9񎅪�����6;Z��m� �\:=���ω�K�����w(���˷�w~4I��㦃�w �B���QC��H���a}��gS��iR����
27���V)k�~����0�`��ӏE�H�,MyiM��$mT<�wT���m}Z�&��
*���`�#��=�@��kĎo3m���j.`��3�霜�=�@D҄�| α��FI�O�~��;��Gfpv30����Sα����s�D����X�IxxR���,������w�5vT}��%������<��3%7Sdv� ���TSs�q�ڻ�:;�GW��e�)|�6&�5����
��s�� ���=�A�"�s�E�GBv[L�0��׌~H�|����d]jڗ�"��O��0�#��-�偺7��xJ�d�3:�LP��K=����܋N���=��xa��b��dQM�T,��Z�>:^�7C��X� xʡ���#n�2��9lz\4��>�{8v���1����� �J��WD���f2T�I@M�jq��6`U-C?F۲�'��c�hҋ��
�Aw�R�R�aZ��a5qé�O���׾�<8��1���p��K����~��ҖF��y��s/��@Ek�	�`�o#�4�KP��J>|F���脄`��.)��n�2Gc������Sp8�q��>ጼ�r:�� ���}�������W�\�6���:����ڏ�@�`��N���,ǟ��N���g��S�La���E�c�SQ� u�����&x;:SƤH]ɪ1�b�sHb4�n�j �j�֍�xf������zB9d�l����m�4��%���}Ƈ�S������l��B"�%�)�DIdx[r�~ �� �wW��Y�4�A˄��j��%}Kˮ�93/��;���H�,\��'�e<��5F�me8�H�?OV��_�Q�*@X��Kx&7bP|�4g��lS�ə���p�l ,fV���`U�������|O�KU��-v�R�]�q�M��|�ݣ�4u}��g��A�V��'��
�R��'�a��7-Db�inm����ꅡ�u㫗�̣Q����ô��BH{p'�&���=þ���DF�k�]$�8�E9.���S�&�"��| 9�'~�'B1`��Ǉj��>�<�W*<?f��%߃'J��#H/KO��c`�P���=�}��ip�&U�/^A�^2���XlC Ӓ\Z�}�xA�wZ�����2�`@Rہ� _���yY��y_�ǆ
(�(N��������"��G��c9$��rٔ'|�������\�(p�Ψ�S-��`��Rv��MS�4�B~�ߝ�J���1���
o���od5�?�]$�Ս�Nf$/�kL Ȗ�
���4Jbh՗����-��|�nqz\�A��"�f*~ۍ!�mA��'�f���+J�R��{�u -6�XL�X���C�}�ʾQ�/I���h�B�b�c�ґbt��sm<{QY�W��L k<��yP��e!<�͏B��MJ�} �*`�?(%&?͸�ጟ���GN+�`0�
�R����:������!d���ȷB%V�\i�4���[i&���~�z��x����[άU�>J���I|y�����D?�7a��m	,�˨�]U��KE���W��[@��Qz:3�/[aE?�#�?��Z��N_Ԉ�F�k�R6fb"5%�>��Ľ��[0+�����1�[����O8��g�	T�]�x*-o�-6���L�)���ި7��Z�r �T�\��{�mC�f��Ql�a��
�*2���g��/n���~����Q��}���Ú���5*��J�.��'I�"VS�w/��(��@?����vpWS0�- ���ո�Ã��W��Q#օk������;I1�ghް�2ɩ���7�_P��_S�B��p�s��h��ؚ( �F|C�v��29`�-����}����8��&@�>��g�(L��HNLE���0q�a��L�3Φ̯�M��)�z�y3����i�#]����v�4F.����CMA����dK� e��;�B�	���9��^��߶Ã�o?�L��+85� ���I�/�m%B%d�6�aa�);�؝�UC)@j��(��`��U��.i��8��s�y�;Ӑb��7+c�!hO{��kC[��#Z(���Ob�\�L�i�9fH[�������:!��Cp(wz�c~ X�����|؈iI����� ȸC��
Fl�>8�f2��
%�d�֧	�k9��X������ĪW��򹏤1��&�]��I~'~8���6c��-&���ٟJ!� �x
#X0.�x-(v��1�L�k��5�܁E���ۣ��%�P>�
+ԌɷBJ�@؛	�$!�zXv�^
AMH��F�O(L��n�fMD`Օ'���?��Woi�����n��t�������B4�r��z�l�`0?�GM7�Z5�d�6���L9��B��7!'x��D�\|�>,�7]�oґ��Ul����2��*iɱ�G '�����q{��ߩ��*!3z9`�+�pPC��X�-]�i�DΩO��	��A�t|&zuHR=�������u�ܮ��XU��N ��{ҮZ�{O4�4) ���wpJ�x�����D���5��l�t֜��Z|'�	�՚�kx��6��y�]���zr��$��%[i�8��/�V�g㗱	L�y�,��Gn���B�mNn�(W�}��T��b��{m�ɒGZ�t)�������ߎj��I_�����?���@��wާ�� 9����1�[�[�5���d� �ֈ.+_���4�S�ǐ>�����х\s���د&i��+����.�R��b��!������/mY0��*L ���+��	�d�~>0�8�Y҆ƃ̉���Z��f)6�PS��x����x�yMt���,��8E��T�����Az59�7�LR�2+��4�A���Op Io7]����WV������|3[M�C!j�Fѧ#�!�*Nmv��FTn��\�,��5�Cɚ�`�������&=3�w:��h0�����̝���|щ��or�&�e�u�LB�ej�w����;7���'#C����8������g�4ᓾV�Ȫ���3Ra��
�kr��.�[r }��X:֨c���d�
].%���V����w�Jd�k8�l�����:M<)5?{��
艭c}-�"	ͪ���T.�E�A�"�|c췘|g�a�w���[+)�P�M��L
zS���V��؟ҝ��~-J2�_FBVx�ػ��7爚'�	~��3�q(���vX\�/C<,���&H���8�֣%!����*����9
��y�M�v�,y]�M�7檚��!sJ���=Cо�Щ��`��d�@S�S;
�'�D��e��B~^uԮ�]���s��QF�y�W!X8�$��_3!��[�T�Mɘ�*��&bK�V�ɲ�M�nnJY߾CċA�h��|8�V�Z�&b=�*�I�_#&��l�Q1�^|͉ⴄ�w�%�	:+. �&��H�e�/�X��Q����Ծ/(d���w��"�b�kV��&��\.�5c���:d �SI`�;C�iyV!�yK�	��D�c���זT�?Y�)-����6E�#�s�Q0}[�̚}r�����S�9��+��+�P��ts���=}�s�z�(4���ՍC! ���)޸���R��N��sq�;tm3����im�hגE-���f<��V.3�:��e�A�_S��:��h�����sg��U�D3Z����j�,J�W$� ��k�b����Ŀ���<g��~U�=]�[������I*���,8�D��̰�[-� ��'���4
1j�6�`�[�=��X��P�8��a�}��b:��}�l�]d*��|W1�z>�x����c(��2�A������8\8�xP׬n<q��a��>ٵ9��A�g8�te`n7�G��W�t�������S�V�E ��n?4?�Q��Oo���i�=>~+�u�-���9,Mr%X���j��<n�`�VN�T_��eaX٤��C�k������L/�ν4'������?:=~�:Ԝ�֍h�n|�5V_�Et4���|4q�PA��X�(ho�=�0ry��������BF�FE(�p��a?�OC/������4��Q�LQ^K�[��h����.��t�� g��=���
$�P�)�Y!}���0,k�X�9��76h�[PB���֠BA�4(����4�^��pA�(�n�7"��teK���U�o�=���&Q���T<CQ��w]��WSA4���U��������1i�k_�6#F6*���Og�ͪw�˃R�5�qP��x�&ݗ�QH!���7e*	�1��w.�.�`�a%�ڤ�qU��eeY		���8/w�]���W��	�e�[�� �,�FwhTN#�ʷ CE�����T�'���$ھmq��������c�|#o�>�#�j^���$H���I����"�#��f#t�4��w�!�Zv���L��i��Ǹ�{v�?ڶ��li��j1zΦZ�^a41��''���9���!47@���J�A݊l�}��GgV��f�H>�Z�:�A�!���\�5�9ɢ��E[��9�u��s�bH�������6�6�\��5�w�fK����\ܤx�����*��a l>!Js@Tx]35������,
�R��H�;�{�M�xo/	X6��}��2c�
��p0��o�eDJ���C����� ��N�Z��E�$���ޕ^=G�p3x��C1$=��/5��p�c��I���̍��#ZE7���%BѨ�45Fx��^s[S(gI�_{qH��JB���;Aq"Q;@M����F��ڝ�iя��|�c:L޻���������"��_M��o�mJ�0oLqc��
����R~�g�g�C���qjH"Te����V˹�Y"~��ڞ�������k\�����6VFE.���_y�Bg�2ar*��T_<�]���B�����"��{i�ޡ����Y�߃�������?�;N��:=n
���y��}7)g���m��ReNU�lX���Xr�	)��.s�Ǵ,ɷoo[���dMZ{�B�*kŔ����$ Y�v��[����oC�Rs��W!EI�����,�����_��1[Sv�#'�����d}�2|�vl�����c�&%�N�,,�tt�������
��"�p��U.�(�wƬ�	Y� p���&��'5a�ď볠�'f�V���������.��~��2Y��^K��,�N�m4o� %��D�Q>ĳG�\T��M.D�I�����F}�ה��e?`]t{���r���2	�si��E����\��\�o� � 2����s��~ͧ��5�"v�{���q�T�:0!����?1~�A�������J�D]1� `�] ���/���㚀���CZ�B��j��Ieb�9����L0��e�Eִ��&q��!�f=�<庯��#�0B)䭪�ɲ�Y��gflYe��.]U�R�p�WKޟ��^sgⱝ�ןez�Z�E5�6�&��Vk�'5ChO��7�h9E�I��eʫ�U�Z�ϖ�xޕ�Y4A&J�n�W�"�J�h2��an�W�U�ަ�({N����YgJB#Ll����k5c�e�5(hV ��r9;uY;�P��� p$w0��*�w��x���ׄ8���i���_"5���6{�]�]��u� ��l@E� }��k.`ЋK�(��F[Ңj��������2�Yxt�� X�k���M��Tu7���������|��iQC�g�L�O��ܛ3�*�.)��}��ƵOk��j2;n���V4奘� b�$��f��{�L<d������W�_��;@�4x��Z�m4��2/�y�TMNUw%�hcZ�#k� �U��,ܵJ��P�KD����B&c$��,&l�Mw�{�&x��2�tZR�O�צZ�&^�?��&�.�O�(��yNO`I��l�#�7S��k-z����B�o�v2��f���_Ge\��q���Y3����7l�uh
~<TOT�,z�Y�,����F�������R��Q��=_Cժ��3�	�L��ª"� ��� [���q�:�~�	����:#C4�0Tg��� �!9����ț�Y���@{��d h���u�g�$T<��.ۂ����}��3�25.�X���m���O�.�΢�����̆Z�u���3�����±��H_W��Aݾ�����u+;�AG���.��oAČ��ZUJ6����E�0�%�u�A��
l�� ��	ן�v_I:N���I�Zo�� �,WdM���1�z�d�8��۠s-|�Xg�0#�.�wS�$)BU��IT��"�Q�B�sB5u��c�z��e���K��HS�9z&m3��^�YÇAB���%�[d��Ck�:���udG�����܂Pō��%"�ܬ��̙�I!��^s�n��k�ٸ�<�d���8���j��fu�OO,�K��[O�an|1�<|��2?Mw/�c^
V���{��P������{o�39� շ{:aP��+<������ ��^�_�x�?�m����u��ڶIXd!]|�v�i3��Q��ve%:��<~�2��h���7TV���3�g5�J� �_�kA�w�K�H؊�&���R� �v�8+��jP��H����;� ��7��oDUS�⦿�i�Y���ɧ[�-�`4��7� G� ��|��ŴK~��C4�[�D���`
.�v�h��Ŷ�S$����˯�'¨0:��/m�?0�~8BCDB�B�=)e�B�s�.D3G�|��[������%��sO�~�F�Ӗ��p�1�2Y�#$98�p��O�J�X����kWȯ��<?��J�{�}@�t��o��'u��������!�><�M��i�JV��m�V����A�{{�8O͡���22����^$ T^�B69d[���-���Ĝh]o�Ɛ��2FL���(�����
v�ۛ���aȽJe�P�9:�i�i3�"�1h��PwmC(Q௭L�<;�P?l�/�~����?C�G��F���4�D��˯�e�q�cA�S7�CJMȂy��* ���V�O � 3y%�.N,���\U�{䁛�_%oM��vX�6�@cXl����o���v�6n��-�Mf��	�����,n8��ո��'��{�J���	��9ɢ�F���O��W�����8�)8�ܤ�_nxs�0�rV�%�^Eel�,�i��ua1ݍ�ˊ�B�H��ֻ���W�TNv3wr�@�?n�;/k4nw��ԍ�#؍!D��bb{����V���W	�g�5������l�ޯ�����8��4)�R۵�[��u�.�S�w��`iW�vq�>�$���VIp$�6:�`mWb�B�"O�wM�O����n�.<���8�9���է��A�bq��gC+�og��ш��B�`�u�E�:_߽��r������fU��2�H��>mEhq�	9�����BZ�^NH�$>�!C�D��?�;�g�7�> �^��Ș*��Z � �cͮ��7هiV)�i�emQ�Wo\�T(���\s��HpNm
�R�T�m���^�N�l�-�c�Q������<ʻ��|���������x{�����Қ~.��������2�����3�!����t��������F%�eB��96ſ���R�c����k�Sx��_����d��z�����%ө9.��*p(��G]��*�$_�?�m�m�4oZ�9���m���	��W 
X��rZ�T`�wr�#b-�cġr����k�v:�����'}/DT��Y��ͨO�9�P �s&�ydF�d�58�
q"-;:?R9;u������o���?�O?�sA���B�|B�	w�SM&�z/ͧ�+������hu�g�,���_��+��K��/�Y�@f<s�#g�p���+.��.�.\�i�;�Ŧ�B�	�8i��m��۔����q�����~k��jͧ�5�@��,���3ќ����Cڕ�2Xc�>&��M�����m�`�4Q���z
3�v]Q&[�k]ڡ�`C���k�į��cz�uP��&Q;�Uv�S���T�;��|?v�
�8�	e�����o�S�F	�F;�x����2ͱ� �>)�5�L��'Ҧ�>C�,��E�Wz����1W^{�q���y���Q[��]���7�it�!^�Y�K9?y�)��|�HNJ1>1�߼F`+(W-�r��^��CEb�y'�|��us� ��꤈}0�a�J�"���C��Q��}k�Ct�_��U�\�`�;v��U����NF�� ���É��UֵX����=y+�np<��Qң�����q�!V(	3`)�;��T<�&�Zz����b���]尪�>y��p�ܩ����PT\.�e��NM�e�Q5��t*���L���$ӿEP�8�l�9��xM)�����^14>���'2q��aiٕ���{���+�]�n��Ώ�{�{�h�J!~5�U֊�7
�Mf�x�}E��o"')
8���&�ː���)���N���+.H~��6Y'b�gnF�ܛ"b%�����=�����{S��3y�T�c%��������d2�`�mb��1���,f�e�h��·�[��(X�y6\܋�`sv�1|�&�~�1��UVn=�re�E��lT���}���=Q�_��)�Wv�[j
��,& �ǜ��J�7yXM�Nb��<�A��?lP��2�v0C��Q_�"e��@�"�EP;�z)W�7�U��<;�C�	���%��֩�r�J�V�@�(t�u�>��"ֿ�"_ ��n���5�v�G�\ک���a��푊�ո�/��_`��AU�AVge�@��8�#$|����V��W�� ����v�c:y\��ӼP��؜+x��J� ����?�&삠JQ���hצa	B��7OS��ΡwF�x����{��o $�B��"D��򇙻t@¦���n05<?�V>\כ��Gԗ�1��Rm	չbN��DL���t@I����q�V�O��":��\�FН1�?�M�i�o�ܛ�)e�ԒI����3,�f���3D�Y���z������Y+�%������;�v6tC�p罆�ŋ�г�X|�V�?Z�H$���B ����Z�En�t�1�?����k�:*��5Φ��~6�v3 �D'�R�� �B����yD�)�x��;Y6���E��M�M:��/���I�\�M��C�v}T��w�FA�G�8��?�˘�~��d��n�+G��ݗ��1�c3y-�PO{�(NhV�C�Ў���0�V��hl�V
6�QsA��Ao�B�y��T����~g�{ShDf&�u�����g7��da���x��v%T�Q���y�G���_���|�y��m�U�����N���7*�Rr�f�dm���O���Q5�W���oE_�=.����T=&��jh<�� �l4R�+���2)e�6�����pY�������7�e/d@����i.[/���.��A���k���}��� ���9ƴ�U�B��X&�ك�k˼ϑ�>�pM�1Bf��)�V�d�{��]S[L�|��j>��l���x��v��~��Ϛ���v�9�\7�Z�x��~�:��V�ɫ�ns|m����r�9������T���|:}�X��X�E'��b�0HIJ-�F�:o�Y�?f?�Lcc�}�'UǸ�<s��-f��id:[���?]p�~Vc� y�8n��
�Z��ڴt���?�Ғ�i�\1��ꭜR��s�P�����\�<��X���Q(��i�(�V3xXH�i 6��!�HQz��+������fo�!���/�r��pa�ɳ��G�q���x��*�4��5 
Q�/e��ng�\�N��ğ,jb��ӳF˶��8�s<ۻ�!d�=k��5�:!�d���K����S����[�3:o�\23L��k&e_��۟��aӤ%��5JzYd�J�B�J	Mdi!9�i�H��z��G'����/Bø��Ê�rṁb�r�m��x��F�H��ዐϞLF��$ �Jʗ��]m�Ĭ�-h��a�����R��93��w(+��B��Yz�O9|��"Ls_���VX����a�����+��\������R�U�8�����-�R,�������Y�*��eB}��Y�'����Y����wU�sane� �CO�c0��ܧ3}�'�$F0FI��n��]�]���l�J�'�|q g�t����B���_l~�����@>�_\��=�����p��
A�[*����N��*Kb�h�q_�DӾ�??*~���1|�Q7zMKd�'��^�Zt��+C��I�oJϗ˗w���T0�^c�o\�c����iL_�V���xT�@"C�7J� �Z d<݄w1�C�D�mWmxa2ll��f�,v���'6��ེJmzFj�{&�x�j�����1?!���)�����O�&/�;�N���� ��e�/s���8b��~�?u0��E'[��E�p�IK�g^iW<f	����F�<�I{�r)�Dn�����7��>��@>v���V]�_��2��}�M�p�=O&�!�?��P�뮳�� �>�D��Ĥ)������b5ѫ��F)ߧ7F�?s��I� �����Ҁ��7��5_p�ὥ!Ƕ!��j�f�}Q��.��h�+���8oMv�ͤ#[�(�Nh~F�{ܕL�P�s5n��`��]��(���8��M��PL�	B+�*K1>���4G�)J�笹'���D�j_Ǩ���}`Mѐk������|"r�Ö���3���n3�e�-iW�+V�������̳Η�W*?f��uV�{�7�-�\y�
n��'�m	Oȵ����Tc�� u��������A�#7�Of&qr�)R�&��o�Vy�� �}P���)n;�x2�cR�A�ـ��hZ%��O1Z��Ru�+I =��L�`��CC�qg%2I��x�G����&�˕:@�}�+���b2x��|��6Xq۳LH����E�A�6>B<n%���4
�rBl0�V�� ҂��,D����B��9`��"|֎q�k_��"�_�������RM�vͣ���U=�X��V<AB�����eS�G�����ǎ����A�L|�ܯ��%���-$0=$��4��e�"2 AuK�Vp�Ջ�9�>E�ͮ�m]��*�i_����wq��,���Q

���	.̤wNv��қH4�Vj�]�N���:M�;h�B�C,�8ޮ�/~�[A6���^�=��d������a>�V���
^���\�fb�q�0�8^�)�J>�|����X��Im�|g�U�pȎ7�O��Q�y��GB�����i��Jߓ��y���S4KZ��>h���:6'�_:٤?��M�%�kt�`�q�p��{ׯ{��e��q`�� 0�_���`
 O�����ɮU\�]����b�Ê�Pa�U��� �5׈��`����U�Ѿ�H�C�O���v���1Ec�	&��
�,���4E��{��LWݬ#(��tNGD�T恮�?-d���m��X &���#5������~��U
d�`���(�2�6ni���fm_��+�48��OA��nॶ��~��q:����Q���:�e{ǔ�3��4xA8�<� 7f�?*��M`�l
��B�X?I��T�e�BS=e�>�v�����i[��ٻ��	�2��W���{7�r�ڟC̴(�*+�~f����Y�+�3��b�kn�-Z��1�Tݪ����x�[?6߃;���9%\'FzeN�<rE��D$������z��B��e�ú�������zi
�L-�%-/pM�Ȑ�ᝀc<pl��b�͋븜3���9vUYR����Bg���(�k�i��B���"�M�r���%��
#��K�K�Jy�ˀ��������+Y(��!�~��㳂g�RV��U���.��v������p�ڻW9J�R�`�?�sk�>#�C{��u�.]	�ʠ?���yE�P�X֏>܎0�ď3k�%+�&7��*���;��y#p�]�>J�$�@Y���V��ic��.cyM	bZ?�����|8j@�]�'?�8}�� ����W��ic�����3�l�>b�;����0�(̴�a,WF��~!�ʸ���6JjX��G;�/������?zk"[����|T�6�D�����%7d�u<���_k#�v�����򕛔ѐ(3�;i�qߝC���~@�rN^�$����@L@m �\�X����-� *��4�;��l�$k|dY�s^����%��]1�M�j��m~��	B"���r�idtX�����h:�7��9��2P]�T�o섅��i�� �J6�
�1)���'R4��i�]�&^v��#��\1��Ճ�	~5(��#�.$��NG�T �y
�^U��h�dE��ƿ���t�B����Y��t#���㖿�<��%���R�)gCT򟄮((�8O �u^�H����޼=�_�ۼ�����]�i����a����b}�Gs����ܥUL�+E���5�WG�����T�<="�i坸��sf^�l���_����d��pY��o��c�/�YLQ��t�K�h�`��Ӄ��q�A�@�T�I#� b�x謣t
m���m�q�c���Y�
�~�Hl�+����C��C��1���4g��fPqp��~? �5�o6��*��`�M
��\F�&Zm�:��F��))�v]�c�4����OK2��f�D�<i'���Y����T��ʔ v�M�X
����O�_�U(N�}�k�b������k)�J�	��L��M%�`����,�:>���W�S�?���cb�~��1����"��%i}�<�J'_؜�RK�X"{��֡�X��繴�]����"��� j���;�������������#��,���# b����TU��D���A���������D4{]�0��$�����Krr���ut�����`[C��kVʘ��h��v�� �z�h�3W�U:���Ј�l�g��9�Du %]:07NFO ,��_�H/��s�휡4�=�{R��/�/����1)-���_�W�/Hr�S�'\Fsb�nZ�yd�ï��i[�X�7�	�S���a�l�k�<OQ1�2tZ��JDo���,�"��j+6�?�W���ՕM�z��5ǦsCV �@0P���`2�[��K >1��z eCg3E����svV�Ds�}�M@[W�k*��5�a�p	O�ɗj���
sp�E�R�v{��Q������N�Xkس�+�ڪ�?�"/��u?�c�<��J:2�?5�7��%*�S���+��$�2��d^��O�-�̮0$�QN.0���b�핰��S|��h�]���(�uy:fMZ*���AԀ����t{X��
�?�{�([��|8`� ��C4������E�Y	�|�d #|��̡sΐ<�W������^�?�ȉ��x\�7Ƕ��_89,f���7��Nu6�.`.9���~�Y� ��și��&У��'�A�4EP4�+�V�+|G����XN�&�v�"W�L؈�{ߕ�-�kWS5΍�z�SD!�KDuh!��Yl/?)�D���E!bd�u��4Oj���w��^O�`v�o�+�HaL�u]8y��n���\��k�(Z@^ �h~_+��I�x!&���#_���NSÅ�ˠL^W��H���k���*���ޡيݕu�h�k�<��Ф&
f$VMk����ɥ�|����%Й�s�V�=�_���b�?2���&&�`���~�~!;@�_�M��z�!�ɦÖ�o A���ڢo����]TR��5^���jLZ�"� %�$-x�!
/2%��F�բ8�L2�/y�9��*b�t��H��}�T�����1k.�ٸ�(�ȍ��g���G��.�3*r���䈦�S
�G�e�`�b<��C:okr���I1]j	���.`7�W/r�u�g=��O��v�a�^���Co?PM��~#K(�ǉ�<�+YO8z�yv��a:�"�hF�ϰ;���?|��.*oO���Bd��q/�����\I2E�#g6�N<��f=rG�����3*�>���CE@s�|f���6�ѲB *��A.п�c�K:�S-7�e�1F�[��-�;�L�T�<��A.E���u{˲ꝙN�𔛿>�w� ,4|�N�K�qH2�P!��å�Iy鬶�ϱ��9܎�1`�Q��"��[i|����u]s��r�sʉ�Bf�v�!�܂(�~��M�h����t���Ť�S���kz�#�5���~��h�sT;�7
K�6
��^%x��S3K<^̀�n��/xv���W�N�QǔB��8�������̠�Z�8Mm�f2����b*���ݘO�=���'>�0FY�!��b��l�;�#����$Y�$oJ��z�&5�k��~�p���5���w#�* s �uU-���|>,�$�	\��#�Ա�n��Is'0��8C�e��,p��e��hL��j��˯P��q���ȡD�X�(>E(����9����mH�J�!���y~�7�O���-Q7����Knm��:\��+V�#0���V�E�6b�i�F�l>�A�0a��$zm��圴��I�3�xu��}�?�jsmu]�9Q�r[���7c��ҧ2a�ł2h�T��0d�%�:����=�=���H�2/�C>�Zscf�,�]��i�QlHp��.���ܜR�����(�L%5�� �D�y6��򆺎)��+���|�I���e;q �(Q�ͣB�Ł	p��$r�Wupm��'o�w�!��t�H4�K�����}���7[)�-:�|��N�?瘥çR�Y������c�10E��@�{���L^ٌ���Y�Fxy��^\��&�i -���O6�,�WR�DL��v�D{��(.��ŭ#���|�_�����d�N� �8��1˪��l�"@R�֠���1�9�pX٩���¨
�@M��Ă ����5 m�1Uy�`�[��	�щH�p�����"����q�j���$��?��Iklˡu�5>���^�7�L���
���p�����3���gr���2yb:��O!Uq�i+��6�"0�E'@�I���<�׊����o�6�Pt�(Ar$2����K�����(�	yHF$�
;$j��3����0�w���-j.��Z�&g���]'W���kLo��V�Q�w���t`Y�"�¸ �ExA�cdEŀuڭ������6��$���U���?�U�uNM���A�\+�G�r�SZ.�Z�����j_�ޏ����X�6�a�u�I�6��{c�3X�&�%o���kR��x��4�}@�ɰ9�e��V���r��ϹT������(�w������gd��!�$�� �t~cLQ�t�Qf-���<��F�nYV�<�ϚKm1c�}L� T>��tE,��VKrv�����Yƭ9b�z�/|/$YZ�E�yd��7�Y���ތ;�t�ݓ������њ��V�/Y'nF�����Ҁf*�%i�	����0_�6�|U_hgB��`�BQ��(���S��Հ�"f�Q�f�հk;����kHd�PV�a�0l+��\lTu�֑1ke}~=�Ҩ���&��d0�j5�
�f��{0��ؑ�nCY�E	���g��S�����9CO��r��m���V�b���3�\�F%ǽ�s]V�(��п1�X��ֻRp�
���kD>��i���$�(TL�j����[����g��C��Lã��:�]iF$D�C{�q�w'4��	����Y'Ib�g�_��n��P,Q(����A>qEu�JA���tQz��X��Ժn�,���_G0\��� ?�-��ў*VI�߄����ݞ����1�G���;y�d����}�[��BGz]sɛh"/Y*���/�-�l�h7���P�R1GI�ј�QwI+k��]:N��kp2�1���J��,���o�\ 	:�pb��ٲ��o��c��$�?�����B����~��ƒWL�'��-�*3� ���B��J���9$�2�DJ%X`A��jO��@�%�뱧ن'�B�/��{>i(�)��qC���_{�Uo՝�"pH�Ҁ�:W����Sx]J&}�F�Ѫ4ϕ,���?OGn�X��o�s�����=�aϺ����p����+Ȯ��}�� :�>�EP$]\����n�ʮ��{D�9���웱���շn�Մ�F&{���+l���6�W�r��T��5�0�&�Xf�.����=T��F���
�M��U��bw`C�-�+ `mX��������$ÿ�� ����dن��}��kOy���/�\��ս��KP�c�O��2���U�p���)�@5�M�>��;.+���#���">R����Z�-��u��/5 [v�篑NPy;�����iI�"�\�!7�sA�Jt���^�3��BNˇ�U��g!6���Zha�}�*y��S���.��G}]q�	��� �oY��s��C��Ԇ������1�]2G�e!)�7yN��ͱ�� _ k8JR����;i,wV�'�����^5�mE��ݲ:���6���w��
dVOJ�d���ڻԞv�Ԕ�0�nA�����4Q�����v��9T7;��*�1�W���Z�,�='��)��-$���~io�{j���.�r]����������2�u�1���󤭇��c �HF3���;�/b/�DNT�g���C�M�;�x�(���;�b�A�}*�A���f������z Mz;�L�����Q�� :
��\�53 ���k�&F����O<�FG���$S&�x�6�\�qj�ul��,�^c���^�+I�gKP�`�������q�n��ʀ=�Z٢Z7�K�����1Q.K$k)��wY;p��li�[!�+9�[ _�j��e3|������x7�
�7w,����
�1M1���*A�8I���&r	i�k��~qZ��o*����!����#��N{�ܩ.�:�͸����RЍ����t��u��Kx� 8D< �짂��vc��kUG� �Y�`�Ʀ�kn���F�UD���PѤ��l�q��X[&x�ek���!yЦ\��ob�Q��Vp;vT:�QCU�:o�;�Uٓ����<'پ Vf�G�eN�`[����R�fQ<ōr���4�[c�^�'0��M�?�_x��i�[��Qg�����>.�P=ǣ��Dk�r�g\g��(C/����q�*��x �..�/(}�'��#��fe\�b�Dr[~��J"1q�'6HU�0C|>��1��C���J�9� .���G������S�ծ�����Sṍ��ʎIبT�!��������| s��!�w��7��{Y�O�oC�N�L0#�Ő��� /xM�֗9bQEQ�yj9J��yD52Y2����j�3��Gk�
�Gzz���T�>B�/h-������L3���t��RN�Oy�f��C�*�o�I-��
��a���<m���!#���������@֓��6.L���>E������2���o���?��nA@� KB�%`QaX�)���X��#��&���4�h� ����^�a�m����Q�����Rk+h��Z�P;bۊ��y{Q��,����E��/#:4���ip������(�ڣ٦
ߍ�ܧA�		��04�Z Ưb��$�y0F��:�:�E�t�#�5��)l1^BW"L�5+��u%���[�Q[}%�o�|�s)�E���ƮJ�3������e���EX�w���|錽������	*���@c��ѼkM�C�����?L(/�"�DF��@#����x��%�6��������ʸ������\D��~g�{�:�M!�s�)my�}C΋�(`i�~�Ǎ�o�m�����]�n�U^L�{�Nt��;�aֻ��ј�(l�C��+�������/"�EV���a�j,"���]_5����RqVC�e��G�#���՞z4抾^��
)&�(�����y���͛&���\ǟW&7�Y����[��Ow\������-M��cr�C���p tA��(,yr��ί���,Qa��Evj�a�+U{a�g�}�T�Y8��u��߀*�h�{D�!N����a����=!QI����/����{^1J����zi�jjk]��\o�t�1��uʥ��>�ٳ���/Uek&�6��რ�F���(4������:��oL�M��S�?�z���q3 �k�$�3F�cb�`�RwTRc/����S��3�l-:rx�oԘ��v=Ɓ�/� �����UpZ1�e_��D���>}�f4����V�tD�w"6�a��\�j�{�K4A:�Aba.8�䉼�@�V_���R���i��H�����3�7�H��C��&�����2�y�g�l����X��=�����{��q2MT����;�
�����1�������'�.�EE6j���PBD`�����!�9I�@*)������3ì � Ǐ^�9�$TU#�V���3�%�HY�]]�����)�	B�D��@{L���h�+(��"�����Pj�=&�CO��L�E�,^^��e�j���\d�K����_��ˆԦ/�Շ�vM������d���C_�e���͹1���M���Xu�la��j�C����D��[I��ωo�q�߯b5̋z5=�1k�xu��&Ԋ�/ˎ�stg\�1䙟�ؗ��_렑4C�۔R^���K�VfQtJ���+��;Y�L$�oc��*}�.�O�B�
��GVǏ��ɯo�mG�'���(V�?���r�h�6��:�*�,D������C�6yS���\��DUNe���|��e�/�$N�h��O����d�>^A���v0��ttZ;�%�>n ߪj��т�=� �	{��H70��MY�\A�r��sPϭ�urs��G6� _:x�5��,1	�0
���}J�ga�Bm6tΖ���r`���p�P�n@VŒ���!���R�_,�--:&.�vy&�	�΁
L�Q�����Z�Ȯ!|cM�3�N#�g\ev���Ku�Γ�b{�����nM駿	�)}�Ib+q�)�|e����^�n�o��!�Ƕ�y�4�����SB�괭���z5�S��(S�W.~2.$��36��R*E����M�g;�D|]���<��t:�̐`�=ڋo�l�H���߾�`��|����-k��%��)zU=�xqmǯ;�3��Gző�9X�9n$�#K!��{7kp���}��J���x��DO]p��)C� &F?H�^}��xѠ�ݵ F��S�%����11�mz��n���(���Dd� ��-u��-/��Aq^�~7�s9Ԩ����-z>'��G���!�e�d%�i<f��@�P��>O:l���҃���XNd���6~�����_���Yx]�x����av�����C������\��a�W�υ�rvRs���\<C	�����T��fT�-6X0A�#8�X��Ѯ�iy��	��j�˴�(�\+��v�^�-����p�7��R��� ,�)�}�cGִD�+��!�|�\Mqk�Ŵ x�_�7Y��R߼�`~ڿݍp�C8�鶡_��[�.@.��>��E\���\
ڈY�y�K����E�]��;��6��)�����/�4�\���Q 1���C;8"2�7ؚJ�?�90�� "V��ۢh�
,�� 6��L�*�"׾K��ge!��ûA0����f��|�����،�6��s앒�\g��K��.�*���n���S��RB�*	��f���m"���u�.G�x�NB�M�:�X����,�.�f�/%�c,��ٽ퉁j`����ⱅP��#*�o�o���h�d�9s!���C4� ������6��#D>���I E�04��x؇_̋��v���l�h`������W/��OS@��s�I�-!b�v�S���<Z�������!!#٪��E������/䇛��{���B��]�N�d�5�pMx�gfٲ��4=��h=��fƲ�E�F�vO��p�ng֦D0J�18 a�ۋ�:�?�%k�hX������i3���tu6[�%ѣ�_��h.?���* ���i����ǭ��|�3��Q����\�9������s�L:��E��3(��!wM!$b�#@
�����9d��4���1��[4����%̡ B�Ѓ
�~��.� |�������W��3���*�pv`|���%VWz'���o��|�=���[�