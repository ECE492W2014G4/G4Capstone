��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>>�Htd�����CB��Y�a	��t�g�0e���������u�7���1��7L0}�d��>�n<ǐu�
�sC38#�1jŏ��z�(��sGvL-�~�� l�W��+��8A4�R�['`�p,/��K#8���U��k1|a�w���_KK�O����㋔n�_�v3���d�J������Yd[豛g�U����AV�/F�GG�y*��8�3�u�����q�N�}���m(�t. �\���!�p��T�q�Lf��� �"��GU�W�ܮ?��7�y�0�O�X��}��E�[�f�/D�*N"�Md�ȄM�!�%���7��@�Ыd�X$7r���a���ç�R�2���t�f�?>&[�6C+o��#У'��K"����W0��G�#���pb�!kV�Xr1�~�&E��Y��E�o72��U�HZ�NH�Xc�Ҙ(=�g549/y^��SS�G�c�Ix�Z�@t��?�������	Is/S��ڦ��7�vN�H�GB�	}�2�)�V�筱���7�)�EޝQ�D���Q䴄`w����� +��*�TǺx�c:uK�z6����L5���2) �xd-��wlY=�G�v��d��'�2䠋"�B*-Z��%h-p�f?�����k��ɋ���Ŕ$D����FhF�
�c��~?�%a7A��̫c�Vla�裎��sv��ߦ_�9��y��B;���"P]�Lx�Մg/�Ӌ���xɀ�c�gPDG	�t��o��E'΃w=�׺0�n��j�R`ʾ���.b�ׅ)VK��?�it"�7�P��T@��E����aG����Rx��Ǉ��M�ʭ�rN�wxrf|W��"�e�G�@J�ީ�xﻗ9�d�%��۫(^>`�N.���'�gK��x��%IЖ�?�ZW��|�����[rf�R�����U������I G`Vt�=y�
��-o&
'����$l��|��j�G�0�w�~�
�S8C����1.<��6��|+A�^�d���$Ev�f���׌f��\j� d�j-��8C�sjE�cګ��v���2
�l +@S���ԥ^�� @�ubo*�Gvd��Ǡt��"�����ǫo%+y}Ԥ��7���k�6<����kQB����a�w�c�B��1������ع�AJ	+���$r�����?�⪇uk��>��,˛��dI�&I�� %X��T������݊��M�U~��
�MsNqU���p�+����I=�}{c(D%�>��b�6?E�&>h����D�/@�O�b�@�h�W�w�A�̨$�+/'ϰ(yF�F���@1Gs����=,���A��'�v{Om�ߚ���{d/�8��{YV�#l�����`���"G�6���2R� �%�bR&fW�kQ�p����Pl��Ì/��l@�Ҹ���r�:SR�gE>�֍�Z�(�� ��Q�Kι�#䄱S#/	&�F�%_�0��tBT�^*3���wؒn�� �ֺ�r� 
uc�y���H���aXk[�5�����:�5��L݉ߣ��H�m���e����.h#�'���!�O7f[��KBa{Ե�-ȗ��]�z-Y	���Vq�ɆO% Jz�����6oaGzr�'���5�S����{��(��C�q��E����f��C͂ ��ҔR�xH�J%b���
0�\��nئ�/#	z�Sv���*��[�*�c|ˣ���:����`�<�Ȉ��v�bu���!��"�z�w�ue���5eRA��)�<-�����B�bym@Ϳ�ԅ���UA��k����&�E��]	�TO'F	z���5uHdv��"�H[����b��|I��A(�#|{�m���~�u�N,R��iEYe���cy�)�_�(�`l�����o*ަ�<3�D��"b�yg�Ax�E*��%���r�F�����<���;f+O)�Zh��ŏ�,��8�����7�:�
iW8uz��t� ԁ�?Ws���6S)��z��U�� ��x�)zA���Eֲ�/�惒1>n��&��|�q�@��yI .`�UM.�ψN�*����1ӷs�F|2C�uY/ַ����4�&g�T���Q����(%Or6�,c���^���qǅ���{}g3P{�[����h~��$�6�vM�6/N��e���cC;'|X�a�M�L�H���VϬ���K�۲����՞yc�FQ��#d��A�0��Y�[��gϔ� �:&��*cܠl�Q��^j��*����K��F�3;g�f}���i:�E7ׇZq���kM���!FZf�~x_�L��_�A�}L��^e���p����'0�=�5]��'�?i�x������L�Mü���PnzJOe�Q8�e(0ӲJ����×����w��Z�.r����]5�������'.@���*r��7�l-m��3u� @��	���MR��j����{�}TTt�U�J�ݔ(������p�b[��
`�w��}���n�m�%�w��B�@N���u� ��[v\�nP��ڵO��PK�$-���Jg����4�\�V�*�_@��$�Ur���4�F��h@{�o)�
�q`u��G�Ӧ�i��7�'�xu�7$�۩�-~3\uc����-���E,d��ߍ�'�=��Bl�2�Ó�ː���ϵ��|���o������
n%4#�ۻ�z�8��i#�kaeS���"��m�*��L���Y+J�+����b����?֚?|�	����X@��ǺSw�-���� �V���1��s\[�\NH� �2Ç��f�9���e�Zѣ�ll�.{�R���3Ã�mX]�\����qB��ydU���UkΩ	��tM]�^������8����e�j	$W����;?�y��#��n��$f���zS��य़2���A9�r1T��؟F3�����V����В�[�@M	����P�*���F��v/r���w�y��	ʑ�<�#õzE�}`�_^�Ƀ��VH)�y��\��Sy��� n�O��B��ɻ���'���ˎȉFڗ�z����zO.WlN��.�a|��H"�����9��V���� �^I��*8�V'}�<�!�<e��i�L�Hf���?��!Q(6Δ��)@+O{���i>�P��R�]C�����Q�	/��nn�4�z�}����
�� ��2�ۇ˴j��kq��;�%�5�V���3S>s����6®L����:�]�q�� G~(ovy��� s�p����5B�O�Q.��ll�QB�eёS$���w���\��zF��e4=��xH�ay|��4h�(��,�����4����ЁXŤ������	h� ��Kϝ