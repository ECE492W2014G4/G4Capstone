��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�"��F9s�`&���a�oq���F�g�O�]�<ݲ����eCL��D���{�5��8̝DFI��Zp\m|Q��
�}�6C���UnF:<�jΈ�2�����<����sf�k��,jڙ�����2��X��Ss�HL��	�������+g?���N�Ż�����|�v7�{M��VNB
��Rs�゙�Ld\��X�'��R :�J���^�����kMkx�Q���3!P}�e���Z�Y?.�U{�RP	�)��lI{tI(S
7ZF��:ȵʁ�wಿ)��ךb��(���R��,��P��Ŧ��t�f=��ς?�#X���5kv*M3H��u��M���Kͫ�%e��Q~L!�t�M��,�����؄��
uz0�� �9\J�m��n�'���Jc�Ƨ�Z�=S��:��H{O�s�H>An�Neo8����Wmt�?u-<�c�.�%ڛ\�
97$�hr����E.�Y�b�T�rW���ߡ��޻��V*��1��"�}�L*�M��NŁt3|���=މ �����{�=�4nœ���NWN�!7�������`Tv*s�M�J9v6&�iC0n�/�z�~j��.�7���[[��B΢�2�Y�l��.!S�8�
�L�l���(��;���X��2JrCf�,�8��^ӿ��С��|#�a)(h빾�w���T�D�*[n7�_����FE���C�
�ViT�XC�I��m	�D����YBKE��FC�ö\x�(J
[~�/n�N�.���-B���UV��.����+L*�s3�뀎��N�xQEH S&����������R�o/|�z4Ow�l������2Y*1=ͮ�����X��N��i��z�����$��%gu�w/9�uH�@N��*�{C�~%�����]��8�,=��[�\�>Lj���<����n#IĄ{�c�3�L��x&���S+'�L�W���o������2S�+�Obb�(��<]o����QA�Y�V*��n�, UL�`Ƃ��k�!0�����#�LC�'s���!�1�})p�����w����7�#�]���NB�]Q��m=a62��ҡZ#�º��l9e�.��P���0lj�Cڞ�T>p�Ypo��0�ZVȐ݀��4���bMk��v(�:��7���@�%���A�oB�Z4T~���	Q�Cx] �x�=?@n��17�3������aI�>DJ,xu�����8J�}� (��A�2�g�Ä�,_�$�h�rI~>�a�m����i�s<�K��A?��o��ó(��NTA�&Ɉ�w �V���si>�,���_�� I��Mr:D-2�0�~�T�r�'�E�O9A ����!�oj�<r��C�<�uZ���o#?�eCfp ��6�V�[v���z��Qk��Cg+���ӇJ'�ꂹo@\���\��ּ��@P��߼*2���n	a�8�ࢺr:��S��p٩��B�ZdrĦ#�3B�\2^Wpa�.~�Jv�Y�w���P~��;���%��v��d2�����s:[.ѓ|S}7T����ʟ���ÎZ��Gؓ�ņ�ly �����3gˋ�������I������"����9�0m��:%H?�D����ڧ}�K�+��ݚ�?��M�ub�R3�G,�hB@m>>+3��u,�{��9R���mQ��{@2�k[���Ifl
�}�3-�
��L��y=��Q6��	��OG!���C��6�C�j�!�q�a"zHΪ�q�U#Dx\b��:)wR]�&�Ҹ&3o��S��$H��P��zE
�ɵ�����Z�2)W�ɪ���f�\�{�]Q�ڻ�gԟ4�=�$��D,��M���|�(�K��+�������+�I |E��o��nr�-Z�OQ��t���o�!I:�J8�OL��Q���� �@�-����`*Q���E6��L�-y����ͥ�fN�s�����%��Y������j�]�{���/�5�;��;f1~F�*����\�S+��d��������0�q�x*Zl�#���H|U�U��	�
'��椤 �j�A:���Ο��P�	g*\���K�r�݌�H�Җk�M��tT���]�׾�[�� �����۶%�r~a�Lr�\K%�
D*�V56����t�{��.�]8I�}YQ&�j.�!������3�&}��`�i��w�g��(��e���h��40�K��&�*�wqv|^�Ҏk��#
T������/�,��Ƕ��?�-6Yp�w�!�x0Q��O��ˮ��O>��~h�ށ����p�^�u�N�K~m�x�i���#qfݺ0��B���H���n�t#OTi�D.���8���.���\�7���������Vc�,��Xb纟�>�� �*���k�]*@��G����m�9E�m��áh����Wh��N��yC��z,�'������N�h
�.t�p'��j���H��m��(����v�#��t���'vq���y(��SAb��^�󿽭*Ak[��q�/��	°�p��b�lY��A������1�����`I8-G�b����%�wz��Z�l�D�J�����rv�T�j'?�L+��g�>w�����&~"�t��8�k��+;S<�;����%����+0!���z�&J��o���O-�&�O��'>6b��سF��e��^�	,����M%�N�^�(�]q)z�D�rrR5`��b8������7����dm�m=ؔ��a��#Ӛ��^����;�7�5�`�Dٹ|��)��l�
J!0ǎ��Ω%/ܤL�Q&�}���%M�r��G0�*i8�-[[�/�%+�Y��O|�e�A_DEΣ�~mhW�膭ݶɰ7	ڑ`g�w�B�>kLL{�?�M[�qr�;��� ,����V�"t��b~�N�&	��1;����2v�C^W��m7���݋{U����_.�Q�r��VQ�2Ps��x�.�D/E���5oՓ�a=���~��bĿ��%�A:�����=�Ѯ#�<Zl�`���:�A9b-��(��l��{�`^;�'.�cԐ��s��������m��``i�Ac~~�e�~^n�K�e=���ݰ�-��},�l����q�jT}�R�/�P�Sx
�?:��E�8|K�F`��(Q��xt�������rMLe��I\��2���[\��)�7��̪�į���}�	v�i@K�-�� Jп��"������SrqTK>���Q��3��ح�ڎ���\8
�He�;C���;�f���mCB���x�