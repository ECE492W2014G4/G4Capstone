��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P��v�"<ߞ��&'��k%P碶�R�ӣ�sĞ������FY&(d���3�&�I,o���%�Rݵ7�7즉�2�Yij�'�ԑ)��ۀ���m����Y������}���%���1^�y���qߒ��?Ū�F�Om�m=HJԐ��	���~�f41�>�+��u�0�2�`��ަ�rr�H����:i]�2z�;��8	2��yq5�?�:�Lg�A��Lz�����Z=�=0@kD�Y�%�m�*k;�{�H?hVj�֛�7����\u��ڻ�#��+�dS���M�;i��E�r�L&K�\����L_��0�AA�׮���i���1�9�׃]�"�ܨ�٨��ˍT��]iMe	
���9�n~I��*փ��6KoLD�9����I�	-dL�6�1@�(?���*����|@t5��7^�&�[GՂ�J}�(�� WH����1�_��'��Er�J*���E�b)�XT�f�#�S�����1��]���a�v2^Q�sY��`9W��;� ���*����*��fnO�~�x��	�o<�G��+��8?��U��暜��D�;�>��'�3��m��>��5�!@��JL�E�Rê�'#�!�"����(ZӫЅ�q����C�\���@��Dw�����;��$��2�6I�e�r��9���CamfP<`y��+f�B&����J�A����5��6Hob���.GZZ7�zә�(^�֕Cu���0 [$�7{�5T$���+p"w����2���er�b��^�NW��E�@��&���*�Ö��y�W
��iG1ƃ=���3�t)g�&F��D%�i!��%ꅅa�S8�[͟"������krLH��z���N���m�w��� k�]}��39��J���@���[�U�R$g�t�Ol��(&E�9��Ae����B���@�����;��K(������1A��3`*� T�?]w�$Od4UH�z磣1tv/A�X��' r������/X4�2��~��`5����5g+B-U��5��<}J�b���������r�������-�#�#6��Ɍ�]3\��'��6��|P���������|o�GY̅�Qö�ETD�CaC�g�f��¾���?���[]"�y�U��(񁻍*�/h��̽��i�d���m�OkNO%Ͱ��>S-�A��o(f�>3|�6�ް�{�{��dg��R{70/�*{L���2�{s���ۀOK��6�Fn�a�	>a�V}ާ�JBh�z�AN���̭�
���#ge6�细��ɶ?YH5�,x8,tC�8���j�g	��"͹0@b_��k��.�	�nј��d��BA�����zo5�$��9{y�ؖ��tŵʖ2{r�w^.��vҬ�7�� Ǿ]7����~[�5$i�[�x@L�X���� >����,!�@p��c��{ʂ�o��ρ`�5�����"���^6ZK9�U���sH����Mm>%��By�}�Sv��a��>��;���5���6�Z����5\]D��g�1ֵ��[4�^&:V�-��_w�j��D`����:��۫O�
�H\(%6u��x����&h��(�(��(w_�V�k��4;�|��@�\�k���*h��Q����0��P�r�}
�dq����o���^:#7:1��1���PrR1��J!�e"B���}iv+��N#�ر_��#o�:?���%R_ku"j���H�l�_'Π���,��1��\ĦC�MĘ�b�m^���m5l�����˶l�3�C,/���V�#��xA6�j���g��+:`7�/��-PEe�����]��<d+ӫ�V�B���������l�Zm�ƴ���@u�y[IeVbl���K��������S�5"ͮ���Z�]�|5%+PSpͺ��/C��E6�<qj�A��v1Ryy��@Mp���r�X՞���U�#D��jc�V����<�`�U�$���a�sك����ݾ�E����D0ھE��Q����������<&]MOBq(�Ky��n'�KO���y�pw��x ©������摆����n�rIn0�Hbr�|.k����:	 {�W52��F��D5�D8�O��Hp�_�M���e��6_4�Vow�sW�Q �-��ȫ2��3m< � ,��+�o���HϘi���M�yq�xqd�r�k3p+���`���B�أ���&���_��x��(�;/Z0p�R�A��1�/�(g��l��㮼m ���04Y�W3��طhP��������g(OE����0<��&�I��3�z�mbZ�,�g���_VА��>�7�����\0 }�U6��W��a�-�+�W�Y��q���~g����.$��y��s��-��?r���O��[)���x�v���[����m�s�[�>���U�%�8a'�}�J�=�e�{+h.t�}�����ȋ���A���a� 7�o��N���޹���DE�"��ϙ/�.GTGfv�|��d�](8U�'�t�����
�h���M�M�ISȿ�Bp���v�����c�����'�G�
v�l�|���g��I.��gē��a m�R?#W���O ,�d-r���c����)W 7&G�Jo�
����L�kg��ǽ ��k���V���iZ$z��X|u������X�-$�@���q4|�ԮT����c�<n`��G;��1�ް���W��c�hs�k6A��i��^�H�Y��H8�W�k@ZJf���K)Ri���G_5^�x���Y��>![�v�zz�)��A�;����@B�Kf��^"�µ�lKDq����[7�Pv;��>&h�^yX@�T�o��6o������ѡݏ1�.0�t7�����mFC�VQ��eb���┉��n�#�"���j+�^t��h���-f0�Fk�p�Y}�|�C��3D:�@���
�Y�p&�9G(>��w���)k)�+]���pb��Ӵ����z]M�"%�TY���jU�#y.�FF:�4��Hg�A��-T������c�g����ZM��o4)�+��/7�z�/�і�ޤ��ꞔ�s�Е#��hWȆ�R�0B���j�
�U��
nE��E�W+2̳���o���w�ŀ�����T�f��Ff���mΜ�(kXHfZЩg�eg�zq�U�b�U�wq���9���dZ���VYJ�Aj࡚6g���h�a�D ;��&�Q�#Ǵ��v���h�r1�n�$�B�hd�6$�!��Ԧ����8 ���9`��O���CO��ڲ&�!L�t������B�䘿��&#s*���}eU��k�E4q���U��P��1c��2�����A�~�	nP?��麃-6�*��Dg��K�帆���`ȸ*H41q�+K��$V6N+��Z_��S��"�v�nH9Q�.�ʙ�� ژ�2���%A�Y>�<z���E��p�xlpcm��G�8lڳ���E�DAŜٴ�0č�4&|	[��+��C�? Ϥמ��b��d�c���y�V�:(�F�RB	y%}��\W$��U�KΚ��׉��}`K�J���>g2t����ֹ5%fY��ⰆN2���U0�Z��2_I[1)�2�.���e��q��d>9�̸�YJc>u��c�Ѻ� P�d�i��{Hy�z���Q��ͽ��C��D�9	��4/k�՞'���}W��rp\�<��B�����jMh�'f-�!�(K�����w7�����n�hJՆ�Ӧ+�∔l({�M���x
��m��`$���9=�5���N
����#��+ʥ^o7��"(~����R����j~��(�V+'����)"n�k�#֭5Ԇ��s�-w��Oڗ�[���/����tj�I�tg��8�lY���B�)���,i��c	P�j���" �#�:�i��
R�����	�@��zk��/�&������U����z<S�B�n
)�<a�`Dӎ��lw s�|�\®�z��^���{��HFń@Ǻ4�ɿ8�i��`WUk!(��'���J�P�vY� %QB<�#�$% F�������u��� 9D�����a!�y>�u��ހ���6���2%��2W����^`����>��YeD�/�<P̻�-,猂-;M���s>��@i������?�����77'ZTs�7e��~�Q��P�zs��D˧�^K���U�֐d�E�_�1d���hl��=���t#��g��OzoAI���A���aX)Be�h�>UF�B|����
b��-(׍���#R����qQ�Kzt~�M�Ґ;��\�S�I8=�\	LQ jMT���\Y�e�G �����;�/!jZ�د�=��<;�z$f���Z �vm��s({��[p�K�rS��9(����(	��8��1��=��� ��7~r���5X_�܋.|�{ϕk���=�o�ti��ƽ�ߑ�(�i$��
�c�
��*�")6�}�T�=�����r�EG\&W!+���|z���/J��б(��!O�m>�.��wE������{��e��,��(�>˖'X�D���$��SQ��_I6h�T�L�y���Ot�cRp��@J&n��W��&���C��L��S�9���d���Z2[�ʞ��mj��1G(���'^�����֌��}��Ǿ�u%��H�{�l��#`�ϜߨWD.�=���ID�p܅'�BHJ~D�O�{���4hm�o����Q%�	Ta�nZ�5�%!-�v���_�ܓ������i� �o���s�
*	M�&Ghj�T�=K̅��zY7�x�I�������L��쇧�����Iΐ[ �L1�ZP,����ƕ;��,�i�60E	�
�gDnޅ�'5�5r�}RY�=��զ���	X�Zb�bW�U+�V���T'��\��_�T:X�{dqX��`���`vR�v�����X1
?������k~L$�j�y��90�<v��&w����4��@��>�0r��������T�a����t���x��xd�e8~�2�O�Tn�<��!|P2�>���}�E��\z���K���9g���H��w��q������ZBP܀
���ѕ�n��1�9d�vV�[c�����:)� |8$(ڊ��r�LQ�l`]�bs;��/
{ۆ�'���f�g=�J��D!�N��q3V+ԋ�L�^9��,jJb6Mթ�*k4����م�0 /~(ﺮ0���}��@�+%{K�|�e}�X�?��*
�^
�Oׇ�ٽ�FVc�Pp���J)�z.���m}�<�AS�(�٘�����
���t�-����M�&���w0�7�T����9��6}bD���-�_�o/���+�A���^�yX��h��ħ�p���:�3b=E}5���}�	��2TU�!l�Q�3�~���`�B���YJ��\��3�B�5� ��GᓦE���	���ނ���~��d̒�dW͹�O!_�S\����h+����Dޞ���b㍫E�� ��oK=�c�ee�W��Y�>p���'���Q��}��CZ�m�~�~_�S���a��6�t��� rV��o�@ H����Cw�2���8~T���bb#N��T6р�ums�F'���P�}�����exM� �* �`k�i$�ͱ�zZ����]�����=�{L�a9Փ��A�6/Z��C���;Gc�^E���(S�g�٤�������i��!T��`]i|��rn2up4����Q���V_�đ4�������]���Ģ���hd|"G��EKA����(hA���5D��*�����5k��į�ï���:+x"g�d��*�_���CA�Qg��B�1D�J`�^5 �l��,T`���=	��ja��*��^�"�T6����NU�<��t� ��F}�L{9�
Gf!�*j�p�=Hj���-&@\���!���Z3��1.�����Fn�7�+) la�xV#��U�D�����^��4�].[FG��Q� &$ۣ)���a��Z�(�������H�����Co����Pob�&AU&��6I��E_I!}�w��F���B��.���Yc�����ʹ�ȦX��-ET)�����Q6��<��ĺ�
��v;TH{W����>�r�g6r�-��wT�x��l\h����Eu~��)�%�8�lG-�]!�����4���זu���>ɡ|�/�o_b�0ҍ20��m�Pku�@�O�M���Ȁ{��M�^H�����ݗ�a�X��ܻ���;M�A�X'����17	A��o(����ظ^�KQ)�q���bR��hiw�r���
���xS���Ulq�,��EQ�� ۈ�)��9 ��=��\���j�95������糂p��p1�W������f�,$	�����b�i�"z}�)��1�ɐs^�ت_.�)e�Zz��{+�L�_,?��$���]�z�&`�S�eE�1�!@�?"�>�q��qiVh�Q��]���VÈ�ϒ��Ш�Aق3��a39�H��Cj�?~���1�����@�~t� Z,o��4W	�M�����o��@��%��/�kC#D(~����w}���%�@GD�[Q�H?蚰~4��	����o�X:$��t�$;�&޶Zݚ7�����%��#�80c��;J>����63�G���V�#x`���<ҿ����V
������dBl���(Te�=�׎�E���F���?y0Xl	2:��MjMr)�������y������9Xv�\�˃���\^���SO�±�� ï7�6�]fd��1\g���ɕ��-�����T ��aA):S2�	�i>.�Ei��lF�������T`���J�4d�]��39U��`w0^��gǻ�\_���{��,MYD���,���d����I���d��s�1pu��3Q4�;#5�����g��bG�>��	0oe/M��H���/,/��4�����`�H�@mv�|+�P��ejF��t��x�ހ,�k=��y�	�N)����g�7ف�s�¥�O�����g���qOk�l�?)	�g����/p��^�+��ݩ:h�z@ ��Bӵ\=�{x�݃Fp�����L��'����t��=?������j�xJ�� ���=b��&�ˬ���ecnzke��A��2Cf3 B��6�6��h��{D�g�%�X�����7������|C��"3�����i�6���A�7�&�|�\�1��\�V���OۃZS���(�,��:��*	��bs�M1W�c�+w�n�Z�� ��M/ܩ�k�%n#�S]j��4��&��ɜc#��� _C�X�C��_�J�]�𠛔��2�PJ�V�v
ك�2�3����tn����[�%=�(�ZkdH���7}���Դ`c��C����,�	�WvV�ِǄ�=m6�ֺ-@�����������c�}ÀDܳ��>V.y�YW@KBDt�"ǘ]�J����~�$n�Q����:6�l�ʫ>CV�O�����Dmz�bk^��G�u&
��0�1<~��>������H���G�'��*���`�#d`����7�Hr�.7�1��2a�3y*L\4��6{�s�p�|�����c�k#���2͎�����,�71R��6;P�D�Np�,�E$!���TZ (��m�k������n���
��g��m�PRSފ�^�zy)�vQ
mfq��\>vh��H�&h��D��`q.�/�۞�b�~{�+U��ҭP�95p_'8@	�4�2@���o=�jP{��@�&�K~��u���]l�4[�2��	��~�G�d��q\��l�����R<�āy����я�(S�Y��ݚ��a�ZǥFv.����_w�:0�#ْu���T]��{�T��~��%^�~�Z.���I��mG�|����?˹��@�/���8q����%ǜ��':+�����mBq�f|���ȇu%���Ƒ�mzY�	t�$Eb�=����Ww�5>3G,��f�t�����l?�Vbb��7�&�NCR{��WQ��Hq¸J�!�(	�%Zc�[�, ]�u����[]f��6�e�)�ѝ0=R���d�&�� ��ػ�?;����K� gT_�~��hz��G�S���)�����☳F���:g�I2�g0����7�@�橖����bz|�c=�pֿɔ��v)I�UZ4rc�|{�Wި���z݆.K�'��H��U5Kv>��~΂s�m�������_��K���
=9��O���W���.��I����{�}{]��R!ѭ�r+B�	�2L>�F�Jӎ�V<���lK����[5Ű���j�KWqD���@׀/�Ds�c���$�7B �W{y��.KG�����_�-6Ǆ�������j�,��>��H�no&����g�g9�!ff�x�7縈1�* �?��L\�`�>;�(�Y���L�2�A�����X9y�ި�`:�+������N�eS�m�8�D�u�b���/$�,$-����*��^��cG�ޫ�m�r���
��&�冠�z�9-��f����vѼH���&�E�T'��P*g?�@Z��dŰYgq3]����=��L���*��4_���7��mDr��"O.�j��\${s�<4"�����N���}'1����d�V���s$A6Q��Я�S��L�`9������������������F���d-E.�Z��q���l���^y�ؑ�?���__V-�P��^R�M�����Q�7��-({0�O�<��}��[!�
۟�`"��w�<��F��?nO�B'N���]���0
/����M_n�%8���l���ޘ�6�4
vơ` oC��՟81�_�m���h�!���v��X|:��Yg�bd�F���4�� ��p��$�9'/�輅,;���{$�E��&�[�;�D-3s�a���@��ۨ-�:��.� M!��$(�j�a@�K������aЧNi�W�~`Mp�qÛ/h�´������>�+��z��S ���B���b���`7Ϛ1Am/�����D����1cfƣŭHc"�Q�y�.�)�C �GY�K��lo�;���"S�p,�eS�
B	�.������O��,���hx)QV͡׺�����j��2�y�Q+Y�K��g�L��Gqڭ�Z-��5]\��
?�6��|��W����֘6�f��pO
��AdOX�k���������i���g(��r�C7�qa��c���p�!k��m?��ӷ�~��vͧ���L���wdt3��<Y��q�j�,��$�Ws�E�3�j4+���ԋ���;��E��YB���{r�/�1H���FٳTO���>�%���9B�*-K�[H�\
k[w5����R�]���da��h�7�U=�H$:܆�UhT�{�<�K�t9މ��P�>�7O3����"YQ�V\���6����l��񄉠`澒���cÛ��S�Zg�@b����-�$t��~Q�!i��l,��?2�ɧ�0W�W��U�q8�J�_X��NY�W�e��R
p��+-�1�a���n�E����>$VYأn��/9Kb�"�X�K��my�dLi�c�~������\=C���l��v����/:��
pA��8
��Qe�� w�7�P�t��i��r��N�RGw���W�G�p��HIitT ��\��	�k��YCBObp/��r��S��N�[���qQ0����h+)�k1+��
Hͳ�EE�P���Ī]k�}�r.��%6�؞��m�I�/@��wYN�ؔ�t%��V~'����Ma9l�f~��G��`&�틻��W�'Η��;r�n� gs�c"|v>�I�d�}U�UÏ��.k�!U��c�?~�an��ِn������y��A��BVg��t_n�O#ui��s���v���U�V&���	��>����[X�7����V�����هĳUe�Q���P�$��Im�[���z5�p/�s�D����!U��d�{Jǽ�����ѿOYg^�����̝P	�,nsN�1�-��(�NW�r�A�M@�M��hNre��9�6��&���IGv�x$����׍���k�T���V_~Y8n�ϸ	Zxg��F�_��$�B���b��g||]�2 �;�dH�U�V�� ��j�5[EW��6Na٥t�Aw�WRw�Г6��z�����Aeiu���߀��A'�֚���soRIjx���ɖy����i��r����23*�f�,J�Y2<��5k<]�Z��]�z�H��ź>�mtB1G���C����j%n㔦����԰,�O�A(��)X�%���Aл&j=�s�;����'����U '%�k~	��L�SV���c��`��ǌ�{�/�!(&I�
z���>m}dI!K�`��{�*����n���L�>�I{ɾ�g��
ߌ-zk��g�g0�\1��%�[i54�Lo��{FU�Q�+�y ��){ �5��
�L�V��"-l��u~�b�X�د����i0�ƏF�S�4�p��8*ҭ���K��� r*q%#���&:���W$bU��Y1�w<���X���^���즏~j�t�G�s�)�il��H�0����k�gD�Q�/���M��?*�נl�OiU��U���t?��B�x�υA:o,�Q�ߍ�YP1$�{�Fm�-O�vN����Le�O0���l֏c3������`�<��v..�����26�i����,�Yv�ݚɩ�̼����	;wE�������
�{�5?��ɚ�ߞ�� ����E�`��������EV�~H;5��ȸQ.���Ӏ��&����T2pQ$"���F��l�Wc3��Q��Z5���&,�q�?;��E4���eն�U�fެܲ�;)X��X�(̅?�����K��O/�2P��G�YU�ĸ�x7~
�{K�@!љ�^{��.y����YX* �)�B[���x+�_-Ng��@�gSŇ4X�,�A���}��sC��	��4��V	�Ъ(nS`<���Z������ҫa�N֐��N��{��ݛ`�u�.�M\�d���SG��iK�d�h�.l�,�=+e�HGn�j��:ݓ	�������5�c���蓨�,Ae&�)<��T����ݮ�Q�7�좹�v�N��)HpdSQ�.�ώ�$��1n��oˀ������������)t:-Q�v��I4�>�\Fol���>YS���Dm����j���}��`tG☻m�_��e��u`(a�mCg�#�u2	�.���q����DAU�n��?� ����̇�g�	��x1u"L���hf蔁����z�����MT�i!�����iK����=S��;��&,<����K�fY���+0,N�t��S@FE#2ޔ9�1qxO,�/�m��0�H��>;g�ߞĒ�NK����F��7��w��I��,��!�r����%u��G`��/�J��$�a��K��Z�%1���(����諲M���@�9���p��4k��4r�BQA�t�CA,�Cpx�#�#��K�}*C��R��5}:����j?���x����� �"�ɛ��:��D5p|��xg����>^�|���R̽�u�첇��,��2�-t���Y$Jĳ�؞=2Mݕb)_�X���)��k�>�Ne�w�u�$����Ż��րQ�+Gk_w�m��>�aZ�;�|�O!��0A�����U�%se�7�,��ý�86%�J�3�`[fO84!*r�_�o��P˒&����U�k�ˎ;3c�+S:X	X������w1C%o�f���mP�_2s'3~4"J΀�#��ОQ;�N��DpdGp�� �@�DH�Ct
b�� �G�7zڋ�	�ݚ�C�ܦ.(`:F)u�_I��^K������NLM��%\�ØM�4AL]%�g�[�3�!,Y�6������Yr@�����5ܹ#�K�+v@]���>��
���h꭛��w����g�)�M2���X�����h����JT8����������C�v�NY�B{����5�(z�3d��(l��ѭL��(�YL�i7?�3��i5g>�2:��o�[p<�����w`t-4oňnhF�r��>���7ZJ&;N4B(k�����<~���T%漆�G� v F�Zx
�y �꬏Y��%�oU��E������D($w	G������`n�Ϗ���'4TJ��TP���,�r ®IU�Ѐ��=eOf7����vE�"����4}���A�ƛ��?�|�E8?�أM��Gou>r��()�R�?�!�D�Q�r�nz1�ny}��A�~��s��i�i9���N�S����i���� )5��~2����hy	:�1�|_*����.�UQ�b%��y�f�?���ީ/n��8`r�O�F�%��'1&�T���ӊ����F=ˌ	�,

��M܂�"�to�ٯaQ�B�HI"sBb7���
�ʧ��>�=~	e$������.�ZJ� �,�a�$`:6v����ؾ�t�
�9;��I��H��DC���gj�F&rMAtew.{���o��@����^M�^{�\E�\o�D�_Lzh^�Q�j�"a�2�UƼ��a�3�E�����e�p�o4�u�Y
�Qf��zy��#��:�b���!�!.��0(�]$�u}�����<Z��m6_��]�&�62��n�D��d��?�'"�����Q�2IB3")U64�$�W���|�k���"�:������Hʡ����JS>|�V��r�tkY^"s�����vʦ07�a�%������j��>�֕x��/j�����"M��ӈk.��;�-"4&5�[v>�.(��\q�6��?Ha��QYL��#��ӵ����	��XM0 ~��~`�쬶�Kƺ7�E�N��+ (R�����:�-\��;�����c��>t���y�2�֮h�}V�L�i�_�%g%�����V�;Ә�e2H�.�ޣ�w�ײ�'S�C��\T��>����GQ�����X��rs�N�E|�7�_͠IO�c*s��1����;�^�å;���Z�ݟ�s��:�o�x���Qao5`����}��F�P���O�`�L+��tq��	��<&�?��	j۫���p�E�ޠ`x��㨇Jݡꝗ��[������Jm����钦�(p��~���&u��|�*���TY!�y�!��2�l��m��M�Rצ� (��:u�ʎ�\� 4����܀u�aV�}�a̶_��jw�2	�z�@x�>a�}�ڙX������g(���v����Q���a���L���iZ�I�e��� �����e�
�d�3��X�e���O2S5ٜ�@��@3�U�D�E$@��� K�Ƒ֏��Ȯ[nӖ� �瘋�$j�}��4�K-b���T��ͿP,�'=y(����sl�@9�����8��Ӄ}�A��A���'�/2�%�(��/=/���J���v��� �h�}��"�c����(+��O����1y�D�����&	��*p$��Q�d�q.^~�nI��۸n�d�M�	4f�ݰ�8)�ت_t8.��2�N��QA�3 U� ���w5:�Qd�EE�����kiV/Z�q��4���;��p�S���D�-{�hnS􀸯���4�-N4b�������9$�����"2&[�2Yw��]�"��Y�=�yy얤�r����x�lg���r��Y�N�|�&�,�Z=S':��¼��Tݪ�^�ٓz6�F�M�p�@ߥMap�en���qn���k�`#7���!�����"X$�6����R��=ħq@�� `���%�B�3?��*���(��v�R�Љ���MY���&Z$��0�y��Ȱ2�%�H�����Wr�-&�$ ��-�Q�
����VS�h�������-cRKI��B��W�
�Þ�+�(X�(,��ޙ=˫؋D���UȪ��P2��W��'��d������FW��j��tF=�"�H�mn�C��g"6wsq��w��oO<;���T�U$���m4F8Fѕa�d\%�6��������44>V�%w[F<��B�erg�q�[��T���F�=aJH�oĚ&8ub���7ti��ME�I��I2�0�y�!�,7�و�y�UR��N�lѝ��F]+�TC��j��V��5�T.g���*2���v*�cU����)8�ڧ�x[���Э��qXx���|���3J*��S�R�a�����P}r!�8���l:���+'�Z�膃vb�K���X��+�V�>�9�ԑ��BaJ	�3�noB��3�����U�>�rFdsg�âjU�dwW�X!6ːe�� �����e��4-��i��"=�;yNH�A^d�5͈�.�E =�8�z&�U�I#}�!����g�9�Tb��f��N�\Jn�싻O�ͫ�sD2�p������%�06���=�ڒ3��F��KD�,�M����da�Nfj&y�JcG��BE�O�O�3����)~$ ����v坊��'�I�O�����4+p�/��%�o���4���?xԈ��z���ac�g1����{�A��������;~f}��4��<(9�|S3O�^IH9�D�V���X:A_tF;���|�n����%�!�)�����<��%S���U >�M����*��g/�?���u(Oh���;�%�}���3� �:�i{g�{�m�
��Q�h|Aqr��x;�#ff�{�W��m;�R����.�G����mr_���I7��;��,(��x!����y�H��LM���	^Xz�(޷۰�V�fӨP���xѧ�T�W�O;bg�<˱���f[�?���bܿ.i�i��(Gӫ}>�o�{lE�"�Zl�����Yo��5����������L"�`�$��9����V\~q$۶��Kt���L�Ҁv��j�  $$��}�+�4���&�`��YLdD����#����CB���&)�3��;۞�p���G�蜽�a�Ʊ*>R-��٫U��X4[�"��������Gt�	�`�\���1ڎ�@�]�����A�8�h0�æ^L̛@��I"a1�iaxd��筝�8���9*�����W�wE��V�)4e�#+#Es�(�k� ��A+�P���	f9��;$�}��	m��[ƻ����^c����pC�9��ţ�x��nhB\�w|=\#�~����?r����R���F9/�84�$^�����
��6�}���^��HӀ�H�/B���ða��,�N�>���%)G��ak������V!����b�?�a��U�d'� �r7W��j�S����q��_��W�m��o��ǧ��i�&M�S�{vX�.n|)�Z�M�R��)�����zh�xk~�ݜ��h�0�O����7�^b�nr��(�)O�#ť�ɧ��#"z�F���?�@\�!���^�������`w����́�޵�B`�3��J��������B-9N�5CQ�Se����8���A�,W�R�6���\�¯'�y�>Q��S���)��q��!\�'Y�zH�vd��/R�T9�#��;�\��P!���JW��>X��P��W	"�vb���㵓/k}ҫ���E��:w��~�x3Zi�^�.��iA�ɲ,!�rQ##>(޾R�[���:�̴)��o�����o	k^AX�6��D����l#�@�$�a�8�Ƣ=&2�kd������`m���'�~�q��Qzѿ���B�yTtڠg����b�{-�?qzi�f�{�7�{%��2�JB�r� �NX�!����,�1�9��\�D`
z��I밬����Ü��DYXt��#ed1=0���1��m#��%:{���!,1r\�a�H_���h_0�������gl�Y�_-��H����ն�y�l:'���%�V��Hr�Q�x�ZA�:J9�� y��������9��[� ���6���'�Y��o%���>[��@}����8J-��k(��h֑�@g�����q<{��J��"���!�<<��
�xְ�6�	70�_�{��J��.u���2w�F㵼Ѩ:pfAj�G?��q�2����2~nW��Yȉ���jM6�aO�H'?)����8��I�e���G�*}�g6i�[��!�+�)C�.sfi��kCb��
�i���`	Wcޔ�Dks�}ւ�o���'h;^�p0���,��� FTZ��hn�%c��)_<@�%�lG<�K6�S��Ǔmwֽ���e(��|����9�i��@��>���_����G$;�t�M� ��9^�;�-��s���3�s9���`b�y��ԗ_b�m�����*iy�$EdG�m�]�S=��_~6���T�)�T��l����F{}+��<��8xNx��[�k��3��4�!)��yn�iT�4Mچ{	��AU�|��)�R*�v��M �ԙ"��u?c����}�5*K��o����Aύ���?�_��~���zB��Χ�ZR 	t���U�)�=�+��=����.����]��K�g��N���I �e@�t� �73V�tw��:lR��#�Ǭ�sC0�����.9k�y4K�ˈ_Eϐ`�Q�u�ӆ�Ku�I�;��]����Zk��4�2��L���ޚ�"��Z�|��~u�f�S�j�Y��ؤ�-�#mQ��Z��*|6-���8?��"+<'	~�σ�1��:ԥx��l(w�
G����)w��Z���$G��=��s�L�����_���/�r�F��b�Ɣ_x+�T#(�Ǡ]��b�E����Վ����bn���u��*��5� �g!���x�M�E6LU��'�=~�����r�S��i�

Mgʍv�Fk��t�^�R�m�=af��@n���?�G r�I���DUʞfv\��"tǩ ����a�r�=����:n�#�Ls��o�����Mo�`
���YO��F`ΰ,\���/z��K j�Ta�an:�: b���!w �O��(ɾ 0�[,��`�1c�1V�_?�m*3a/1p��͛���u�����FZMC��:�]E=�0��]��xSbt���η����|�C8+������b����R ��Y�!@�W6W�繞�oB��9�����B�⦅v�R@IL'��G\D������5vl�l6����_e�7q%����F���Z����A�8��K\;��>��;��)�rQ3Ӡ�Q�<F���5a�.h��(�}�[x���}'�я��=�>;�Y��K͞X�ڃ<~�6t8B��q?��խB��U<�9y[<A�����+l��Wz�gS4`��a߹�}r�/~ܱ��c�grM���2y�_�A
)�C�׎����V]�g�pF�a�ͼ���@Y.Bз�S��z�@��>o��d�ð<O�;#�:�J���C��ʛ���)]h�z��*L>v����7ʌ��ow�>��Q8K1؋y:+�$�v�p��f1#�,��G����x��U�UR��s�(y����̴�A�6ˠ������Q�6�jN%�a�K�]3�[���3g���;��4�Ae�[��4]�L�
�����Ϡ$��K��/��Eo�S0�Hm����`�
	�K�&vB��b��,��6��Z(�&��ۚ(^��+ř��K oRwwξ�B�,�^K�ac�&��7�O�'� .����f�t�ңY3��'�=GLC$�l7�k�t��+�[���K����N+y�a��?I5תmձ����]�g�}*�(���ue����^�G�Q\��N�(�G6��ПDjջ�QN��bu���"�$W���뫒��5/��!���פ�o�9�ZU'���w�%��R��iB8�+B$�l'��6=����u���a�P�9�n���\"TS/�MmLj��F��>Ҽ܈�?KΎrj����,|j}��/��'�w��4GAr��1t�����gD�\�Gc�<v:Ǉ��|s ������I)��� W���E}��y0�ij�+�0J�h<�PR4;�N��c\�y�2�}u�N`�ѧ�~�'_�o"��J?ol%��ET6a�X��?f4�9��Z�`�PU�s�|�q�Z�6�Z����42il2�(� T�M��p���a�; ,Pn/��f���cui��D��U�w�5ʍ�2�xneFe�-v������d��zݎ$+K��S��RdU4g����f�/ʘVkD8_Π��;�0�a|���a��!W�j}AH"��Wi����5�(؂�
8-�Mlo��i�RKuJd��9[��$���N����5/*����	|+�ʔ��wN��^��l �bx�}z��<�.2�Z�q��ׁ&>ǭ�ř�_�Ƶ�oWQ���p;f�c�Ŵ��Y-'��Kh9Y�[r�I{q�&����<d�i,�u �c8�$�q���ŀ�T<}�(	T�9�T�E�T�!BgB����t Ěm�"�N�,��򸻲.T["���v�xO7B&m.��m�Z>�c�Z���M�yEe#�Z+���K�j��e���ZΜ��B�y�aF��))�=���1�1��(��{�)ݦU�.U� ���'ާ�B�NXz�w����-����΋���6��03��A�Q�'�eZa��sU�1���`�H��-�ȥ�at0�Ո25�g��E��2��
�M�`z�r	�dg����r��`�s�y�� 5����fRӃ
�ֿ!�u�̹�S�;_�J�x����a��J�+����'�d��d�����qo�閩���Y}�v����ۧ���P��i��a����nf��8��[�{Pj'`�㸇dǔ%�����"I� ���R��Υ��i�&N� x��q��KJ9%K4�*2:=�������������d��%l�?�����&@1�3�L�Y0��?̷����S6����8 F"��z�M���+Y�x R=a�~��q�g�?�4�INL��1�-��گ4c{���˘e��U>�dV�,b�"P+�6���ͧ ����Yg�T��������M�Y��W��Zm �-(�;]�6�w��4�௘��	��O���Y�3������k�:EX� �8���Q�fG��k*��3`�k����;Our�l�����;R�6\��5)@�E.J�]���+a��� ���c�4#A����_��� DH2�4*,9�u{h��$��Ζ7��!{'�'C��0=KCHE�@����B7V�%^K^���^����a1���@_��6��>�&��
R-���^�nW�;i_�)�;%����.r�s�'��i �y�k��\��q���b�����l�1� u�ŃV�^�h�Q�ף�0����c����Ϧ��`�Y}�@��
9Ǭe]�p�JX���9�y�a����z=�V�;��-
�eh����>x�c
���E�Á��=���J�$.`�UW�$����tq�xT�_��"�S?�T�z�B`p:��"B�c����l��\5�q��P��X(��P���ٿ��y�8�K8f��S��k�D#�A��1�<ԃ�K�)#�z���`�����}z��}tX�)"u;>�������0+�f=)7޵r��V�d��`8���XO�7k�"9���b�I���*f�7Ʒ0���o?�n(h�~�I��4�&T�X�����I�S�UNLh$� �-7*�E0:���>~.�u�ݳL�e>�_.���k�r��������QTE�6��=_����-z3�P!7`4�*=�vX���H��1W�����d�1^ǔ�C�:"ޮ��SKC��zC�%H��av�H�� I�T?�֯�*w�e���N����X����?3
a�C�ǜ�;�)��v��}y"�Z[��==�8塓�,E��m�ٯ�`g9IL��N�/�J����T��\k�M΂�n^/�R@��&�����8{5�/f��(���Jiy'�*�2kF���%Q�C�&c�8f�{�BsQ^N-�<��-d�Hf���M�7u�Z�.nf�	0�#:3}�L{�LՃ¶��ͻ����n��B�EJ�9�n��wI�o�?q�y�q��E0x��eo�$���Vn���i��E��3�U����";��/988�SIî�ޖX�5��pk���
�Yc] ԇ�*p(�� ��|���	�A���x�<�C������,,1�ϟ|���^m��]�����9N��}��?"۟/W� �Ԏ L�s96�(�O�fvKL��L�YV�V�\1���<���htT��=1����؀ϐ~��\��<,r���R�vg��zCAĽE[�����[k���	YDK`赢��v:��e��W��p���L���ѷ9oaTY��Ԍ�B� ��<�M��|��� pΎ�.H�'�:��4%`�L�� ��\n�H$�J��U��`�j���.����V (�y?|���Bkx��ϰ7�V�=��[�M���� g��Cԅ�ބ3��j���;,.�mV�-�!�N���L�ü�99m0�^`�q?7� �f�e͍��~�Z��.ǫ:gC���,��뮳�	ȗ4�W�@ş9����J��/�L���גCM�0�~�4�c�% �:h���TXe� nì#L(�{�9�^%�4���ho�
��[��L�,2�KOPdru��_@�%��*��Qq��t_�l5H��^��@߽��G��8��A.(��?���𡕤G90,oR�A�6�s~��_Ϋ�8S�Q�q�K��!�mZ�coGw���o{g`�ځ��z �&�of *�� qz��ׂ&�32ro�s�ñʑ���A���U���h�a��M�l��ͨ�u���7�7����}B�墭��W�`�zu77#}�X�-n�i< 0ܟ����\��릜������t�J�x� �VdOA���5�{S��~4s;��p��1Ou7�����h#h�-�i�
���9T�v[q%s �,��G���� ���=Η]J�ӛ:��k!�EXޤ'O`���g|�"3RS�H��m�۠,g,��-�+��:�%�FYP���{�@�����4"nѨ}�9�Xe��kh,<)g��g���{���%�����Uԭ�rMQ�8հ�6E��i]��7�P�T�;�C�ozb�s璧��tD��Ggi�+�`���H�q�p�Y���]���u����}s����!Y���l�fE���OD��Wz�4��O_BIa?�3-2�$��x�����%O���H���<X��q�A)�"+>�.��u���4�i0��A�ژ�gAw���0�fm���4��e*�g��$^H1����d}�]��EpI�_�d+8Lo�%m�?焐��^}E�O钯��Yr6��D�D+�q�%]�O�������������0��7,V�wvUM�� �@�gP��J�)>��W��+��wƙ�\1��:�ip/�M��x�ȅCo!���=(Q�i���^?��R\U��Rk���7+`��>=��͡�S@�������!;� Vo�L��d%�Kq�μYk����z��2ٹ��op���2�W��C��}��^��?ٞ�����d�W������$�,z�,�2�1x{��cx5��qK���l+��_h�32�ةT�����S��］釙�c���w�0����"�MԜ#i��.���-�$Vla�q�wn�1�8kg�@�H�f��r'I�1��-���7o���	���m/� %� y�r�p��8��M�3x�' �8=���sj0����|#��:�өy�+��,�Q<�h�O臝�ܥraH�lQ0�"�N�R�eV˭e6qP0�3��5�H��4���t��i�N��\���a�~��]��j%��}�ߐ�.Pa���8E�+5�J��|�ZâęFĲ�(�G�D�-ZZ��G�t����h��v�V	'��著���ԝN�X��⺸��k{"�1aNO���E�B�]����9X�6�Շ(����)������vr>_�����A]�Z����Þ�e�Z��W(#]X�03?Ο�y c���mZCD@'�?�SP�!�;Y����쫆��R<�A�x�E���&�פ�_^?��T`֟�,��g	�� �&	�|�g6�H(�� A>v�!�A�G
��׭*=c�6��ש��!�?/�1�Ǹ�v�eQ؟��)WÒ)I�����\��(�ÀR�-�з�3�(��<���xfP
iyvCP��3\T��ư��:�q��1�s�JC���$��H�,��_T4�+����� O����=S�u�@Ĝb)�q��Ir��%L���~����zc)�m��Xo�6�N��?+`#R.Ό}Oa����5���H���qJ��0�K �v�ͯ[���OQ��;l��{��Lb:�K� J\s6����5��Ss���3\շ1��=Ь��hce���D��M̪$>.�"_�m�i����,p��5),5UU�*&0</lP���.~�Zݒ� �n�����0vR�m$����g�U(*��tɠo
X�t38;}���0�S�1�	_~��\���S��҉�����3f�����&��7p��!S0�֟������5V�W�:���7Gb�ކm:q�R��ֳ,����%�S�?pCS��-.8�y\�%�|��+y�d;�ޒy�p�)IhQ�qFO���d�.(B|{�>�2�V�V1�a�d|�<��8d����c���"��0�D7��v����r�������ȇrgc�h�z_�O�񟆑�כ�!4��x���s	^�7�ӖF�2v� �v^�B��� _{U��ꧨ��QR��^�L�,S_�Q|��L%��$E��?U���2���*���',�Kx0��m�;~�q%H.P-ħ4Ȼ3J���֦�V������>��
G{�L6�����m��C�U@��y��1% �'c��ck��Ǽ�R,�H�u7��ZIc�l����N������0ؚ��^:���l"{>E��P��]C������rA��d�w)6Ur5� 
���8��d�mڋI�V2�#\d'̔%R�4r�ӷ<����֙Cu@�� A����ځ�+;B�h��J �qI&O�k��=+����\(o|�`��B��玭fQ����>��Eȡ�2ӡ:k��\�E��W�A&��g�7�Yn���?��X��{��}�:t6��������s�����L��u����p��0�%�#$h)�]�)�x��9�J0�w���"�b��umPh7����9��>w�f�^�m�+���	f	���^�]r��K��l�_1����7׊A����L��D��06��z@��lb������R܂(��,S�׳E D�G��ݨ�9���42��S͢
��e;�߄�,>�Л�d7 $�q�pt�y#��a^o�r�gR
#�#af��|� 3'�J�S"�r¡K��]J�WE�
���ʏ�ݚ�j���a�lz>�"h��fN����:� �+l���3:�<�ş�L�w�ŏ�7�L�H]�*��e�� ��%'�QDA��xo����Z�O��&�;��MB�le�Y���� ��DY^4M��}#V���3�t���f!Rc��r2���WS?����`���U��h�gG�m�i+>bh4먧�H�g�<�y �v�x�5KJG��N��)~k���X{3���(��=Ȇ�bS���VE�j5�M��_\R΍���<�Z�e�*�E��($FB�ш�5!��L���9w�D[Q�j��5�i�6́d	��]TV�2]�="H�r��%6���/�u!)7(���+W�2Z�9���('�8'2����j��ֲI��w�`�,g�H�0���A[!g9El�z$�Y	S�>e4����w�;�Aחu9��ԣ1B��=M$#��� ���߻f�����DI�dw:��Z& �Y@�hT�k��dU
Q�e��L�$�A	F��ZG_�M����;D�;A{5���j�n�q���Q�y@Xp��-BU��+ �k���ӟVﶚ@_#�y���$YV2p�Iu���i���"�S�����9������O�8�@��pf·�j��?���qL$�z�����X�r*�_j�v�~�0��oq˧Vf뗍�qJ�]�ǻ��;f�2!�1��j�'�H���!I��ut��1��ܳ�OTK��7c�9�g�rD�ݠp���5_�qb>i�pD�x�t��m��x��3�3�_�&+.
g0PA'���,gٹ�Ab�6��[��UC1y[��v$�����gX/�Ş��%c*w/NŒLR=d��f-��&�賜�W\�÷���~�V�~�N@_���WS���5ŷ>�������Ȋ��-�s��lnN�)�r[��
+�2f:S��V`��61�0��F3��]�S��'���it�Q��g/��L���M��A^l�O�s�b7���x�$_\j(O����Nh��3��(�&A�틃��z��nkqG�*&fEJ����ɾ_�nX�T`��v�� ҿ"<rě�";�32N�N�8H�������V}ܠ�n�_dT-�e{%�"j�v�N?��_�	�K�lz��i��
U���/���	fj'2���@�+L�:���	��2�&���5?&�4�B�WZ�'��/D� �Ht-���fv�bG�ko���\w�C� ��j��[3�F!&�>��V9#�5_��{�*��/��Jz�CE�����W���YT���A���wq�M.UX��b�I�v���Vi8C �%��.�N���?Cl�G@�]x0g���ǡ���Vǰ<dUl����4��:���8t��6��T[�.�Yj#��+~���wM�r��W��ۑ����#���:��hg���D��p��yH���ܔ��՝�����Qr𞔥�w,��I�CҔR�����B�*E��'�<p��_�>��i�H���ʃ�zB��Xϟ}�C���p`b�2
+� ]G�]G�b��#�-q#���3 ���ե��w���q���杜�镨�d��r`��Hn����$j(<[�fAz�k��ֹ�!!4 EJ�$rT^!,K������go^*ݚ��.́�̔=7zn�9X�A�C|!�{R�`���u9�и����$BJ�6�c��6���ډ���)�%8T��'�>3uڨ,j�˲�#Ѝr.hq�gy�@�[N�m2m�єk׬� �.�kĔ�dH�b�QG���P
���A�so��?8聧c������_�
Eh
����``-Y��C��T���d���ѝP��x7�����)<[2k���0)P}��ӑ�{-�8N�ފ��ɷ�Oԫx���� ��a�����J��R��ό����.�(�O�/%I�r�f!]�T�3��w1\N��[���R��
Ӈ�nwEZ1J� ���ۀq�q+���vvc�G`6��(�j?�̳	�X,QR=�d�]�F�
�X6n��V����/���4)���d\qƐ���Η��Up�_�Ld��<M8�݆��jz�vi�Ԇo��,��i  ���hμP�������_��O�x�J�n��	O��Cw���֞�M���xx�qpu��w��'��$?{j�eS������9h~�wi�p���'�1;��Y�>Iީ
_&f/�:��* }���jk�ƍ��fj���	d�N �(�wFq�2��<\����!b%�p>�F^���&���Aj/�r OR�%{��*�-j+	����imk�Q���01[�KWZ[�!ͺِd����v�U���sV��l�g�g����(;m�j�����IS���<��P&�V��3�%�z�a���_���*�<8���]��k.v��d�)F0,�T��Y,Ȃ�=S�q��̏P�x��Y�5�=���6�rܫ��:��^6)w��DJ.���vIH�{{��K�.U`�����1��Bu�z?� f=�̘�ش��u�(;����1��NS��\�B��!'���r6�(�̓B����2L�bw{��	���0އ�V,����TW+dX��lc�������2�L/��:�)����Kl����[�C���s��4��C��Eh��X��e��L�GGZ��iy'�6.���%�{G��ǥ��#~����I#��~����$3o
���ɰ��r�-(�r�t�Z�0/��|n��|?�2WU�RM���<��ϸ�S���A�y+���ӊo�Id��{��ynv�����'��ߴH�����o����ovp��c�=����1��-� ΓZjĶ��x�	���E�[�
ٝ���Q&n�Q9+��+A�Y�����{Te�\t��4�Mհ&�?B1
\��j1��n3�uYmoJ
�C�aȾ!a�7���#�
��&b��%� z;C0<���� �"���~��[gm�|�'^2���ՔU԰\xK69�=N��s�m#�j���*�����!�cm~�R��"M��oł��cq"�nnM~�C-����Y���ǝeUDa���
%��M��`FƇ���($!�%�n%d�*�T���0Td���!���bA�~��}���қ��?�[��
CQ��KbI�TS�FD�RKXCܧ�Q4�cr:	�m͘AR�������̰���ä���L����C"^N��L��R�x�O�G��k(��`ܺ8���Ƿ��\�"���w�v��{Pnޫ�"�V_|,��C_d�
[@m'�O�q�s��D����)�j�BLl��c�hj	�5�M�d���$�-��TԎ��U#����w,�D�����y�}��8
�����_,��8���ϫ�0�C��#�틝*Q�&a��i����`��H�f�ϑ骜��Lʷ���
?��\�D]=��(�X�W��C,�����
S?���V��	g�)/:Z���B�)�>ě�n�WX�`�NNN�)�������]�4�X�&�i9�Ia�<���@��󟣖�����;1��!0�Ia����.ˆt2�93=�F|���B�O�]m���NL�c�\����F�'5��(��Ќ�+����9&���&�i���5���O�.�|59�>��Kޑ�</�W� �N�~m�^�9_�a,�1�mH*UЮ`DXavh��cr�)3믄��粜G�##�q+�������r@Q�\�u�=̄2��'�9�� ݶ�5C��Z�0���eeL�@Œ��5�q��ץئ��Ex7��K�<|��l����=�G��Ԣ�7y.0���!��bH&\��&��uJ�~�)ň��x��3�)I�]�!x�ɘ��y�Z���J��TzK�qS�����]�D�
��H�t��_����)K yh$}�%���P%+�:��FF�M[EP�mf?R��["�0.�q2�]�L�9�I��CEGP�+sVP��y��W/a+�7�`�4_�c7.q���a�aZ=���3��s��_Ǭ�eGb�S�ó�O�K����k|�{am���a�d�<�?�GnpY 5y����W9v����Tߟ%SH���탉��ޤL����'k�O�	�<�M^$���mP��Z�HǠ��D&"2�_���mvL�@��6q��~:� Lo��2��v��r{������m��!H�_��n���Ŧ�v}Oɭ{��`O�c���Ҝx,�9�[-�R�$��k�ը�j����$(��[2��$��#�#鐁U9�HA�8���/��P�`�3�s���&�mW4T�C��ݏ�T�.\~�f�r1�G�
�q�B~lL9�W,��mMQ� ���j�O2}�T��[Wq�������
���B���p����1>[We��𽣌<�&�f�tӆ��k겸,�P�a�QV��j1: ���$r���bb�@NK����K ($����6�m͍_�3j:N=wSg��s3����D֥�r���HV��%��F(�<�m]�&RF�����PQ����X�|�k5]����6��<�i�����}I�զ��f+��'!E�V��<gv4b<��ٿ5e���/]L(�k��a��v�^����gZķ�������ɷш��?}� ����Zo 2��[��Ʀ	�LZ�,m�5֑"�o@l���k��y�B�u,�.a�{�
��~o]��N��2��������k;��j��54�I�^��N��^����JQy+u>8�uڣz~�Q�a_�꿆*_��k9;<�3�߭d�(l�m�A��	Y�`��	Lt��&�{<������͑�N�d�`q�R�t�p��6{�.�Z�����K�X.���W��R����?.7f=�>�g@�M�ŏf�WP�ρ�đ�+�o�_{k51U��mrN�c6�O�$�%��d�f1�ɱ� ���WN�{�h��!ƪ�_a�=��� 6�M��tp����@��V=|j�����0�ڎ�D7�'��_���6��d��.�X=�${�n�9�~z�b|��$<��&$>aǓ_����E�-��h�X��� �G���tPٺo�h�(���v/����!�w��|ި��O���|
������-	!��H|UXB�O���=��b�2��Cm�����yN�2�l����,�SEgT�rJ<��������wյYXǃ?�,"">�mJ�Z���$U���:R��N.�)#'|Z4d)IUxM��E4���Yy`9zI�SUZq0D�֖pFjn������r?���� ���
[���?�<�XJ���C��|5��yH��c[F��4�mk��JZ���뒦FY���6��n{��C��T���?�l<�I�Jp0|/���h��G�2���g�S.Xht�ݛbj_�)��&5
��h>[o�6�7���8ܾm��ܽ?�*�ZUӍ�����-F{����I=�Z��Z�n'𥡗i\��f�SuIg�x��Q�f�!�q��r2��X8�ă��5K)k�9���)����
��0���|.�a�TBek���+@���QzbZ�\q'e,��5b�l:�[I-7�(����ம*f߽���יd���V.�8����Si��6$M��	N�$�DGA�x$��KBu�49�{��q�I?�- \K�Z,��x�a}n�5Y�R$AҒ~�vɭ��������4\�c��Cl���rq���H�	h����!�2fWSL[ːie1$Y^�'ǁ8[ԌO�]�
�X���}t�Q�v�=�>�E��F��5�W���)a���� sIC��Q|�so>sRZ��N�Z}�����o�����0Ϟ�·G�1/J��k��p$���l��А�Ăy��	NǕ�[�!�@�=���O��g.A��SK莊0��xZ��}�s��j��j��ُj��^dr�1�n���z]	<��3VC��S��0��oe�W{��9)��n��Yu}��k8wZ�qELlY'�X���*��$́K|⋜�|c���Ѿ0�\7ÐN�����<Z��}�"0���x� 䩋��Z����ʺ3
{hN�ބieq��mAa�1{8��9�qL4�:�C�ih1�*�4�E|yz�>o`�UA|J	��ʾ��`*�#�b���3İ&ņ�w�.�C�L�GӾ���\�U����j�&=ϙ��-8(h��R�*�B��+�I�8 ���&��P�L�߰7�xl@�'�@�A�+CUp�CH��^�WΪ�OQ�O��c�%S���y�k�t���YX�<��E�?л���l����'<�
�Lc]X&=(�x9Ur��5\	����l9��&��V�7?������<A�wb�Cr����$6A��0�6� :I.��}"�I�=�Z/�}iUӊ6���MI�&�;��u���òB�A�UɱK���V=S����}K��n�PY�
;�R�Hm��R=��ik�G�B���.��8������2��*#�&�\���q�B
X$g��;IXh !i{CLE �����J��P�%V���sv��X#{�+�I�T��T'�l����g�^J���\ZT���:�c5Ah�3Af�VB^����X=��؃�:����)t܆������h��>�?��&���Ǧ/'Iʴ�+Md�
��Aׅ���TV`�B�VJ#g�dm�g�n\���0�b#0TT/����e|%l��A#%���������@���`<36xt/"#�!�|�M�%��	��M�&y���_Ȧ�7�`��9'��Z���snT2��D��S=ş;U7�V~C�|�}��>v�/˸�ԧB>��N��l�{�J �k"s�d̷�V��]r%�~ƨ1���qL��$*?H��1 ��ڥ�����G�h������02"�<��[^��qXOYwY�>�^�>��*[�=��Z�a:a\�6�.�Ƴ4���ɽ���H��8n��6�q�&�E���0��#��i�>����N�{	ji�+�n���6O|?�w�:��SH��1j�t_���Y��Rheye�������Bs�ɥ�3�+�i�	��X��k:����Ļ��Y���z�r`m��'�5�R5<����������í����e�J=2��ܴ�з�L�^�IIw(� O���=�lZf:�)�A�dg�
.͡Cdl�(T6��803r���i�|��/l�p�C#�����7�z�x��o=Fи����G3���p�h�8b�9�q�9�]��q������z��3L��m* wO?��t\�A��Co�͆������[}�u����y=|r��y�3�����k��<��W�M�1��F4emP���R_-�������a����B���/B��Z��$����]j�����Xu)Fǹ�q�7i��Sҙ��K�Ϋ����u� �(�.�t�3��;�h��?�m�F</��
F��&
�$�}��/�U�S��N}�:z�����[��A(���v}j�`K݁�p1&���ϖ��Z��9@9�"=���d���� ��hl�}pp���$�Bi<�	s����ޤ�S�lh����Y�;L�*@8cP������R![󋳉f��(x�)O�5�����o/h_~� >21�ծ�e;�d�D�l�^�������v���X76�S���I�
�Տ����FVU_!e?�=v�����PFֵǥ
�� ��0Е���#=YxH��eGNo�:Ʉ�_LRA�O��)�8��Z�J��dٚ��(3i�UqY�����ލ��:v�,��t�(kxI`����n�6��3--�Ӱ�;Ǔ�uuW�N��pė�.1<R��J�	�����q~rǒ^"���c�x��tA����֟�Aa
zN�p-�D������y�s[� [?K���c�����	<�l�؊�m1��g��/���`+���]��t��]�֜O���G�-FT2TY��/��Z�1�że�W�.FAR@O c��֦U�H���/άtü� �x{��bh��=a� ��iQ�Hڭ*�f���zS����iܔO�䳍��=j~�jg��4q�)�0�3�;� ?�_�1L�X����S-��4����M�ڭ�C=Y��i��3`P�jJ���U�w�2OOh����7��R%�-��s8�,D��e��X��*5�A�A����g}��L�F��S��ɍ�b+������	F\�� �l�����u����V	�R����
 �������4O"���w-�͋j
 �C󷶂� ;fu��?��k1InnP�a5!�\'Yo��_��3��+�	F��a�]��H�������⃰,CP��Ѡ���'��,w��S��ߒ�F=�/eߕ{���! �G��,a ��)�D��������١ӎ���i���' CE�k�O�/��}}g��fD�@Tł��JY���E2�
jM����oӟ�&��-8(�����4�Ú�UЮ&����>l1h�Q�j!ag��:�_F��p=י�}��
.2���ژ�匔�_+$R���68�s��p��'�:ƅ��NU����EΓE��W���(��# 1M�P}4\{�!\?Y�^�%�.�u�&��u��˽�M(�x��5���}߳�M�y�S��	q��`�0`���H�jUَ��Q��@R�iM���M�Ho.$�~4Z�L,:���C�C�<�\��}]���K{�E%K���R��9q鼯d�����k&�ےRc�����[J��=��Z�(��F��>W�U�U���T	�w�J�s ���qs��uN��w=!	|���[[~��|-�*hn[���d������X`n{�o���#^�U�As���OY�O$G;�#&�3(�Zsi��a�S�06b�ᦡy��R6Ʒ�����ɣ�p*%s�>�X�
�2�n���v�k^��i�ȑ9��2���N_��E�"1��\$�4�|�Z�D8�fɗ�ׯ8�,s��2��f*��������f��j������0������AGVʝ�+䪸� MpUԑ���S�)l� rPm3����L�1q�G9pw}d�L���?�F�gaE�d�6xXF���7_��,7}|����R���Di� ��M��y:�jԋ�ƣ�ӛ�xQ��9���o*r.���?�����\+x3�@�V�9r�|�.��(ΰ���-$��<�g=�������5��["�i���Ԑs�U�aN]&��._h*��%БDd��+��Yb�/���+�
�AoO��.|:�.��=愤�P3�q��$m1M
Ryr;�0Z���a�A���;���cQ����C��LuI�|f���'��7�]Ρ�\���H�\�Ua�Wj�]��ވ8!���p1}��eNW�?;�Vh��=�@�4�P���\Hv�%�M�ҩ���Svl����=�2�!�LχԼ{b��?���G_��U�>��Y��3bJ���'�5�\�r�d��Р�H�}����W��B�~�7D�x�_����=��C۰� ����Ś��a9�:��
rw��zUKF㇐8x���S�f�C� nΉ�s%&�����������f��UMD���.���2 A��]s��י�Q�)x��va|����'�˛o����\�C�8�JM\�C��k?7��WS���`9.tI��_Nk�	�ڒ
(�]���au{�;PVv�f��ԙ����P�1=��ݠ]�G�he��Vdck.j��~L��]��)!B&C�����]�"#`�僇�ޮ�=�������`�0�m%t[�'E��Z��R��� �QeSk��*`tC,đ�rU�0U�tο^����� GZ(��Hu�o�
!�T�+(]A�E�j���Q�iq����˲�;�AqMʓ�3����)�z��Ӥ��)8ZDOB�)M�~�(��O`7�-N����W`D��=OH�sWWF���52:��o��+�w�������~~�5iI��ܥ�4+��{���!y�4#@ �'��~�w��|=��ﻣ��,�تM�%+�-��X�<����@�H~Y����LQ*��4T]p�ZX�=�%��|�M��q U�ۍ�sL�ޕ���O㯺`�Ӊ���'L.����qA�l��l�ėI����PrE��~���5�$�(�j�"�����~�+�'R��%�:Ig/l�� a+'K�7-vD��bO��L��~�_j���}�di2�2�"	��(b��.}�B�X!�O��=�y�A��b��^����a!�Y�:T�_\��pz�1z��ogFr)
[]��鱜ao�D&���s��+d/tMR-�!���Q\�O�P�*^|��sb��6�������J8�7Iy����� �(<q�"f�t������X����9_�b�sn�@��`�XC�a.)���%�� ]�z��N��?�҂�1�@����#��i��_ya�pZ�سcI\�C�"`���� ����2��*5����A'5��GU�1���g%���	�yM.�T��\�<\�q���2LB�@]��En'tE=6����2/Q�����y�&�=���l��5;��t��dH��E�e��Ԕ�o���*�M�L�����u�R��/���9�ͺ���� ������_���|3�!Y}�
֔<��]|�
6�PK�%Ho'�I?xMfc��e`�R��L�{�n�W�������a�|[��{��)r�r�Ӭ?�3S{\T��X�Y��T���a;�����Q�*y��g���D��0�i
�5��@7�I���/;�U�%Py9ysy���5ܵ4�"������)�<�$��
S���S�+�<w+a?{�~3���ڛml��#h��lL���滽{��whz.�z�,^^m�6�.J] 6�a���hB�㣢1�M���6J�(�FT&q7�Zp�5�pr\����S��'+{XM)l��� �ps���FUB����?Y A`q����SR���'�7=����<?�Ҕ�F���l^�`��u�|���aTAU�V�ݐ.�0B�W�Ҥ\�	�ݠ�T��s�{T�M@��NP���п[X5(��Ǉ�P���M�"�Q��(C�
Q(���<F��)�LP�գ���)�9��)@A��+|;�N���޳��"�1makK~0�39G�/�
���;"�S;�HB�6|��p�]�ΐ�G�1����x�n�"�����t�1o�M�m�r�owg�<�Y谺5�/�:���3Im�.f�Q.�1�ع��k�BL���ŉخ��^�W%��[�����s�s�r�+B*���.U=��H��{�n�i��=��ɲڠS�z���M0�Ψ�[X��h̻wl0�}r�W��ژ�m����Z�I��:��2�2�t�"�F-��ETqf�U�&�q_̒d�R$Q%6�2��9CuO0�F���&��A��C4E�dGe�����ح�*������߂�oS+��{��Ǣ�v��$Bm˄@�a������Ԙ��Z�O��E��Ih��g�a-p�~.�O�t�"�g��n�?U+ߊ�8���Z?+�#ר���(¿M�Ar�'|�߶U<�j�2"孠�������C�_s��t��퇎~*\E�:���Lk�w��r��c��ā�`�ߏ�.y�#������֯�-PԘIU����f���������t$�u���i�x�C�E����.���~
��
m��Y�?] ��"�&�w�e9\Ɩ��/c�������I�"kGqX����TqѾ�	\,Ox�S��;�	�e:~z ]�\���>���WS�xqU͓*Z1*:�)��(r�%S���B������P�{]Ò�xg7��7�A�Y������{��`�#߇9]q��2ء�:��#Z���������4������!�}*@��#hMq�Ė�!�>�} Az�ρ�$�瘥�"�s����O֐��4{/f��9��E!�2�B(A��A��b=���e�]��H��$�O���\.�-��d��s��$_\J�D"�9݉"���{����B+�k3���c�U���ζG���K�v��L)�ȍUO$�
����h�J	�fK<~5�R��]��a�@�f�z����T����ڇ��h�M�)��&��w��?0���r�D9}ݐ��?���U��1`�dn�8�ӵ	���?�.q������TRߴ3�иs��`[�AH���Ȇ|���f��4y��kpk�ݰNф���PsP�ٓ��+����-q�	���A��L��J���ՌR��u�:��j*�d���e�}]�3��y���G!4tc���p�s�D	}�Y��s�eW�y���Y�/��TIظ�T�6��:Ä�#��;���lE�Eh�t= 9��}�j6�!�v���<���%�@�bX����e�V;�!6��h8�<̮Wǉ�3`s��U���w{W|�-P��=\�B"���V��U����l̞�X�#�Q�F�,��$�K"Ąa���� ��fXZ����x�2�/2K�^8��X3��*7�
�⌦G�@�~�/���oUp�J̏R�,����A0$,6�WM��n�ti�f����'�0��]���5�TEHh��٦Ep�#�UL5�����Wg���^\Aao|v��K���Ʊ>�L!5Q��}P`�w�q�_`M!���q���Jo�ڽ���F��wP}�=<[�<r�aj�v�5o�Ӊ@\g
2[��8㿬���wU/U�3`�����72�MbD�%���\�%p���,�V���cF�w��A'�&�DԀ惭�W���y4��dc�-���v���!r���@r��UY�����e�;Q�oXh�u��3y�*�����hh�>L�WjR�Bk���c�ƽT��PK��i�2�n�$����v�����vA]vT�h0qG�tB�PK��g;1�����o�>����?�Y�* ���� X7��э{�jM�\l�q���q���rQWx�.�½î:=z�RXG�<Ry���qa��I��ÿ��!&�����!�[���\�A�=K[p[d�&�T��;�ɭ�:.���_t�i�x���;�����uU�_�ޕ-+0���!�/��:���M���I�:[������HI�J��A�0�={�rkl~V9-(���!b*��4���|©�4y����'�I���ɔa��������[C4@(�ؙG�B���Kߌܧ�3���V�L���f5VY,*�-F`��"��o8ΥMZ㲀�)z�iEGV�b�QS���B�@&�|�t�փ�ω�UBxfdoV�0�����&ʧ!=)z�����^�YE�y�<*�{>6:+���s?uk'��ũ:,C�H�N`��ֶ�Mˣtgw�o���c��v!r3
��O��3���f(F��Й�������tnD7�r�GM������������� B�9�G���٠��0`�2�^�����³��n�wJ�\5c�E�S��^���i���)��(Joe�5�XЋ���q,��Kk�}�Qjv�'U�`R!e�4� �'u�5��X8�E���78�Q͟Vx`�yU,z�� ������$͙'�<������as?�{$�틘�G�a٥��~�N޽��-���,���&���=_��,R�M�5�!@i�^[2s<�E
'S2�ײgA���N��k{-��~�y�Ѽ?���xuSL�R������c$�����Ս��i�{�`\�_�g/ymǰ҄�P�et * �&FozΙ߭R��8m���֞�5/'084��~?L��;|]�HwwAkF�=�9	���b P�T��hh!/��e��A�!�4�-���B��M�V`gcc������$ �$��=�q'=�7\�e�;~��Y��c&�6-�b�rc���/k�㨽/`�؊K���>J��Gl��W�c�3��"&J��T��M����+z�9`J%�UI��:�4̝�S�p:�J?Z:�y������۫�������R�_�m6�w�0H1�
�,;UTUS����]:x�2�ȡz��O���6ҏP!y�YQ����9�P��9 �,�4�*���!B�&-ɣo+���}=�8|g#`o�[-`t,?B�Bm�1����t6u��`�DXX�4U:)�� D0:i��<V�#�)���F��K{^w�Y�|�R����D�C!L��G�T�[{_�>>,���C�_�XJQX��M���,
GK@Z�x�Y>~�/.[@F���Y�2�pԧcll]�T4����E�@F��g�P�.an���ߥ�kO1A	r�7*���-L&M���m�P��< �M��]����_�ս��9N6�ў����O"�mG��N,�(]�]Ű2��UN�؟)�%
#oqF�s�{銝r��O�G�t!�Rx�i��V?��*D���v>����E��ޏp�������nC��N��Ȋ30/��{��]�V�N4�fڄ�f+�h��}�ʛ�ǠӺ�Q����b�ŀq���(�}ǣ��)0pr���D1G���*�hq�mY	�p���N��Xu�^<[w+0G�
��|΍�f����q�����ۆ���gL$I���7v�;S�⚣���{P�aCzV�EQ�
�֙j�+��
��u@��f<��s��+s;�Y��iH\*%5W�!�~H�d��<u� 9������u�E��꺜�:�6��T��z�������'F%�(?x30��f�$p�$��p�bLu�g�BQ��  mǒ�'��<�����UK��XK+�˽[��2���׉b���h�;�����Xr��z$��+|��}��E�纺��p4x?x�t8n��޹��=z�OW��B�/���Y߳�ҷl��@LR������j���e�������W�D�D���!Ӕ�+��-�����S�! Zh矜����Q���-�ܚM5�X�X�����J���ǉ3lS{#�@�_�iM�xwЫ��y��A����+6w�ה^yG���XZ�=O���Fh�qC�x�f�5���+�Ѐo�B_��o���K᱖LO��g��|����� BRN��+%7��b����k���}��yAG&�V�<�O���s���0Yq�H�C��b������^9�h͒&����;ƈ���vO zs%
�!�%銄e����c����^��u�-��YS=�Ym��M��N]������{ߣD?��@w����
y������+�;���{�|ŔB�ߥX�)���Ы��K	�1�Jv��ُj^r���������?D��fydx�Z��)@C}Q�YHغ�*��6L�����7��>A����$i�u*��%rMXa����q�d�K���`'L�xB�_���D~��UI�ӭ)���Н&=���Ոq,d�QQF�P�?�����I3#����x��8b�˞�v��3�����Pȋ������r��^g]x�c������-t���L8��[]&�n�C;������<��OC4�\��.�؝?z�I��~�(]�s��Vj4Y�@t�V r��(q`�r#��-�Ϛ�M�i��qtk�Pjk-��e�.�_-�w�U��h�}glL�i^�k���3�	U�bj*� �-�ӷ1��%��؎��=
U�pM���bk�}Y����K�~�xR�M�t��o���zB�^E�y��,߇�Xʖ�n_���BE���C�&���z����p��C��Bu��s�" ��bʂ(?&��l����F}!�=�6��tg(��jU���4ϡ� ��k���D�x�NSY꩟S!���۵
|O����'y���h��	>�Ռ$Z3�]�)��fΐ
B�:y<�0k���gݞ<G��A��Uקj�ߧ��8��G	��Zͅف���#�|*����i���[�aϟ�2d�)�4�����fh�.u���`���^�F	�~�
���B�\3i{���Tt�$��o�#)�;�hWbȎ�+e��cj]���Ql���4F�A���Ŕ�����L4�\Ʒ�U�����ׅ.�Ӯ����}��(
	��n>jy=��4��b˚ܵ��[�}�~a^���no]����ؤ�>�B����t�pG���C-P���?��=ls:��79��{?���w�?���~;�DV/�J���,�J̱�.M�sb�����E:��q�6'AE~㒵J���Ys;1�sT�Pg��k����ӂ^����#�S|��QJx=���mhN����n^^��M��E����3i����12�M!�0z9ʧ��k��p�hD)�Y8���:�O�3@���a�<�����p|bkz�����VjO�Ê3?���֫��!|�p�&�܋tᩓ�Oǆ蠊��F�Ⱥڡ9�a�f*������](l΋Jv�Ѥ�~�T	$��q׹0�g�%m�} ��14NR��gX��¡k��-?"Q����j�t��O�h=$�HK�\�{�/K7�@�"�m�f_r�Av���x��jwG!c�wD["%z��JX"�=�a�����C�w�����s�ѓ�=��%Ɔ��U���~ �lg�u��7T�&��]�K&\C� ��HxȢ�L�訶+�_$�}_��c$��&=����F6x�BIv�[5�.R)޹��!!q��|�*m����"��CV0^�/̿bKVl�ס;�2�����!-�MU�����&�*N��"��%gP@�	�3j ��O���&�5q�А��e��J&�$��M�?��AK��r���-)�ǻAD� 9�"Ux�c6�o�\�S^o�T���o�gi٦X[Ũ:�1K�4���W������{E�u�6Y�#����s6��{@=��W�����W�����L��Gp�^ ��*���X)}����T�m A���R���W�0��>e�K�p	����Z֜��M�$.M��k�M�C�P�z�L�$X
oI���Q�#��=o�u�X0�<�F%�LZ|������f&f��`�+U���lȂ��3�� X�jv�p0�\��n��\k��le0�h����G`'���,�d�3���wj�����
�Y_��qZP�it`S��ܒO:Ǘk����;��-c�<'�7��2����׿0�H�G���V�t��T�7]�,��,!~��%੽+VD���n��漶 �$��/y� ��<���X*p��Ojl�,re(�Q�k��^�*QNA����[�n}u��`����$�ݡM ��:�GIwb|w�o�g�ʦ"�ٞ�~�9&%�7BGw�{��|����v(��Td�K�=�k������C8t���NDI��7�����7��%����Ş嫽��O ,Ęꤔe�?���4�y���u(�	�@��h)�J�z�-�!�T���ǫ�Ƒ��_��K�y �2�Aѯ��S�B�0��]tMN��N�`�XR�㦞���m����ǯ��8�(R]�����F� bX>������r�>��X��q%o�N���/�����I.Ќ���?&���9X��S��]A����ȋ�7R�����Dwc�FPI�f��~��"1����E������G��G��g�'�2{�sUy����i��fʵ�]�/f��(ǐb�\��b^h_`3��AI��ܺ?
.�P���F
LQ_d�U�q�T^�)� �� {|1֐���\�׮��ԀCI^����>�l*���O�)��[T:�R��"r����g��/�����?7�n��ŝ��:ř������ȝJ����[��*#����%�G�贗B��آ*���tH��G�cC���Z�,��֛�w����PUq����F�=d�i�s�B������a�|F�l�z�:�4���I-��P9C���l{�?�H/`WYp�VJhC$�o���f?�-IH�\_�>�jj�1J4q]6\���B����\��M����]e!u�&���0��2��lQ@ź�@�6�TW���١cO��g��6����֊t�ʮ{3�k�G��x�p]�'*ck����a7��e�-#�6�B7�JhǿYLq!:��&����A�
���
@���0
U����ē�0/H�Yߙr�7�8����;��dʁ1�}�����&u��,����%�r��F�㨻�k����������lT~�n@-��\���V��&���
����I��p�W��N�<�R���5��O��~<H�`���j����*�;���|P�́��FP�(V:2�
��6�;��S'a�j���8�I�.�pp����qI�]�I_��+��uUEm9�x���7�Y�ߨJn�la�>�N�c��wC�%�Ad��B�M\��H�I�� ɭ��6���o��� e�!Պڅٍ-���0=�F��-=�X��o3��hk���D"`V��$�񏌉��/���i/fI��:�2S$,'i����U�䳳�,:\:P~�"fnE*�X���͇��}��V�^`=Pn^o�&q�:j|���%�`GP��:s&)�;e��*�OaT�����U(���&J�1������6ռ��=�[�= #���c�����9��H��[�H`B����m�����k�5�듦d� �a���|'�E��I����� 	�+�����1�r�4{�~��c�IF�f�:�cۏ��T�,��	
��3	�d��oeZ��]��}�v"�د���^���'l4�W?U�gW�̯RF1Э�l��]��Rb�{M�u�6U�3����~����#����JN����Z���`�O�������\i�k���=��؋)AB�4�䊞�T(ގq�������3����|�=���g�2F�q����؍��bcth�YJ���	W,|c*/L�y�ʵ���
nЗ��E)������;.���s汸�"�r�7y�ڛJ׺2��M�o���HP�=W`�O������)gn�{�6^��v����<�`8�T9�)+�|bZ��M�wȥ��X��c�i�?;/`��Xc�hQ�Q5�k�r��O#�P=���|<�"Z/#�7���JnI�0IK���E[�ꆲ$a�����@���"�(��[>Q1zd�ʖ�@�{�Vf�'���u�<�����+��L�( A�<y˗�=d�����l�7�^g����:;j�VJ	��&��o� �ˢwxo���a���R�PJhD��;��sV��gf)C`���@K����	��2�^�lR�
3���No/v7:��>�5&��rت��r.C�fcL�B��N�M��
��ǒ;��:��N�>/�����L�kn*�£Y���4)c��>�;��D�˺�*?ncU�aܖ���X�c�o�K%ӻHkR�)�i�?:�����E��kg��F�g��[W�K�\}aJ��!6�E��*��*�lɭ���DA(�����O}�͗�B����'f�8 �Oe���}���������P�	�ޖb�ҡ
C+\�{�d�W���u� ���w����AxJۇ,�I���k��Z��Q=ZF���X��&�7�;ʷ�R}�p�#�����`�3�
�װ���dᡀƘ�	g��[� |�Rj}EH�T���2omm�Rtyf��x��|u�5e�0֢J}��b8���h�[�n`�lO��?�"�~"١�'+  �m���i���/,L���P��C*�� ݻ��D�����,����50!�]]$KI�N���V�%N�#{���=�uR����y@�b��ճ���GUA����)���)�),�՞T��~6Uyc�~Y��T�+��P�hBS��ӴEU2�o��A��,�bS8ذIަ���>3���0��Ջ�s퀋Ev�� ��JW*肤L�5�:�_l�3GҶ�PxĬm����|⺿u��f��B�n��2������jT:�$Q-�_w����,��ޝs8gSybh0Yd�e��1Lx���D�
����R��N^J��)�;c�j�1��t������F�Vӂj��V��^�Z���"��8�O=��#F��Cr��
O�'B
�׋�;��v-踟��0'����{�hv~���OU�y�;�u�����]Xi�v�%N��c�KUI���䮀�A����"ǿu��؝@ �۵�8n��@��m��O�gɌM/���r9�¥yal!dj/8��� ����}/)��W�J,����!��m �Kï��[mqp�D��2��RԄ���#���4�G��G޶��Vm�_��Ü�-����G�&\����&��wM���%d<UEIBf3��K/]�/[�{��0�Tms�q� �ڙ_���$�M�N����j����/�Ŷl=���@����l�m�t�5��v�͌3�@C�R������eƛg�O:���?�5h*���5��G�~��0����:Y7^<�5_�c�~��7���Nq0jG���[z�CkɝF��L2���ZD+�YR��l����j{�����i6±�P��۫n�L83h"a��� jZ�k=�G�ڄ�$#��Q#�Q&f�/t�[����t��>�U��oH�[S;�k);����x<h�7�VN�jꐷ�l}��ysiy��>!��Cb�bj�gG4/��r_��u�5��xD�}�M"��2Q����a���
v�� `Hᠰ'�z��z����b�me�A�TH8�4�I�o�r
���y~S)
�9��=u�KE�9�]��LS�d	�¯Ue���]܇��kHfqEA��}Y�Ux�1��L�eOy]�	�~ȟ��ܐ����{�O��/�|AKtmL;������-nl���������_7�����<����G��mPE9Z����*�[7� �w����hΣ�IOX�����T�C� ϋ��ʂF�d�l�-�2o�
Z:�j�`�2��KDY�E��K���"����6<d�lꄖ��;�҆�� A�b�s�U�1=�+��#��e�w h;Z�l��o�*"���DP�nz��{�!��,'��e�-��1���ȊS�	.�^0:�U��Զ�ݿ���B���o�o�+��3*��(��s\�����G^<����WÃ��*�5��L+|ި���h�5���S�ɻ����d��W�Ps-ء.s�]�<U3Ky�����m~�ϵ��IZ1Y�Y �*�u�y(r=B��0������Fm���t�~u�M�T*���L8-� Dv֔&�K<ƧKt��Y<t��<ڞV� G e���^�˸��������_WJU@��|��4�p�@�r3j��5����1�͎tY��{fP.�u5c�yCK��� |@9��zB�\�ѱ^��x5銖�]���b�t��ː�>0��Vrc9��H;t\ ,S��l��${��E�N�cR�҆�"yM~AA�1���WT�Q�gy['Mo�������� ���
����<�y$ sAM�L��2}��u����I��
���\��l�����4'Np��D<v5�3'Rŧh�4�I݆�H����<���	rtCONj���w��'�J��N�F�(�S�D�讶�3�67Ȫ���!��+�
�}��g�����j���L�*��f.~�Q���{�rh�]:�Z�8ɦ�`��܏�"+V2߼֗���}�W�T{c�\~��]S�W+ A�Ӵ��N��������<n���i^�ޡ�%	�m�b������D�L:7O�+� ཱྀ�����<�#1?�<�0e.�:"��T�z�� ��v���W6�:��.�����Q4A�vc�kK�V���~.�w�}9�r,�"$��<%*o��'��ʇa0c�!�L��:x�1�m">�w�9�s��2��<nע]*$��Q;��߿$F�5�Cx���9Hg��0GX O��w?���M�����I�kP��~�K(EѺجD��Œ�ӷs��'�ԙ2E�`�v��X9E1�I��.#����� ��}!9'F�OI�𙠎n��Z9#2&ξZM΋�q��0B�(�n�&��GxM���
�-�K�N�#����@�
r)"��_|�NAZ���3]�:�����A)l��
�����`ڪ�h�`�AÜ��w˱Q���:���1�+������JH2�Q�aں����g~٤,cq��6d~$EO��gsb����{��;>��tR���p;x�5^K���-zD��_���.��H�^'[Zy%B���u�`�!�5�{8ƒ:�I�rpٚdlj��*�I6�+�L�9dP[�_~�R��B��qƈ|�Ľ�q4ݵ#Sv��W�!�ΠO��Bm�������M�j���L$:q��C�X�Ig�����=yܨG1�hK�'x\u;�04�3;0�#�8D���x�� flP����y֝�x�Ό��F�Y�a���3��Z_�&�3�s���BI������Qf�`-7�.�qI]K������Ԇ��k�j�,��ƾa���}�x��#�M�Ѓ�޻����N��i��{�y��08!�������*�|�ݶx}Zҋ;��6��:]���R��G��$��*�T��H��3v��Lׇl�1����+wФ�������9��r�F1w5)f/u��{]�L=�CSya�$ X�R �K&aހ�xz��>~@���3� r.�0��Gp�@̺b��{t?�t(Ȣ�);�e��"+�>�c�붘���읊����@x�
t*���E����1�מ.xb=����_��5F�qY��Xk���f�A��2� ��S}�`/y����3u�(�,��b���3VI��QK��I��z�}��a�6O�Mc{;�Л��&�ԙ���A{r{bXJQ��:��_9^��G���V叁����ca���b�jj���ϖ�~��6��0��QJ2�A�(6�[%%�ck��E���y�d�MΎ:��'qX2?!]�=��^]gS֍�<g���QZO�YcU^����Pn�z�W}Y.��Fǰ��v��!����$��,X\~�p�"�pY�J��j�j�����z���|��(����+����� g2c>f�o<��q��i�Æء7�f��NY������Flf8 ՛�4�D'����1���7�����o�k�m��.T�7y
���οr,�h�$L��CI�1���y͒��3��m�N�	�hJQqH�:H���}�u�h1ğ>cu�jad��q�?3���#�V����]��\N�
���D�Kb|i������/ oxQ���(6$������pu^�R���!q��T�yV��$�+�W:���Cn�b��s���C�ܤx�lo����{��XT��>C���1 Y�� b��x6�0���3
��?s���9:��v �v_P�~7�-�p��uJd>�Z���GO������a�m_t(�`��n;E��n�����C.��C���r��Ut�ŋ<'Y�J����n��a񭅅��q����w
JhI�ӽ���D0g�3�$����6�!M���"����i�l3�ՙ�?�u�J���PU?�^`q�6�]X��ׯ�}?�`(�~�������0�c����W�S�N�ڷőD=�j6xʎ�Ѭ�>�G$őIR�6��/?��5�Դ�2n�A��]���N{��yf��Ҟ:�N�Jw�x�NE��q�9X�i� `2�NO�!�ƛM��x��O��}�F+��);l����T*y~�@F"�3�G� |��̩�%� ����٢�>�U�d&�tG0�6*&�� C������D��be�=	����4�q�H$ؽ�g��^�����$��Y�N���C���Z ��B�vr�~-ݰ�.'=D郞N ��h���A$W YvjThsg�&-���K��I�D�C�DX'��z9�������0�[?��όF-[�W��G����Jk��W$�m98�x��vr8���*[�6�9D���eU5���$�D�a�M�����B!ھ�� �!Pg��*<EF�-SKI�Cm���/�Tz�O�]�7Mk���*>����IN��r��l;��UhA͉�
�=0'8�Mr˕�񞹍�G��-A!���-QZA<j?��ne�d�{s��Y�1��-WgE˾ɄK{n׀g���K+�'�?'���C����t�E*�k�i,R�[x�U#(At�[y�C�����ݛWB�%�5h[6��C�������6p���:r3�+t�40<��G��������p��֥%�fn�9��:Yj�
l�.��{�o�Y�$�5��nй�\vy� R��`b�	oۯ�
�
X����y}s��!@�fVKU�~��<�v��܈�cZ� ��2E���I/3�/߹q���D��S��q�k{ޠZ���<!-v I�6rI^�?!ƞ�������Q��]����ON�����܇��IH�^�٨~Vc�T���n�ʋ��!WbEg]"��4Z��O�0�j�]����z�Ť�!]D��,`7h3��[o��&0��l�S�_����e��x�,T�3�j6��V�( L��,㷗ë�^7RE�/�&���(m����D�G�7W\_��sA��O��զ"U$�~`�>��D�LR�I���z&�j^vT���Sl/Krs@Ȕ_Q�u���������K^_���S���&>G�@W�R�����XY.�v�I��V��Y9���㨑"K�����V��򦶒���>���4>J:���.�]^*�M����v��Ḥ�d_�9�9 ��3�'�W���RJ�������4��j�M"�c����$��i���(Ϻ���֓�5<�K������Zy��g(�Ǳ�Q�����m�z�8�$?�����PȰ�3���&HػbXޱ5�0F���A��<� ���5{Q�Y����|�T��v��0���=�ku<��@���[�Q~��C}��~�ׇ�������Е�{ 3�]N����4�����<����Ew�r`�b;������"F�iT��*�R��������A�����{�����ٟ�~{$�J�A��H�+�=�#.z#Gj�#IMm"�!��6��T���c� 3fb�_OC������ͧ�c��~�ʉˡ�K�)5T���s@�G��{��!h�o:H
ӊ�Eq��7N��>Jkt�N ���OoPNQ��!�F?p�t��Iֺ��&���]�= �

:�0�ș����)�{�2a������-� �o�>l|*%�5�]��1p�0���.:�m����Wب��['��6{:!w�0ˉX�+3�˒I�'�M<��|�e�u��g�����y��h��Y8X<�[��ۋ�1vzv�
I͎m ޖ���D#O����C�sW�Tk���0��,���D�*4Om��25c��2J�7�F����m���i��dw�� �*z0���ͪ�<�t>9U0+a��]`8���S�T�����D'q���mT%����X��W�B��Խ[���\1�c"���1�}r��U�v+����@�iP�lqH��ۊ�a��/�	�!����R��!�j���g��$�R�T��<I?���x�m���)�s�s�;�e�7h��p��0gA"!�m�5�_���ݑ�(q�9xT���M�3��p��V���b��
�,��gR�~��8P��z�'�P������k,���{�l��*��9��mɦ[ݟ��6��T~\��-�p��V�7=��]�v�5U{~�o̊x��T�e�r�_��f��̣DZ�9�o�i��Z�3�|�3�A�u�u��nL�ly�t��s*���Snh��`W�G��)7M�7�TMyJ��&h��Ğ�{¤	+�\��νm��n���k��V�lMCMwT<g�0$,�6pEA�HB�9���B^��S�jM�7�,�(��<��l���_�G�il/���$�ߋ"p�Q]]FbRئL��#`ߜz��N��VFU��Sۙ�g�wa�Kd�r�y�ۊ�{�3v�Ҭ5��ʄC���LZ�sK�O�U�h0���-��]n �����ޭʤJ�D�300�Y����F�Fեcڱz�:�&���ÐxK��v�t���Ӷ��6��H]��E.��q."ze���1+�'��b`�ޙ�0��y�Q4����2�S�a��f��g�ɻ�Ջ�"M�G_��.�&�KA�3Z���rLn�r���U��U����tS�o��������P�fC�������|{��؀y�
�ήk�O�.o�Z`�*[U.f�ˎ�N�����'�B��*�V����p�4 N�T�#�Ż|{N���q���yӋSˣ��L�宝�"�Q2���Vv���2�����<�'	��l�S;�$��+�_�:Ѯ�9��3$k��&��;�Rw�؟vP(�5��94�4�=�:��Ft.� �&�KҾ\m��D������ PbT�f�a��6�"X�H�<v�uw���U㪔��.�a;t4��W�n�ex��Mo��b����3ˈ@~��:TN�:-�zԂbc��aW�n�	+��F
��&ي}g��Tl#SW�ؑv6���p�ta�2��z��I��g�c�@�)o�&���ް�C����J�-�?Eq�7����']��	�z7H)_�4��ұBt�_���F�<�sI>�m�cu�	���C�g2�`�yTAT<�|�e�Wi/h�Y���RN�z���וJ[��e�~!kL:��즢����L6 H0�������8p������34��������G��S�-b�Џ��J��&M����'��u���t��h��A7"�X�����Dۤ�iE���g�pV��*a��L4'�#e`�jӅ��V�`>O�Y�T�:L�E���{C���5�'�;ݥ��Kfy�vR���6��GX��/�Ro*��J�w{BU�(*��ʀ�E/p&�O�����b��X��A`��S9�ioP,�ܳj����k��>�v�ߔW��9��4���z�R\�;�	;���t�Xw>EՃ�-���+��.�a�Ք�x;����f5j��`|k��1eN��6t��`���+��?��~��YJ��nQ-����B �.�P��*�������X�r.�w���%�6L��'|��wդ㼄|8O<瓟�`#Ai������t���Þ%S��ʮ��U�6FĎ���^<�O�P&)}E���X%<�G#qClw+�0�f�t(���F�êB�X&EZ��n����n�']���T��w��^Isx�F�-�uD�֒�hw�X�^Z��@��K�:�mߌ���,]Zm�]���,|�����Z ���@���.YTB	Jyq-E�R>Jq�F	��[���b���aȴ�}�I)M>���@��0X�ت�"CC� y�1�7��@��~/7G��G���'��p��$�Վ=I_6Yz�C'�e�Ab��N�����+:鱥܁"H���	��އ͹U�|�Oq�#HF�t�߾:��[�4�'2�x�$�Ĝ2}d�'�j����g�y�+�l�̶���}Ɯ?w!A�;����9�=}l?����OT��ѓB#i�����eOSb��#RO��z�L%~��#�#���X�/.�3C.Tū6(z*{6!lWs�9�;GTuJ�U[p;���,0�V~��w������2��+y<�cm�{ I��끿�s8Wo��ܚ����� �W�"�;�V?a���j=M�k�P׷0��PϿ�6�E�]�g2Џw+8���w�ѯ+��	��>�w;�5�?g�k[F
�[��r���%�ņ��DI��# ���K8�%x-m6y��y�)#�l�G�T�jN�%��1\�`�4�~��T1��[K�.Y� �K-�
��+l���VUP{����g�Քo9,4kb �u�h��-?���l[��������$��ms�bAkʄR��k��A����8�`(7Q���5c�����7̽�qY����%����Հ{����a���i�v�>�2j�
Q86������b#��S��#��?z<>�!��Ǐ�)p�Cӝ5;��4sd��܄�����:��5����L������PJ��V��kTsF,�_��e%i�pG.PW)�3��3�Z�S�?������f��[m�-�u����1���S!���[ޒ�梯�	,�DG'd�I��&Wii2*�"F���Z.'{���_�J�O�L.��}JAQ�ey�1�;��|x��Hc�?�w�w��F	-6�ZS�w�Z>9GJq�Ĳ����3V?�Ǟu�MA_;K�~��?`��D�xc�x�E#;�!$�G� ��nD���l�1p�ϋ��)��GhvB8�L{]���0�1�x�x�P������=PdH�#`����%x�`��Z��.�L�x�Ⱦ�VªU��	�kh�����O�'�("|Iڝ��[h��E����"�A�J�S�_��|B�͝e(%����X��,��M�S��ŵ�K��DR�B@�~m���yl��l�J���2�Y���@v���hz�҇C��z0����?�㣪���쵯1��Vx�U�vl�'C�D	+ek5������G����;G��<�G1�=]Z@��ar�^/���9�v�-a�1|��8۲�o��О0w&-I��p�㹷�a ���xů�����X걁_�Q�L.�-w�O]�?̺��ک�SSP$F6�9�� ��+Z����fl;�*�ⷬ������M�"1ɯ�����	g�/����[�M��h[�W@�^0o�싖f8��mqn�7��$��[_�S��1%�����a��l$�)i,�Q�9��źZ6����.�O�qG��+����a�w��o�gl��G�~֣�� ���+yB��ܕ�g���3���C��=L�	�v����$��-�(?p�B���N�x��c�]LU�b&7-����}N��h$�H�6d7n#_�
���EmG+�X��&;�����ñ�6�ȜS��.��N�x���$I}���"8W�a��KEPF�v�7�D1s{����7�AQ��Z�ddP����E�+TP$j���/�6Nr�|4����2_#����nZ�>�T�ЃQ����_��^:�ă����=�Y�� Lh�b>-�SX+�:�k]���F��aO���/�v,�q�XL�ʚlm��I��:sOA/�o�J�b�����sCU��*��
}"�A��z�zg���x p.� ��1�K�u�#��WMk(S�.me/�Y�⮱���>��a&Q4��!J���4�G�ߓ/���jb�u���&�;�Q_#_�	M'���V���t8��a������tT�O�t����\1Iz���Ã$I�ۉ��1�T����A�'�m�2�Q�F�����ϓrioI�z����Mz��h��,�m�������A���N��]ސgR�V��y���\R����["�m*�A�:�
� ��c7̒T��뮻WB�f�a<���f��h�Ò�Rvȕ�D�GL�r��/��/��kCtQt���>��ԣ�����f�mK'�"uB<���#�~�c�9�A��Qpo+�5�'��o�G^M�f���>a��#w-ƕ/| �%�Xz�+9�����<"�_gR��k�>_�<��M/a&�B��UG����B�����]�����<��s?����vU0�C�9�PͲQ �j��9��>b`bɜ�%�
0[cܒ�q|7���$�V�·�<V�ʫi_�z�p2m�Z90�0q��3��y���ۚ�����2�kF$=��� �mf�d��	�*5����Gk`c����K8-X\y�O�TsS-?ɍ֯cGf���',��V
/�J�L@�g`�uG�Ε��jӊЭ�Db����::g-uH㮛5��}+{H��J:���B����k	��F���r�����1�D�F���α'�S��D#8jy��%8�!��P�@�L�^A �U0�ȡ9C1e��>��Ą �>;��4kr�zϏ�N�x���v;��t��t��v���/:G�)�B5���5��s���_���}�a��TDҁ���Zaxs��S�agh��1���b&������'�~L�~�&+��pש�~��_م�?׺|��dNjݐt;[��޲�����c�gU���)�Z�2�e�[��&�Yr�ų��//��w�
|�ɫJ�'�q��t'p}��
��)�OT�#���L� !�SE��dr=�Y�J�e*9>Lܧ�v�M����#�4Y5h��d�A)�G�~z�͏η5��\��3ͤ0���|�_I�H4�S}��i'��.��#�$�J��J��
�E���cu~-�Y��� F�� �A�vؚ�p��R<o��M�#T�{N1Ou�����6(;?��SDJ��/)��P�ƃ;��;�!�٘�	�)({��ggc�n�� ��e�|�}�U=�~8S�ϡ��/���8�܄����4�ϭ�V�t%C�5�k�@Yا���0���:�-�ƞ���%��S㞛M��Ǭ�rX;�_J�xG��[��U��3��yLv޾�E���x���"`ywN��,��Kl�M�}�B�3b+4��Ӧ\��~��8[E��� d,K/:Nh�yI�+�m3n�wSpD<� �-����Zs=���FP���o~��Lk��_���[��l߄�[�GM�Y�6�6߭Ѣ�l|J�㺣��-Ǡ�H
�B|�D���G��KN�8�`?���b{Rt^��L3��A�����\����&��̉8ε�~@0�3�����w��3GQ4��1���sy���UzX+'���s��`�Tʃ�>^�j�a��x��-�ɕ<@;�r�X��=_ �1[����hw/�(��#䆖�׋
�!�&ߕJ��y���,��0C�,(�5S|Ox�G�A�2�p�X�K�e����	�p�ռ&�y18�^�e7��5�2�
T�ݐžYu jBvx�(���(�%#���d(�[IŦt�o�{��7��M#���!̈�5�U�A�7�_����O$Rt�Q��DM�yc�&R�k��z��m��uk�Xʤ����  �����np��ovU �D��@�.�t6l�	�H������������a��|Ť6B�F	��~#k�[W�Z��u)L�Ht����<�T������ؤ)�u@w�����Z�D�(U���C���!��ٺ�tqre��.��v��~���P?��R�d�9,�ҥr���Q�X�H�{.=�B���y!@��}����P�������!x���y���y4sU� L�dU�j��M\?��BQF�HRb��t`K3��Dy9�p��p-�hO"ҥ��T!	�,~���'�+p��7�)R}�-�Џ�n�ه,3�c��;���ԣ(�NE�Ц�Q��k�z�,��?��-��S��^�A�`��c���D��Y���J���� �>?4�Q�����+��0���i����hJ5���Ҭ �8P������ٺ�e�c ���	w{׃����/�����~�l�Y���YϮ ��ӝ�O�%���5�C�v �H���wJ�C{�'����{���VIA�B��A��L����Ts��fq��yg�>�h�s���ߟ`��=O���}15�}
�Œ��y�m�a�5���H�
"�'�~V�`�P@q���A�CG�9�d��tH��!6�W��	���\��X��W���'�������;E�~�"!�! ϣ&�����#1"g�e��G��]�dE��3I+�8�Cf��e^p�Bo��F�
7�\�4���9W�n�������!�O�@�|�Xd����)	�G[|Ǖ��i\���:8$8�]�wRZ��_qSE �|�tx��̫@�u�f��:vg�߈��͈�~�y�9j�§V��4�|�J�G�4�`�?��ήȮm�Rx�+"���j��_��h�N��g�$��_5��u(�N�N������`�T�\J��>��?{;��=;�s-�`w���@�4���U��#M��c�H	���<���G������G��򉋔R���1{�!4����l��'QJE~�`�gw��a��x�}T|z� aV��+�j��}�{��Phn�VN�v���k���Ax$��n2�eoE���-�g�;D��i�sM�5�$;nB�h2�%I�������YlX�_�g?�<�e7i�yu�s��X�Z؂�����ک�6!U���C��G~�v	���yl��
x\��G�X��T��j ��#kc��=�5���Ye��uO��!�C%�����7d�57�,z��,I�rW�Ňħ%�����Cj>��kԐ����8�I�`�x�jK{+aN�qΪ�rP�r�Ƶ�{=��f+�ot&���?��r��c�P]R_(@�	�r��G��z�J��S��g�ڷ���Ʒ�*�I'2��`E.��.��Ɉ���~�S����
����P�Ř��qF���қ�WZȡ W,v@�M���ucl(��Լb�a�]eBĞ�X�H��~l^x���:�#+�5�VR.����XY&'5�=2
ؚ�2kǷ�-�͸��\�>��r���*�i4�E�����Z�� hṣ�9ۑ�=D��E��ݬ����1�G%l�K�����ձ��h+�ɵOH��c5��X5�����b�澤����E��O��(T/m�s��a �V�H�A4o�Z�_�F|5F��6Czzo7/�X�U)����0M#J6+s�����ȣ3'��cBӭ�>��о��%do��ݨq�!�l����dQz\�ȩ�')؈����c|Q\����n��ͼ;���k�����%�G[K�J��m?Z P�y�B�;�# W�VѠ*Ovt��G�D�7� �'�I�}̖�"1f�Z���T�o���ߑz"r{����u,q9�tY�^��@����7�L%4j��N���F-�x�Dq`ESeb�t�lP����o���Z{��D�:q=��p�HT9P	��X����;0e��e���{2���z��BPîČ��d��e��3e��(�.���0�a��fP%6���+-��n_�N��]#最'���`��(��Za1-�]�^q�Bl=̉�g���X�ZZ*Z<���&�!4��U���HR�d�˾(zFTұ"$�&��䷐�����K�_B�F��m�Ry
�"lii���
˝C��y��<a�qj���d�8��x]�)+�>lw��B�X m��p)N�� �)�ي�Qg�!d��8�P��Oj�|�'g�.T입![��
��w<�E��`�0�=n���n�Y%�u��~�p?��l�y�	�>T��W�uy��A�^~�i�ɫ9�rH������gF?p�>����g������������*v�u���L����b�
s!N�J`�ޅŬ��4r��/�����F�|YXK�T&��E�/G4���{��H���lj�bx;%�e	��Q�Q�� ,X����+D9!�٭0
k���g�e�Q�I]uE�	:����iٮ0�hT������9	�R!�v�X�T�:�|�7��nD�>�
��q�tc�
#��Eo}�\��]O���g�'�"�}�����'����sV(;�vA��L��,�����T��mֳ$ƶ�(Y�c��`==�3d&���U�$},+��i?>K�P(|�1�U� lp����5|_��~��/�À?p�:S}���']C6S\�F�tPBT�4�fS;X�Xv`��d�'��ം�Y�@��>(Rܿ$�|0�O�U4z�G�:�o��@_*�*׈���j����WJ&��@?ˮ54,%���2<�/���r��N��F$������k�zϗT�UZs�f���b9gQX�%�t���/���w{��y �|E{'��F����@�"��GSLo���51�������-'X�ً��A��Kް��!����z 璏��M:��nz��ϒNI$Z�G�<��I��@xYKM�6r��D|�UyH�ܓ�k* �>�:����]Td�idQH���}<yū�b�h���=���^$D��50�Hk�>8��E�	�`#��lط�ldڼ��b�3�#���c%t�UT\�J��a��ϊ�����]�ǒ�����fcds�h��(7����F��J��>J '��*�\�q��
8t��} �C�/d�@�-Q}b yiy���RfB6�?��H�uo��"��-?����rx�q(w�x��!�F�nP���E�g!cl9&�$�[�$��V7!Az�� n��4`����־$�9C';!h�r��5wM�G�@���)���+�����@u��#�~���bhY��_Y��0HK�5WB: �`x��<�5*����#��}�`�W�W��8+	�}��᮶c�^�o'��*�� �Kb�փ��p���/8"?'?��0���׌�(S�{qy�X�/�d�O~���%�os��XTI���ݻ�>�l`f4n���*!��:�=m�*�o�Oɍ����
g6���emmG1�#�Q耖vTP9���M����IR5>�`a��{�����q�!���[�ucn^/׌��o�w��!f������#�]'T��t&Ǹ	@�*Ϳv�߬ɫ�G�M�F��~�=�v�.U!���?�{���+W���.���{́熙� h�5�ZûU���'0�����|�n����Q�����X��`?�eX22���TZYꁽ5��?����=oT@��Z��S`hf»w�R�UW��!��X�=n��0�0-1�Y��6u�o7iY��P7�XaD ���9&2w��ɽn�-'��2���K�˒��
۫@���@,t�c	w}� ��7���(f"��/]���9�hNc26f*���f�'�w랫q#�Ueq�M�O��}27rvl����Y�
v(��zA
~
�AE"�4J�����8l�H6��`YR��'�<ǹ`i��y��u���;��$�G�:2b^�����z�ԷQ��:�H{�ܮ���ԶY�#d�G޿��� -�1��,L0v!u�BH����d.���)/x��l�
	Y���u�:Vg�����l��!�Q~�kb�m��m�0VǾ�<b�EC�0Dh���xcXG��ֶ>A#�"mY�U #	<A�w_�����]}@�>�3�S[��5��uG\��qOo\�(�&������`�uw�t_g`0���۱#�ls��5�X�2�-E*����4�M��TaN��H�v�;�FZ1�\��qYk��m�)tx�p�'���i�� �O��ά��bs�� ���)�c=�j(�BQFިB����N�J2�j��~ q���`�q<�����?J*�X��v������lY����F��$V6/���	XM/���1�?佴j �ό�0��sI����8��ǵ���"�&��TUw$s����x��]�4���<[WO�g�/i�Ro� ݑn���6ܓ��5;+w[��?������i�q#k�>C�Șr�]w1��W��N���tj4���,a��gM�쏡²Q�U�S�¢� g��ς�6�A����������H|Y���*��rs��j�����h���H�+���Ȑ�t��7QO�.(�9k��
��7d� ����*[��].b<vW�L����L6�%�t,�k6B��)^���bc���j0"�m#P"�e�I����掽=����������t  #��R�J��joBU�i�	�vJ�|ҭ�Z�G�ӜR��ܠC��Yˏ��$��ڛ�h5�ӊ�P���-LƙW(�&Z}���|�2�1�����ʥ��6�2����Vͼ�Ր��#.XW�à�Y�����
�g�UQ�OW3/*H*L[��Vݙ�!�YI{Bq�5�s&ٰ��IػC�f}�-���G0ω��ݡ�^`� B�r�p��}�� I>�� _?����n�&י���bn*EWr��+��G���0?'�3���)mɺJ9�����Dh0R�u���|����Y�k1h��d�9��k���.�)*_�0_0Q�orGj�O9�����?�*��È5�>�R@��i��9e\���g#��WBi�i���p5&��a2? �@����1F�꘬�(��18ܺ�go� �hf���T�m����K%]qg%3+��R"]"��dU=J��}�����>K�{�4�������7\�%'F+�sPgt+	�J��1%�5~g\��*�P�r�20��$_@]�p�L|�D'�8݌�M�4��]��\����U�8ޢ���AN.�7w.ǥ]�_�7��)���Q~r�4�ma��r�g#u:�<2zF�`m��xl�ш`kȻdd6�< �OVVKq�O��	�P�JM�Q��"a�����x�?�ȷ}ƽ����E�����-�N(M/$��JQ�ס�٠����s�Jn���G��5����Qe��F|;�Y�!����U�M�Sm��4{Eܟ']*pfP�ĳct[�0�w�;<��������,Wb�!�,�7�!*r^�	�W#�!-�0�1ɬv&�|�!?o�����?��>F�����[��q��}_�ʨ�=���W���_�u�K�`�*v�u��UR�˟�{�9�7�&'/!����xG����J�u��{w/M�	�mk��#�Z�i�g�]Ź�>U_�q5X�v�ũ�
%�նC~|�:8-���}z��b���r�R�}W�<�(�Pf�S�2GLP��l'�~ᶄA0�꠺ԝ��{K������~�Z��d��fm����	���R��O�.��_$�M걳�'،ƙ��(����j\��ʨ(`�i�1�w�g�������v���&?�#��c����twP����>Q&}���{�%~L3T�&�?�y7��a�d���ӑՠG���A�.uW,W߮G��),CRx�͎m[n4A�=ߡ�����uB�@� �����gg�a��aA:Rߐk>���K$��]\�C�R�����IH�%8�mq��A��	�|#�#��D�2�#�A���������Sv/��0jc��K{Ff!��J�n5��x�x�I�kwh�J(�T�I��Y�����3����@�X�ܒ�3�2������d�	1y�H��a���M�*���Xr�����n�����4�� ��K���kn=��I��K����7,����u��h��&{�ԗ`��!K9��-w �&��jI���e	����TW��'�"8�[+��e��8��"��Z�-��sbS��Q���(3�B�Wt��p5?;��2�`�%�*4�e6�a�3��)��௝��u1�72���Eg�pq�4SOT�ˌ4pOln�V�~%�#��VT2�!��[�<	��k�G4����o������>�SG��~|o��b�h�2(ÐiM��l�����ηnՍ�9����]9�Ox � S\Y�E��5wLU�
VI��>�0~^��f���α���D��<.�Q�'v���v$���^���.Jc"�f�,6T.��[/|�/�����S��W�s;q��2P��C��*�k���\%λG���;M3eb��k��x��,r|]�g�l;M�%G�|�N�+��h*��w�'f����e����)N:�� �w��0_#�aB����!<�)�e1�7�[�K��q�ۡA�)bT�L�^����7�r��(��7!����(Xe���κ��h~�x+�fO�B���Tp�7r9$Ģ!h \_-p}jF�������]���G���s�����mڲ�eXY�{���:���3,J�@��[��|��CN���1%Y� ��,���ш++X��=	�Cz�B���J�(�)��=D�.�̖���b��{��b1�=�sg�#�����炧@�o�l2�]7 [�WŽ{b;�`<��l���m��.��i�tI�����$�jk/1��B��L�ݨ��Q#�A�]���Y��`�^=a:�=3�I���swҢ�c����8w2�πL���6XkmI�����Nl4b"�WF�\nb31��d��w=����4�g�rA]������5�@u��ޣ��MEx���	�w���W؆��7�����f�r��'.Z�$8�d��f#���_�/�Md�U�p�:��H����5�7��M��b�2�w��o�b�)7� � ���VU-`t����a%c�`�_���3f�c���VŠ	�����k��Ff42%�Ƕi	%��u���^��W]��y͂�́����D �~�v���a�����ڐ�@�ɥ��I+�H&f0����q�o�"�ktIH}�d�6��g-���.��� �>���cOߓi@!�� S�0�R �s�<��t^ϓ���3����&E��0�ffw������y�Kܟ3��}D�/6$�ҳ�My�Ţ����
�2�I����=_@�Y��9D�dRܸk6f��b$�Fv#Xt�*�1P����.	�������rG�v=�M�n�>����L�����U2 .a���>y���0��A�"�
����L��>!��E��L�\�M�7V�S-��)S��`<(�R�fvl���\
yj$dH�B �".��.��pBKS2n�73��7�����!<l4�H.�:qo7wz,(1�W7��_���ͅd%�'�%XO�D6_�p8�qU�I��(`��z�֟g��-�w��u�ѹd��a�0;��J�A�����gT�� �@��C���9Y���+]�Z3f�}$���}�Yb�-��7&c�a��Ơ?���Tv�b�,���[L~��W�\:k-��=�'��9y ���GPr�̝U�
�3�۔����p �8Z��(�:�N��NU͵|��%B���S�K���ކj�����e�d['��ED�!K4��mLrE��!���8��-�D|���-~J_����@��������/��n�ʘ�w���M>�Z�"�e��j�re���9A%�X�Ǡ�3��qC�ɺ��:th��=#�����m�YJ�Jw��"�_��E>¹l6�)��֪Q�=J\˖�!�IUh����ʆ���@ܮ�I+��5������d��I���۟��~�:�P�b���d�/���%�ԓ;��YR�f�?�O��hA-M��c0���ʘ�| ���;�c�a�&�)��W)�	>�� �����O�l��\6���\�^�����à����|k��A. �[�ޔ�/���i;���T³����ӽ�vM=sһ�����^�ܚ�BeԐ�����[���G,%��Y�BJ?JuX�{��-�QE$�Roa�t�40h��j���(�zJȷ�Vѩɥ�_�W'CuĢ&�ð�S�h�����I\�\��Gd#��P�{T�_�X�9�4����UN�w�阒��A����C>,��Ov"�'?���q��3ϕ53���9��d@�M�d�ٝ\��Z3In	>��3M͡91���C�*�N�"�C��U"/�xlJ���JY�TY�0=�D�t��~2�����}���afj��x5M����Y'�	��`q�z���o/s'�#�}9�~G,F�l�*v����67�	R b��E��w0�\�I#��s=6�ɵ�������eL4JE��������s����b?r$q����2�U!Q�ϙ���D�-i��2-Tx[�K\��v��;��b�����C_ibL�j�	��j��)�Q���;����8���h̔><G`��������1�mH{��P��(tm2hn �>���y�^��57!A {y�����������`�z��(�W՘�L�4���\�o��|̄�(짜�}��u�
WBڷ<;�V�]���e7�B�{4o���QE��曹��8��z�8p��1���e*��%���~��
ՃV�� ���4�>��E��o�����0x�3�G��l��7�?� 9	�_�����I����|�*Hp���Q��:}>�m����+DO��d�J1���v�]��r�hl+"����󣷮��-��2i@�����Ql;I�k�`��*�^i�F(� ���g���`�*.����z]5�~���21��x�E��;|G�����F�VZj�[�aI�%%o?�\a��&�3�h�<�:>OCy(0����ҎNG��;[9J9m�ۮ�4�5ס�q�Xh���@D�(�n�D�e�[yObi����r���*�nm��9�5���5����u��!��r�o�I���P����$7z��F{]�if�y�Uԅ�L�jNN�q��%P��#ꨶt/�&?���3��W�%Ҽ�ʗ,;o�'^O4�;\���cק�7ge�i��),��ܚ^s=�5s�����+�	��9<�oR���P���mQ�p��=/\����O��iC�)1~��S���Nn$Rt�$̟c?ߚ9�����S�X��0E�dK�U�ʩ��y'�Q9�-r��I<�A\3i�>igN����zZ'7w}=��(ao��%��)���W�3�B���On�|F�������
ˏ�_�'�4�n�����q�'����9)�/�/�JB3%A�T5�����|����e�h��9��J'Ͳ�(F�/1�� X��!����~�w��NN׋C�v�	���p`�Kh�+�<�4��ލ�n�)h�:�Sd�4�i�f��?VMCp������Q�$X}��5]L��
��ڹ�+��;4���[_,_I��3�gA�5���1�2�|W�?�ڝuk�ZTy�ు*�*^	Ic�P�9<T2l��U�!*��~���"'I7C*'��#鶽� k絯��ǫ2Vqu�ʫ�N�(ծ���Z�}���E��0������W����u?��h�M���#�_N�Po�AMw��ȧYU$�E�#ك��Չ���� [�
�!��^É�Ϳ�|�q�d��|:.�J�P�Qo���Ę1�C�N:2rmW�[��,�c���[�Y����rg���Jf,~a!;��z���(̔�e{�i;(���-��P� �ĸ��I߻5�d�5V��t�!��~�=b�2�U��X�]~�᜗�s�O�dQ��=9�x��)#Q�Č�@i�n*߹�x���w{u����]X�Rf=�9 '}G�͍^��vК�M���$�b"���j�l!�"c>��7��
[�%C���J�S&��YFd� �.��ݙR�%g�8	(�<�V�A�if��T���J$hK�u+����j����Q�#i,�q�9��p��nZa��q�;i%E��Tl= ,�L���;Esi�Ԋ�}hG�ά�u�X$��Xk�fd�\ E;e����rlJ-�-���;���Q�}EU!l�@O.j���"2r6�R�7u�>���θ�� ㈨���ֶ�Mk]�_/%qL��Gq� E��A2�������ENtYu}���=TA���=�}uR�ɟ˚!��3+�j
�xi76�zE�D|J�j9Յ��鳐��>/�����-��tUƉ�q�K��S����o�Q��X=��pxnbc"��d��cI��"u���21�ב��BgC2��Ca%����7�S�����g���v�J'�&J�80	Di�Bi��m�
lY�_r�tW�d��*W|��A ��B�W�V�x�$�o�H��ޯ�Q����O�Yb��R 1�m&��w[�K�6g����D,�Ë�I�)@Bk������5���q����� �m%���m[�TQM*��'T$c�<9U`�`����\��KP<�$A�LWW��l^g稍����m��,��6U��.������E:��������U��Y��2�k�߷� #�g��qk���p��:�W[�'E��ߗY ��Є^�CDX��Q��7���W��i�R!g�ڒ�&�1B�Pwbo�B��wq}�����Z�6Ī{j/X1�IB �~�і�o*�����:t�"\w6ڷ����/QmR���k��>O�<�xe�UE>�`/���@z�������+��~�I���l2s@ Q�)G=��ײڿmR���c>�n�hW���8B�G�I�|����x�/���N��Q��8Z�ƛۭ��Meg���y�8�Q�71u���ԮK�Y$͉	=R�8�/D)�1'�G�8�B�	�Kյ���:׿�pG`�8n�2\ٲS�T��gR`۩�����O�E%]�}H�}�Lw��� m��I�����`�9�{�o���c�0E=��!�D�������j o�n��/� ��I��[��؄��)H�P( ������z	q�����}�Vt[o:�eԬ�
�����$��Ϥ��������gǚF�}N���^5vE4�s�!�P��i#����M r$��T�g�|�4�6��tM����	,�+��8�/.'�jŇ�҄[y:��ce�)��I��;]Ax���I�x��E�B@��=����͋��O�O��9����;���Y_�(0T�)2�x��:"�.?"/���3��2Wǚ��1�����1�}��I��2L� �� S�Z��j'�����p�<zY�s�����W�`�Ʈ�~�������ЛNpH_������+.��W��C���"*+Ɔl�<�٘Cfʵ�#�q]EW��@-P���f�����q����L��5968���c�N���� i$�у��w<O[n�E�~���PzY���n*I̽`�,s��}n��� x�'�^G�e-�eA:�`�3��s�YG�=�ݳZ�݆Ȝ+	ş��{�~�_����v=d�٥��Onm{��G`였�z��+mF�:�I�?�������;��'��`�����#wS�[���rպ�z�� CK�S3DX�k* ��b��S�7�a�Ҵ�υ��vt����8"a\�����|o���L���g��r:��2ٲZ�{.s���&��!`*_�X�:9��>y�W�U%��H1ʗ7���%}UP���l�>s�p߸�p�_�7#��W�V�^���YSߤ�pB��_�}��9��͕�!H+��8��z����Sb!>������,9σ���Ӄ�E�v���{���B��#=��ɨ��#��!����J>�]��RDq�cZ,X3�h0��̛�ǲN��P�h�Cv㨞�Umۿ��vy�q��A&�LrȄ	F�r�/�fЙ4�k�NZ+�I���04({қzlp�+�k.a�F������At`'_�]R���'d3!��I!g�P��d�wCx���[���v��Yy(�gQŸ��ޚo���2#��-;��9�R)�E]��C�����1���P7*	(�8Ck����E'F����	蹅Q� �.b��3z[bu��l'W�Cz��Q��j�̯�f1����2������х���O�{y
QIo���7�����]EÁq�S�&`��׋�^�ܬ'fp��F�u"�����a��S����iZ\j	�X�uP�i)L�%]!~��kB���+�	M�/}��.�pFh�9����'�U	��Eeѱ�yچ����4؅�Jm�΍��S�����2���[,R�	��X�*Ƨ��U��F�����|�V��N�Z}�y�����A���O��*����R���dz���mј�_����֢��Q�-j��<����kL�Fiǆ�Y��ܹ;�x�ay�Z�׳~o{����
[��Uーj:����M�j�ۡ�zrEMQ]��F�������Bٰ�
�Gp�%�E�m#�6/�M/~��A3:k��Ws�����H+�H���y`^B%(��ب��6��������z���Q9!�t��Ȟz)_oB��-��
�B�{����>5\�~WN*Al�UTr@��m�-n_/G��$�%���/:����E���:Xԗ%h�֗ZE}�˫��`�i�wJ�W��t���`��A`��/G��tKWY�E�q�> ^?^�9�dcNpE����9�B+^�,�}�j*a�i)T9[�0\64q%��v8k��娾��6���4'=��9�2�� ^; ̟�o���1$-Y��{b�)��y�Zy���U�,�t���ޡI����1<	Bo(����f��9^������v1�9�JO
��ʂY����=Go�����{ά$�)̝���I��#z�~�ˠ.\�C��d_=������)w��a J[(�`4��� �q��٠a4<�B��F7�8\��`����=����\��@��ƅ|x��\�_4���cJ�$|�3�CN����a���F�SE�=��;@j �mJ�o�,���hpcȎD�*��e��\���k}�гf+���+V�S���`ć�$3O+�F�1("�/w�����W|B�-����l��4\R�T��u�۾���c��@�>��#y'V���?���6h}�(!�Ofu�7���F힗r�"�C�թ7����ȋ�%�heΨ����]TcO�g�Ln�����o�7<1d��BkQ�_a����,S~�O<�@:,��<�6"�9>�2���v���}�\NX(��3,�D�2c�%[�8F�mo�WO��d*�9oe�@Y{��8�vdp�����D>^IN�W�XGpeؿ�s�WT�v�{b�d���9@�H��Lk�͋��wנ�&�����"j�,���$� 6�M_p�ց �J/4?��g;�e>䬝�c+�.��m����]t��Ypt�D��B*�����I�"v>�j�7��a�uiݎ�s��db��_Q����z���	3eMgӌ�x�S���ׇ�).�>���z��|�ہm
�*ʊ�dg���iaW_���V�~&���q��
�6���r��Jȗ�C&��&.�(״����)@��2PwGm�RY�����7�|��$	v>d4��������a*�pAa&�'ϐ6�csQC�+��X��φ�̼�Q����6��<�O���f��k"�o3���"�>�5ob��Qo�|�&C`k���n�~�g�G��\��1n�����%�˶�;1
�+�^_�
F0�gZ�B��
���ː���jr�NP^1��R\q�Dn
�E������bh@K]Ө�{<b����@�
���a�(Q��(�KQut���:k2�렪��Z���ϣ�h镬Ȱ�7j���&-�h_X	�6l�3�~������G�F*/���4��Mb����cT_���G\�Z��(��h��W�C�,���w�n��;|��4�~s���2&{^�,1��p����ϖ��e@ݎVx� ���qM�����C���������Xt����ԄS�vƻɣ�)�H+J�$S�k��t:o:�z�g�Y@Y�T�#�6t�G_�j(=�Q�>P���!�(���g���ӨtՐ_���h��_E���q���Û��<G"b�����.�g���hԦ�F"��� _8�wj��RrK�v���=�Aw.���u�U�2v7i-4L8�u`�x�d�~,�/���D�,��1tu
��@�$bV�R��F��H5�N-�`���ɒ+ (���I���8y�0'�zK�]��E[ۉ�L���Q�$����,��Ǝ��0�F]0����S$�i?��d\���i��Ę`xK�9�iZR��կ7;@�Ǣ�&'x�J�]��P/"�["�r��ja�X�B���{�=:εY�pl�=�+� �8ћ�P�)��%
ò�ck.)@�4n�͸�"��;��Vf"��� >J��FT�iAG,��w�q;���h>�G�~i��*D�N�r퓓��v��o-$�k�ƞ#��_"�S�C��q���dRۜ-p���m���Gb��H�"���8����������_-Q0��o?&VH�^`�>[�@�&F=���c��US��А�[u�]�/�iL�e�^���M"b�Ofn���0hdT��� ��6?˟������`��'�='�i򴸔�<����\�Y�]�g�b۩g��?���YּoQ��D�6�`�mSR����P�1�s8�cdjEHh<�"t�PC4	:f��M�&2A5͖���Zإ������~�G����#	��x�'OAg�ձTyV8��\�ŗ�AK���8+´��,��R:gwٙz��+�_� �x�\���痟qގ�C���ܗi0O�]����M�ҟ6��L�K��1F�y��a�H��Z�Ng�.�c:J�l~r�������O'��yl���v���Ku���V�č��mڗ�`F)�>�t���"�f}>�d��ۺ`�n(��;쉛�Z���(@ܾ+ژ���� �ɉ*�ū*�-Z@][�*�*��с�a@��m(�ѿ�!�?h�@�1�(��ē�!��$4z>p�b;d�
:/_��MLЯQ��V�r�G�-���]���ȋ&&4���R˔;C��U�7�E�槵����~�9�V\�"��:����4+�`���ͩ����Ł��!J�R��	��2������Q.*e�Vӫ�G���V�9�
����ܴ�fH���=��W���-!����R#�u��
�4Q� � ҂�u��u}� vL��y�˱�1��h-���$_B�����o]H`P�Գd ����Y�;���k��Uµ�p���| ���ױ��#<hd��L��Lf8�Y��]Ȓ�F?�EX���7ˁ�+K�bE��XT���%=^"�hF*ǭ��u�=J'<zQ�w���+$P�W�ɰ}�xx��;q�.�JOF��3�|�F�����g||��_iBn��Gnl�
*x�~�
~C����^}i8�z,�Q^�-�35�[�Qy��΍^d�g��Y�G4��J¥��T�k!�+���W^���ꃀF��d�N��{S���I�ͧ����U�vb�}������c����[)QG�7)�iDc��!�|'���D�b�W�}�إ[�Mq�g�{���������=�=��,Y����^K��l	o�q�Zp�5�y7����s�T�슥�ܯ5X
����y�b�F���ԅ,���L�1��"��,�Ie���
�����/�
��I=�}�Jq����[��*s�1��^�����+_�,p�d�\��]�]ko������|x�I��J!��#^%�ǝ⺝l�P�'1��x1�w��	Y��k=@���gz7&�\(�U]s��`	��p�<X�V�&(���ZL�d<Y�;l%�?��)*���=�8��� �CfMU!�?uYOҗ���F��Δ]�_7h��2� ��	��.�єg����dA�D?=ak�ܡ��2c�i��Z�K��9�e� 3��/wf:2���{{X@d�o!X�W�aMaF�qby�[h��f/�u�8i��`��E��P�/�rT�Sp�VX�?��\��f	5t]E[�%�Zǣ�Mv�����ǽDa4Λ���	[��g�Ť/�%�N8<�U�8�U0����%��Y ]/�81`�p�E➌{@�.J�~�n:"]�ܽ�JC b=�X���o��g��y�����o]���nc;��&Z��܁�K����*���*��z�!�(	ނ�{a����w�w2.#����8bTM����6�$܎��)[����ip���pO\ފ�2i��`"W�Hi��F������%���x��%)����揩��g��ʸ`~�|�Ƌ��k&e� �5���
$%B޿$H<Wx���K�T�%�p�HuP�Ÿ+Z������
�ML�a���+�'��?���ϛ �R�9#;��Q5����H��2��rĴ��#�H�Z�8���V�p/(��7��u�k���L�\`1�?���<rn�I�k�8��G����BBO{�o�-�W#��k>H0�:\�N�.�B!���!"����#��l�:/�A ��/�ĉ����֗��/T����^=|�x;����C��i�Ø'd^O�?��-"�e�U:a�@���c��U؛�r�T*�wl��׏,	�^XQ+%C+*��PNA�yG�4ʃ��$��i��#�^Zd�;���"�����nS��9���C��A��L����f$n�\	��1ȵ%tt=z����M4Ek(v�9Щ�u�}�Ĭ��׋�G{)��a�������CĖ���=�����>j�䎯?%�����;CQ����~��~�`���YAE�t��;�#�i~ �q=Cm�; ��4߷\3騇QxK��) �~�[O9f�����Kޚ��Hp�mre��2�^}ʠ2ĉxJa�EX�h�J;/��B#m	��(%YWЇ��|���m8b]�P+X��	�����:�� ��T�օ� �A&��M���$����^�C�����X
��vvu��<	w�q�8�4�BL_�Q|��R�ɠ�GI��/�f�^x�P�����T�)��!�X瀺�'��O{�ֵ�8���L�y�gxh^��#pty��
���'���)���X��`���!�k&Y�$��S��_���#0+g�1ݙs���?I��	e�(c珻�hd}�Ϊ�׺�����/(@^x+������̨lh[�����l�D�����^0ӗp�l�w�ο��i�c�}[��iz����W�y4�Z�I����p�YM"��	%2�]Ťlr!���[�ّ�ANC��T�)G�.9�z�@�DK����m�@�5���k��vu�/��-�n4�C����|P�iZW�/����hx!�	����A8Zr����>_
���V���a�F7 mXm�WB'�s],�Nt�&B�Rz	7F�������0��E/�쥼M,"�O��kOrg8u@��}U��7�(��Ì��_IG��(k��f�w��(Bu�]V��<�g+��	���e03����#x�<����W�h
T�O�E! ����*?E��4��%�~�&~������XC�f*Y��ٹFc�Α=0��%���vw�s �'=L��X)ڨ\�����
=iw48h��o6�L�D�Q�ۦ�(�IJ�V�e!�d�a�UJ��d�kS�Ic_U���O���M̛E�=	�}����S��-r5{��)�*���G�>۟�|����#��%w<q��`˛t�ѻ�rU;u.���qwj��@`[�E��ɺ��
�m�#�L�*3�Qi�\+>��C�8�	m�i�=O���Bܰd��2&e�D��5����K�j�{�P�V�Tp��A�8�v�D8��J�*Z�ҍ���z�R(_����/�&\���,�]p��~	��\d��Z�-"e,n���MK8��'j��"HH��^�.�@���x�?���Q�+�WN{�g�\��]
�j���L�=-?�k)nW~��l,�za�m��ꫠ��J�}N�t�&�:������DR�Y�
�	^��c�o��?��[�{�e���� ;t0�ʈ�8������2/`��_�o8cL 7 �n@��섶��q�y&�=R��ù��Ty��˘�xj�װV?�O�t}7�Fw�P�w�����T�)^O�_�r�@�ӕ�M{��:�j)z�1Jz���Z�aʅ��AF��6nV�}���,g��|�S<FW�4�
߅�;����r1G���m���H�+�:bs/�% t����an�K�oW�?�Du�w�\��P~��&������ĝܲ��!9.0���I��� T[��f���F�4�e��C#�i�ry{� b�B�2Q�r��m�l�T�M/���k�oQ��c���b#X��v2�v �i�$�Sy�=����t������ص��#��?�~=4�^�A"+���4��R5���S�s��nQ.	��Xǉ��U7�?]�t�Re�ӄ�9�E�Ols��B�|��T����@=����o�CSl�j���`��g=4n��7�Y�0�b�r�$�/nIq��߿�9о����.o�R\�&o��j�9���p�F�v@���4��N�we_���������$�c�&����&5���[�j'o;��h "��7�u�}n�(����Q�֫d^h���?��@��?Ƽ�Ɯ�f۠�]�/��E���1������kH� �6JԸ��l�2Ȣ~�0�if����W��x���vjf�H`�K~Ji8�p��TO�m -�����ݳ뒧�Z�I9�s��f�����=�j)�c�װT�r�=�n!%�pg���.�����>S���<숴�p.�_��-N��������X�y�F|O"n���l.iF�����?��K�B2�e��PZ3\���"���:}ڙp$��f1����F7���9���_S:�c&j�(;X&�%�yI��ДF�[�aʑ��d���%�zI���g^@���k+�`�6���
S��&�P[�헯(� �i�Ƶ�7�ç���/���YĬ+b�����Ly_�L�,�*������SEO��H�JJ����>앲�w���.�/�	T��0��-�d��� � �*uD�d��ܐl/�{{Õm��E��t�Mi���Y��S��X�0*D;(���5o��W���<�[�<LR��4�����N�e�I�)�C�@�����d�ȼ1�CƷ��ҧ]]�k0}��1�.�9��A�@ɵP�<�֙P@Ρ��2���R�3�tE�7r�8��j0���.���������zT-#7�} ��	J,t�Cս�u�z4�ٙ)�IOa��3�.s䕌xM~V ����r�;l���ڽr�)��1��\�#Lm}����}O�����bO��-��'�[�-���R	@����X<3��`�;-u�2��A@�Z3��Ƽ�?�|܀��#����n��GCЗ������~��t`u�����[���������M�e$�6L�3�C3Tm�dO��NB�6����g5���<}�E�|	�IZKx�XM�&#	���$4�lq��y�!�N^�W2IS`������;��T$��98�O�����B��/��Q#���ҎXƬ&H�6;O���v�}t����TB!K|�J!�\w�Q:��Ԃ"�`�k�����b9��3��'9;�/��N�4DOƵe+>(֨k�򠟭���m9?���qB�%*�cr]�|�H��!:<�I�f��!������t�~Ю\ߑƲ����
��Ԇ�����;�m�-�6L�`��|�f�'��h����a�jp��>��M�#���>�j0�JyD_r��#�������?�y%os���ߓJwB'�x�}�fEo�y,b%(h�8����$S,Lh�G�6�U���X���+_��+$}	���Ϋ�8��l����U����nل�`�KX5�^��C�U�ϗQ{���L��t��*�w�]��UC��?i����I
/;�.)ƫ	�W�~�D�ؕ>ܿ<�W�4(`ȋy�{e�n*%!VZ���������|#g�1p�yw��72dI��Ro���(L5bE=��֖�Ż�@�~�i��{�92.���0�+�֥�-�s��Њ�U��m���=������P��G2��B񥻼~���ŝ�>Kܨ��������XJ�t��P�Ԍ�Z�@��ب��^�_Oi����״�,m%�������1�h=�m���m����đ*U�._V��_c"~��I͌.�O�X�j�EKXgg��w��8Ҏ�M�w��5�>M'o���L��Ek]��L���#��l��j���ӆ}��@=,��T���:ɤ~��9+�(К�S�:W��zHuV9YxԇCKS�����_���|���2*�� �o�b�?�	G	x�3���
Č��-D�L��ϻ�yU
4h��	��Wi*���T1��N�۟,= =:6��l(��K��N��gupf,��?
��Y��A{��LB���Ϩ.I�R�a���f{�SI!�B��Q����|�gH;a�����?
��n?R���ڦ`�E�n�Л�<`��-���r�Q�������iB��|�(^z�p[�(霗��D��3�S��$s��^iO���'ua�?�����<+x(t��m��IL'���q;�8�hd��?�%[�|�����A�̷��f�0D����0�j�?��,:�Yx�b��",���}����xڼ��Ys��=�tBJь�L�2s��,�N��4(���1�w�����{��8�ؤ���?F��O[�F�gw����3>�61n����z\,�� ��6V��p�n�/b�VR,�G1U%����6���Ǚ���'���?%����1->雙/��O�Nԏ�(wJ�<]#�Lz��Wܧ|���t)a�Z�Xǈ$��ک���'�O���3�]9��
-P������?c�P��6c �w���!l��f�m�`���\V�m�5N϶�s��`��g����*&^�@���A��ܯ53�
r=�E%�գٌȋ��:4�V��L^�9K�yz���@�iq�"a���]����-���=+�~�!�)+.�(p~�+��k%#ƛ�W�n�)U�`o�8���\�gĴD�9�k��Y��Pd��+�u"rЍ�����Y��k$
�F�4�qp�I��azHd��
����-�6����*�)���$����+�C���i7�My$C�&����Q�����M��]	�R��=-����KR7����_Ǹ��u7�
�& �)5�e��wvA_G'L��0Cgs�aĸ�$���å=��D�̦��G�z�3W��YD�/�N4aƥ*He4!��$c!����_�m��/>%���BJ��!O)�
�D1>��_ଳQ�[C��&z?'Ǜ�2���a!z�=a��8���O�$����]G��İx!n\�]�o�����t-a�2��򽝏2A�%�!�iO�/�U�LF�Tu���M�
�W)�5
S޼� �rcʒ-��t����@���u'�-��C�#�y[��咅Ԃ��_KC'��x��;y��f-�t@��5Zf�xb�Y��^�ZQ�q�PXHr�&�Bȫ�i؋�vf�O3\�A�����t �ЏZQ�<=�A&9'&�^l�f����K����S�]�i�nw+���1-�v�K���a�ќ����0��w�	���"a��o��~�n�|�2����~��a�
i��T�*6���9�\e����Z[��Cl�ԮQ����������%��y�؏G5H�_?�UPǋ�[N�
���j�-Uu| ����c���s��̿�[��<�u���Ú�kt<�c�-4*��Q�`JW�?C�#��ff�ǅ?���7$����H������i��%���uW�k܅�$.�Du���|b���ɥH����T���9m��<x����_;/Yӄ��E��1�Q�$[yq{��PP����9~���W�Yrj%�(�KF.W�G(�g/�d�����[gkwq���NV����Ko\����	����N����Զ�?���ûc<��m"yU��<D�����U�"s'_ǣx��X�ɱG�7l@;� �"Y��ճ�6An�Zi�#���byU0˓Ps3�����,6_�!�ī�0'"Pg�(�����u�Y�/1�6���S�Xޘ� ��Ml���DG����o4��3B�n�'"ofl�
�|��S�]}��L�det��d��Y�g]��4�e?��N��Gïd٧2���!to��$gM�m"j.�>�;�\:����b�b���>���.�Y�)"�$m�7#Y
[]��SD�G���O��Z<Tڷ�[s��!��Fw�8��0]}2/|��9���@�C4�@!�5e�ҝp"F]K��RƳ���� �$u�ĩ�apjbn�����$,*����V�^�=T�!cm{*f��~�=R2�pKf[�n����V��G�˔PR�ǒQ��U�H�cځ�"|��)�o�S��'r�B��m���O�&0Vxc�U�R�I/���Γ>��0T��:���ј�v�-\r��KL��9i ��l ���yk��+Z�IH����*�W!�v���D��M��k�"���Rw��A>�,"��(�^�ؤ�n�Z�8C�n�a��L��D���bKۢ�=*%��:G�b�O���RЇ��x�/q�2��
+Vy�	X9��yB���+p���Y�α�X�5���\�A�
���6zR�J�:�� }Pw#��S7U5�YgyEV�SGN����5z.�At3��)�RJ2DI����<�U�P�w����F���X)l��D�!��\>|%b/_ �)������P[����t@1�Е������-dJ�V�g_l�]|���I���c�C7�^����pP~���D�&�f	������AZ� �S�p�R��<_O��$(J��X��0|C�[���r��2��^`�+1���W،� �X�~��l�3���l�`R�KI���B:R�ԝ�\�QLv�|&)k�맮W6���/���oh� !N����vŚ�-@A��[GĹ�3�R��cYBc���<җ�ޤ�����]|�U��~����؄gu+݂RTs谋źy�r��_m6�Ah��yO���zu��|�ˎw>��~�f���.>S'��?�<{tKU���������4j�F�_��_)F�rg��.���l/;�"�Xk(�W��@7#����Ŋ!� �n� Ю������B�2~��.�$Iq ��ڔ}V�<[Jo>x)Dql���� �k�������{�LI�M��=�ǻ)Ќ��$���`W���)A���DQ�Qb�aB����xY����y4�m��*W�y�H���܆G/W�njl�a~Z���>_���NZ��b�x�0���H/�&|��w�ꦺ ��)��^�g��_G��T��}1.��6W�:�Wv2���yF�䬩���ʆ�1����r6�t�۵Ȇ-�a�H����E�}�%*E?<M�U�	�(��G�����y�֒ٽZ��w5��u��i�V	-;4F��z�B+�<��EEd���c���VssY����)�%���z�F~�!�ӄ����ퟃ�=A	��5g���Q���,�z����H~s��1���v_L��g�t���@��܇��`(��Ii{�C�I����]*��Ti3~��������"���(<Ùq��Y���<]h�I�e���~��Q��+�VN������/&߲�uF��imX(<�
�b�~}`&tQv<��7���`����d�pwQuɑ.:��`#Z��uXE ��O�y0�"��-}���M�)����ĉE�#cVa�13��*p)��e��ٌ����G�O�*1����.�n �ٟ��t��}�RL�s'�]��):�������}�#�6����,������'U�屭E�I�p�(�Kϻ��^k<��/>!�
ވY��l��-����>A�h�4�ȞF���.4m̒�3��;�,�$vnZ� 	��!�Ǫ�5�ץ�6��f���	��-'�}�
��tV���˼�>`�a�}
�,�򆦨�C8h@��(��{� ?V��2��]/��TЩ.T��eD�x� 9p��H[C6>���b��c�c���J(
L�˝���"t �B6�~2��S�4tK��@��S'u f�z�q���SqPA�N$	!�HQ&��\�/��u��#]��FӶ�tp{����`��e���0����̵���u}a=g�x����1"Rj:>bS���l�D�UhV���z��'if�Y�cP���/�.{�m����+�9&w�=%�zE:+7���y�}4�@e��������]��n��Uk���*�^'V �ALE�����=����:�>sZ��כU�(L��,F�(U�I����o����A8���'k&���dI��.��Wӭ�����.&���z�Z7��g(�ʜ@�B�P��VT�043� �4贮��11�HI�gC��&8��z��[��*��'�.���m�N;8�
�o���Z��t"Y���ȑ>��l/�	��"^�H�{w��`4>(�[��i_\�L���m>ou'ZrM7�.�a���2P:׋�U�.�(���\���)�ҮTZ,sB�E2��?��'�O�ʮ9�c]>��630������%��_��ϰ�>RvG'$6VE�Hr*#>t���}P5�V-��׎:F��ܸ˦˿��MGajF���z���ƀhBm�|.�ߒ�|��Z����5g�}/��|��%iT|I�m�^н '�$�Gb��?���$q��\g&�׬m�̲H-�U��=�n�R�`���O���W|�@�<`J8~���!*�w�z!�-��"?|M�]��Ǳ_��@����%�5���l�H��k��օ6�S��(�ϔ;Vf-bF�'�&�#6�Zc5�t�C��!\vm"Q�/�~�S$�#�y��������#��Y�K�9�y�ՠ$�/�͚3��"�ʞ�1<�M���(K�<���^�,ƥ��Ո�p�E�6,9D��(�;&�9�W=0LGXOԲ�V�"2Ѿ:�g�1�n�\�hg^T1��KT��İM���nV#o��&�	ww�[�r�--'aX]Z
*��C߇5� EU���Wq�w]��+���������'-��h��#�Za�ϲ�r�g��(��%��D*�؄��8��/'��af*��n��zK�3��M�I|r��2�S��߷E��"`�*�ɥ]��-�Ui5�������M��\Y o��^�kh,����y��M����Ce$�GvN\���M�&����6��?U�}���P��ROBK��&��.b��Ƨcա�g%@9�J�W��	itq)k��{逃	!1�W�z�{%�.inAR��K��$���u��p�f�y�Y�S���a��p�T�8's��o�2-�I�`1�8o9�$HQ�⦅�|^kF�����C�i)���8?���gj�t�Xj��ch8�^v�J4*���V��6������x���`�1'�J��i�F�V�y��悯�A7��)��>��\g&P���X�u��O�bY�zjF�U�Qq�#�x�"����ս/��%9���7`��񫶄�X8�k��^���<~�=v�Z=%�	ɢp^�v��M.����㹢�1��w�n�J����2���C]QfT��uw0�Ds�\��N��j��̝W�y��s�������_�U�R/���^hq�����=D	B%��,��1��᷄K%���p���ɗ��Q.���O��W��|����`�F�,���:�Á5&��_N[���H�X�
�/ס��B�������Hj��IG�_�@y�8��fpNqel����̫r~������0�2ʊة|c�^�7O�:	)k����ǉ�٩�j�L���f��	��43�R��\�R�%6_c෱�byFfmҨS�fX:���ۜ}�%��R�%��>un�4����zk�0VQ�xM��(��d�D��I	�$�a���~��������\L=Q�P-qA؞m�R9����19�k���t	���^�p&��Ŭ4eQO/K�r�3��~f_2|>^Q9��, sw�p��7�Cx9	�s�A?g���O�5ƥVa[�5��xԙ�U��1��+�=�#���.LLg����GJ�ʚ�����9�N	?�K5�	�~da]�K/9Ux)`<��~�ƙ�A�J^1�a�n�m;�}�$g�W(�||d���;�a~��	=�녉M���~G��h����H�^��/@%�c���6dk-�F�ֿRc1�ow���3s�X����쿙@�ü욫T>���������6�7�����*9 �*4S����J�? �ڿ�`x51�e�� �+�p�  ��Z����.��O�����n�S�Ԙ����H���$=~b�hMBZ���ú�U=^�#�F���;"��"Ky����}��h�=)TP���A���+�L�:���G�-%*6~d���t����\�l�Z��l_�PMU�3$�XD�~Bj\���P#�J��^tN�{/�W�{� 2YڵX����3ۧ_/�ju�-�����{�k-�?oV�&��
l1��mdj C��`����eD��FdQWY�(z�����J��g�|�JP��Z+�2@N;�〻�Y�7��p�6p�/�|�Y.��޶��Z�s�{D���M�g��}�DFqS���t'���z��蓽�/0�,=����/G���xG�i$p3L���2m%1#��N�g0>2ˇe��8)j68����9�3_`��1%9XD�4 ���`��ҁ;��$Ť;�����UR��`B�ϼ�c+��D�~��zj6'ۧ�#�|�5�q�ǯ������թ���9�� 7z<K��y20=o�f���wN�,RD�<�'��.�s�:}����Y�F<�m�f]X�b�����O�����b���a�<O��RǙ;��4���mQ�0g�یQ>�Og�*�E�\E���B�`���0c�f�owO�e*�����kV�����Ӷ8=��ՃS���1�N褅�3�rʹ�l2B3D�}W�s�Ė�r���ݝj# �s"
<V-�;�Ɨ���p�[����mĸ�K�����SAz��j�$vg����P�i�#`���W���	��(���H�#�#��o`��p0�$63������63���S�l�y�ӓ�Jۉ:?�eٌ��m�]��f)!��7l�fsu����<��BC\�c��ө״��9�^��n6�a���Yc��n*q�W�7C�	k9�Ύ$���cZ�,�WO�*%��>= �����H�4�����EH�(b�v�@��U���L�J_&x��]l��)�k9��OރH�u��=���a~[��9R]����=��$�l��Qev_�!`�I)@�m�� $.������PQ7�"�UދX }s�Ȅ��UC!J.#�%w�����T� �t�F��x�ܭ|���W����_�M�zif�4������})���6!����թ<8$��6� 0V��rƂ����"����P�d�J�h\3��[&�!��[�
�/P�(0|�|�<��9��;�ό�����ƼϼKI�F�޶�0A�]θ�K�kQ.�Ke:J���+w�NU�X��h�^��K�6�YH�"�}͋��?i�&�#�|�}v`���Y�p��:�.� �yVa�X�_�BYp�M�-����B��h�7T�X$�,8G�u��\:!�E[泌��)��+�F��2"��U­Q� �"�\����`s����	o���FbV����S�� 8+A9ohd�C,��!��7b=f\�f�jFH��o��#4��j%\�Uh�a8SE��s�X�������voBMRS���b*v���Eg �ߐg�~�_¬wlB�}�Ha�����Ow��߆"�cЃ�T�6�tA�����qM� �P��3H��9��-6�O���y��py�MY�@7�9��=����,����P7�tM��K>:����/��K䖋V���?��<g�-�1���ΕX������㿰	APq[��u}�L��a���H��H�	����*�;|&��$d�٧ԫ$j���!��g����b�D�M�&�6,��ڟq�?>�B����%'��ivHz<z��I���wPR���Y,J�q�����L��[���)M���w6��\����XB�q���8�����
Mmա��U��qQGK
�]��M���Ʌ���P�A5��=�@���ߵ������E��_�N�x%�yՠb�q�2!�VX;��V��/�%9i;ls]��t&�5��b��7nz��WqIH��� ��0CaN���775��RZ�z-�Z�;8��5���twb��9�m����&&�x��KlԊ�����-Q�hK�x�"F᷃ݵ���(�h�j�y=�-.�gɐ�p�a�Mq�a�=ݒbu��m �װ�K?�?#U��\f�L���������!�w����~����<���:�3Y4Oԑ�?�(�������Q��?�]T2*�?\d��f�68�����@����e�2��/O.����t�u��|¶����#B�U�%7-A�"������=)C4�L|��_����e�%�w�_�=ȭ7K�,�^u|ªJ��#�E�is����C��.%m%�^�z̟�ćbo�T2cPCTN�"�����
���)��HL�U�N��m.���1��5�ʎ��B�:��1}�$>Mo�\��>���P=�~�K��Z>j ����=,� f���ڈî��j�� eC1�4� �����34C��K���i���~Ǟ4(��r��;u ,Ց3��a�c�B����Q}�m�{ʭ���yy4%��#w '�:9�cp����wJR���u�3�Y�1e��bb���p; �^��N����o�c�"JW߯H��r�A�`D�O"���ӳ���.C�+K��<c���6n���Ǽ�Жj��%#C`+LmbF��l��H�˚LUԞu�_��}�S�[��3Qz&h5�3M2=�):�.X�����e~ɀUo ��)]#ޮ��)9w�6� C���\�v���:m����:q�!V�6Ȟ ���	�@,�Ŝ��Yx�nb�mPf��'��/�V��D���=����_i�o�d�7GO÷�4�m�.P�u�Ph��,�/� �VE��	�iߠ����,�)��R�l�CNWz�y�;K3q�CĜ���Ҹ������uc�����f���oÞǸlD�w�9G�Ly"Rf�>�^�=�:t�!���0B!7��}�LP�w~�2�v%�kn��Л�sY�Z`�v�6�@�^�\Ҥ���y7Dj�~}Ư6yu�ˇeg���_�?IʜH���"�6�a��&o��}=c�*��	�,��s����+���4��Ły4�_�4 ���0ؗ�g�	��"YƴqZ����_�w���K]L%=��W�e9���{Z��,�.�R�p���$�������^ݦcه�˧N �ŧr+��#��-���S^d��%�F��=����ۉ$�쾋��gX���}X��B�o(ya|?8�&;�է�\n��a;v��\��EI�QAU� Q��,��Y�J~[ҏ+�	M�a>V��4U�Kz2N��#�穖еU/�t�I!��P0���TYy�p+�0Ϊ ��t�s �I^�}�m����bhY�����䩯%���Y����/<�� ��[h,�3w��0P�t�����%b�Y�>�:`����������A<X5<��bn�z�l��˃���p�U����+4b�M�1����Z|�6>�`� -w���Eܬ���9�Я?�75��s��C!�J�a@�`�$7����*#�:���� d�t:��\U~����߿�I5���?܆MM���e���wJ�ӣst�c'okM�,9���	*� L/�G��v�z!�aq-o��b�΢"����=p^UiEl:��*�(��A��(AR��G.�2�]<�D��	X(d	w�'�����������0e�u+�����U�C5��G�ڕ�S���؋.�TD.�~�[>����t}�#��0sY�9[x�L�^;fY&ķ� T��QDs�p���L�{�.���fw�=m#�Q(ewyo�Ak�n�@��'�sы�ξo 0-
��.3�^�"_	��&�����;j���(��q���%*ʕʳg&v�C�=��̙{^�S����	��-�ra}>�^��yS��v:s'�d�!��pW�jy5�Fa��9e��J�!���j�N�v٪�P!��/O���b띲�Yms�ɾ��&���q�-����/��a��1����'e ��H�~���ѳ*n��c:�@&�9��x5`cF��lo���6�'ʊd�����3�W�n���u�IIx���(��6[wA/�?���k	{�Z�!�SOZ0�.��!d�*ju�C*�ۺ�j\[�p��UG	����+$�=�v�hF�/Z����,^i�����]�T��-,�G��HC��A~�UK�R]���H�	.mz�о�t���,}C�c���uG6C���6td^���Vpf�j榙o��z�G�L5��鄟��c�	uʿ���$W�(���t�R�N%���[fҪ?�JTh&,ҧ�����������T�H"��ݕ�T,aC89�$N�`��F�/j���!e%q�,A��.ƚ�+O*+��H=5Ʀ�y�By�<�oJ}��z+���w@������S����ڲ�
"	F[�<���T��)��6CW!ij�8D� �:L�d<D/��' ����H�斈j�i�����tc{1�� ��R�C�c�zȃ9�'�d�x�ڍ�n))�kkMݘY�%x��SF{!z-7�	��Df�A���7GO`W�ﵣG,�@�sn &p��Wpc�p�P�E6�U%�y���5mN؟���*��_N��8:�J?�A�-��_|��xO�C����i��2�)[Ar�Yzq�472�
vwq��E��#v�E	�lt��qN��(�J���m�=�檥��� �Q�ˌ�j�}��AϷ���*Ajhdf&�'p�X�FSx&xf ��L���C�l��Le�+`(Ta(� Q�pP&�}t+��b�T\6S-s@�����ݜ�tN9���{+�d=V����S}�,X}���o�`�y�g�������/����|��BWX���a�ʮ��x	u_��e��}��T�d#������O��I3\�=Eӧ�G�	��z�a7��PJ�`$��4Le1\�?��A�@>oߢ@A����e.F�1	C"f��\9E�'C�_��_2e/���f�pi�"�MD�p�����g�u�kjn�C�%$56})mU��a<��t���Z�9�|��{o#c�Y\����u`k���y&걢��O���Z]z�0ߛ)b�k7��ح3�DO��-/B2�b-���n�*�����b�i��FI��[rV&&�'�Ԑ�+6I]� Ce�K�-t�BAb뼞�����~�(Ґ��Ԕ8��Y��(�NsЉ��V�'S��"�A-	)��j��#3`fR�w��#}~���@�w��J��F`2�'�m�=9�������l���Z�R�$]WȨ�%TRO:Б6k�����8yy\�xa $j�
ީ��`�_��tw���Zo	��e��(~� �K�Y35O��|��Y0U�������	?�a���\�%}�4�i�l�$�����(����k\/�*�E�{����`�7�ߘ��+
@L�:vR�(DXxP�6r�h�G��0@śt�B��G�93�$�8t�Ue5�~��H��(��{�lx�}!X��"�d��%�#'���o�!�2���֒�d�*3?����<%�N�y}�����*3���5�~=����	O�GE�]���:����d�fN*�U�*��܂�7 k��F\<�S����cgh0*�]��Z�v�����y6Mk#k��TC�q`����ef6�/�d��I����97d��o6����Qy�ȃ�FDV�
*CM�ok�8����ܱҙ�ʡz= O��;bwg�U�]l�{�"��������O����a�L.��n�Ѳ�4���	D
��	��m�F��Ӳsɩ�V�*�M}����H
Ƞ��i@��]MhG���ob��r��uͣX�T���J%ŪƼ�����/�*G�%੠
C=u�;�H�y|�����{$�7��Yd�k�V-g��H5�0D9�Ǩ� ��E
��tF�'�7RA�2��9�.��W�60�O'��G�mjuHh���/3K��qX�A��u1��t�،n�=/��gǋvwZ�U�qޙj�5@��ch�!��!����4��Ĭl�c�W(o~-d"����{^*r9��@:A2C�M=��cÂ�����ȼn���`���x��A�j���_A��s��@�����0�5@"���g���qt�����R���]��Y�'�� }p�N�*��uǜ&��A@f���o�OP9uS� ���^-��zP
�#j�rl1hb����ɕ0���7�Ӌ��HnBU���Q+f>{W�C /z��9�_�zU���x�9���ry�wS��q�C]6��੪���jX��
n!�c��ߡ_n����=9���;���Uڣ�����
z� �3g*��峌�u�T�Vݽ�ި��qR�l�@#d|��1��K��̉��UC����8VtmZ_���d�D�S�	�&��w黬���a�M����'��&ҼP@sOA�C�o������T3,ݧD��u�.�Y�г�iV�s>��e�ΐ)��k��bx�������Ҙ�s5=���3+T��O�K�Y)[������lz�ߏ�Z�hx�3E��:�kr:����2�߲@1��ˢ��&p�./��F)�i�K����>i�{������}1��H_ϳp�>�a֪H��JF��P@���#f���B�J?ƵzP8�x����9_� �m5F2�g�� ��oR�RFO�������f]��"�y7T*S$f�8�D�1 T��� _��y8��hbo:�T37�'��?�W����[�9���#W���;�x����N-���S�tʞ+�+���Zn�i�P���坁�5,���\P�bϒ,�
l�)_��ŕmC�7G�M��5����oF�ƈ���Ou�$����a�@�A�4�uKL�7�\="W�B��ܔ�Hœ{��Ie%��IU@g���[��Q�NV0�|��g������4OB	�M��`�ZM�W��g4��2�,�vЌ۟e��)Q�+hZ��1]g0�s[z��'1~�l�D)�"��0`<��͏ �o��$�cˬq�7"h�%�j��Ο�G�&�&�d�=Z̗{��ެ1	Kjѽ���3�n���?c�8|`4�K�P�EAQ�^;̘{�&Y�����p�s4�j�T��.�ތ�O1��c�ԋ��&��H�Aξ�F�5�<��� ÊI�|��xN:����p����ϓD=�����EG+=��<�m��psw���2�/����3��4t���.u	Q�EތTתh�9h�&`��'���i�hMA����ҩ9�ը��qJ\¡���Ur9`ܗV��8�[�'>��kL�&�O-8D>�ixv�%xݞb�'�&�{}���&i��%��� ��y_��P��aE�qomp�=��y��>�?6v�br6����FC
���嫻���T��A R���p�B�l���q�i�FV�Q�hr2��=O�Փ��L��=�I���j���xdd�CB���`�)t�#��J)���bS�o}�IF�Y����IǕt�f�Y�M�*OsH�<�kA?܃u��o�Ty)f��WH���{��y�pj�	t��'�]s��j߾>������=��g|be�I@&�y�ᢇ�I�Kπ5��f�e���43~�&�*�1eJ�~��Ь_�	>�+sd��M�_/���� ��p�M��G,HP9��l!?�͕	����;V[o4��IV�twv~����1����54Z�-��K�Xnz���ia�^BAb�]>[QIv)ᶇ���Da�y_&�y�f� g����5Q|?��^�5���v�H�t�����p2��eݣ6P	�R;��")�7~���h{L{M,↕u �^2.%��-��p%�=�&wS�\0�������� �ڌ�+�/�[���ia������U��3k�8<c9w[�B"^dS�b��3��H�v�<(���:|��r`f�(L��+{Imo����������2}%-�.�'Ygkٟ���kl��͐V���ԉ.m�*����#m���9�͗���t�r�$��0;�w��E���}`���p�&�U��Hļ�8�=�:�3�9^�L�g��rSN�C��`��w/1J�����g�d���qeͱr���Y[{^K�2*���� Zq  �=M�R���Q�Hy z�x>�W��{�ߪ5�����j��SF�����$� �!N��8�ӮN��Ҹ�����m�?�9��ܶ�|��#9��(]�y2���|$_X<���&��\�<��D\��6��
ޭ��
a�XS��ɲqĈ3���On�������,5)Ǌu�YWXt[�)�#B;���1?\�L]JC�!}��x�	��~�V�x�	Ryy���i#[JQ��L�����0�Z��C[+<���M�T�}Z�fuhfC:�ɵ}	W����_�L27���
]�[�rk����q��6���&**l4��ot�z�O��_�1���"�3J*Qtb��)��'�?�n�_�$�.򚗦$�u���i����}!��;�D-M�yS�rP�C���=�A?9�v��{�N�n�3�E��EP�)�n�::����J�*����N$�g!���H?Iu���	�)���8�����FY4a0�����d��bz1�Ł��J�2	��᙮�d�4���d����c~�~�,u�}�n�^��S ��J�!�cL��#�.1�V>�fR�����;#���iB� ��T�P�n�H���PC������>���	?7>.�Y�b�����h�Zt>."H��f�
"vkс��"4���`'�V�v1��N��]�
�l����u-�"h^��?T�i��J��~`g�O�b=�b���� ��D.��Y�Z���K�`�u��m�//�5(�K��o��ƚkjIfF����R�����z��Lq�B��~�`�iB��FS���R�ig�����WYE>5+�2'�-�����%$F��BR���b�X-IG�%����.w�c�T~���K��Z�+�~7Rn����e�>G5~����߾�)E��wNe4ԝ�.�t3
���$�C�$��+�Ȫ�����ڥ���f�R��Q�M5FQ���o<�ð�ꜹ�vi�E�� u��Z���X-���\
H�Wa%LW]�rr�s�73��0�b����?%�R����#�n�����D���w��ͨ:�	2Oo=����J�u�:��p�U#[>L���:ɝ��f��[�>Y��]�&*�J(��O��˖zn��X9rG�(~'Ɛn�仯3�m;�)}�.���7���N�3�^���t��(�#��0��`�G
u1� �k�&[��ne���x6��>��ķX]�/���䮭Ўͥ��w���.���m���<���
U)��W㸭�U�~��Kes"]cipPm[��ֶ�J�������jY��n��X_l�:W4�<$
��i�bCq%�WĮ�$�Gs�8Rj��ѳ��	˄���TKa�W�;s�
�+��k\��x7y�V	��:�����Ii1֩s��Պl��s�����띤��]"�'3:�1��z�r�D����7%/a[0��`q(�{�A%WSEu1�G�y{��&��8��+��ws����vx�rGbd�sˡ�;Ep%NlIZ���תx��9���K��gT�:�J{.�`�D��g�}�C�,��rؗ�P��@�F~�ϫ4�E�,!��u2\����Y
����0��˩����Ȅ+�?��JA?�=�\�a3�n�|�4�<Q�[��r�oQN���ט*��k~�H[��(�:C��c�<��5� ; �_���>6A��Y����R��Zr+^� IvjF�X�@�l�#A�s��֏i�1�����u'Jۛ��7(��Ϯ�t�}�R��j"�"�����zc��O}�T�`Fڨrt��M~8��ו���ި
��(JE)�����IT�?o3��U#�z�Hm��_�J��N`��.�z��>�[�R��@yL�!�a��X�c:��#�ٰfո���$�}�{�N����®I(��oԱ,l���3��a���Я���.�Z?���%�Y�f>�%�_��1'�}ȥ��#:�t��Ȗ�I٦v؂���ˢ�s�:��쁙�Uai!�6I�|#��F:��l��K��� ��-�&U�68oeC#���x�qYt,E�D�.,�X��hG
{U,2:I��=M�M�$/T.2��mPps����ò|YF6j_Np�!�0?YI1�H+��VKD0p�^�ܑl�}�;��x��y�O+H�R��{&gz>�4gEd��K�ٞb������T�Ya�u��C�Ѭo�B�L#��h���: �<��������|���^*h�M¡zS'�i9�LQ|ap�>�R�=J]���J�;�e&a��pY"|�8��*Ҭ���%�ds����,^�_Bar���t1��#�������|�8^,c�V�%V����Mi�~�-h���� E�ekq7�⵰����+��)�M�)"�P����2�Z�q���ϻ�ӻ;-�x!�[�:����N�0H��{�����k�A�k?�P�x'@�40�	�����[1�6ƹ�Z��F�9X�7��g�ְ+�0�����]
�E�[���R(l���{M+�m�)�~[�9��j���7�7r�v�,���s��wIonE·�/A,랩wd����zD�5U𧽕o,�T�z�Uf�P[�W�z��~Zn����'�2b2�GZKs ��.��K�C��X�J��O "��Jl+��ʂ�a���f:jX��㊀aq�a�c�hE���T&�ƞ��r0��O�i!&���S4n(�y����qg��[������n����Es�#+�Oh�pvH���
m�Xb��O�+V����� ���L'�K����*��f���}ł��]!�&aAT%_�@�qi�g���
A�K�+FS�3�)��P�2.��d��@2Y� j��H#�'�$wX��Z�����o��<M5�fߌ�ؾw��~�]q"���L�� ;5�F,�e��Q��rS��4�f@�F�G[-�] �a*���7���l�
�=b�ײ�;+"���s�;d��7Lf�|� �is��!��ī�$���L=WCqϷ״�����1�q�_��'�W.�ݧ����K� ��n�T֙p$�2��&�F��=�!4D�)1:P����
�����]pTv��y0���rV��0�fOhP�n���y����ń��vC�I��*c����d���C��9q����b�Y�ă:V�����G���t;�n �+P]��Ok_�=��=ng=6����f�Q�@a��ƪ��V���w�0��}���xU��KpD
�scp��}t.��rg�%�q/�b���X�{zi������^�`�a��Ң�)�~�@^ᄌ����a���|�Z�9;�yݽAU�	0�k:f����t�΀�\�>��1�<�䢕�� DܰB���ley�^s����_�
���6���_)�&���`g+K�+�����v8`U�˻��6�pB[������K|�^��͑1�Z�d�����C7�=-g�����ԮڼSUJ�9�H\� ���z)�<��&>Ӯ$c� &[���\�5���h��x���% �G	W��E������ڋ+�L�G��TE����ͧ�TH/fj�q􆴇�y�M��nX���J���#)�zm6{�2\}m��u+x�o�E�ep�S��KqFwU�7��@>67ݾ=���P���3�0|�b'�����Xyظӄ�S��,�U(\��I�=Hc�Y�(�E��S�/��=��i�F��n^0���|�`�r�w����3x��PS�ۜ#��(~٤��Cז��'6��Q������۟���T��)�f�1@��=��)td�p�Y�P��0��g�[-�b���P�5�.��e,�M���f8�go��C���ʻ��O<|���ZX��$����fe������aa)NcZzm��HQ_ܥ4��;�s�7��ek}��7�D�t'���b�������d �R��"�,(p��~s<�y@�#�Z2�f�,����cB)����!(��&��]'�*����~̂��V=�H���i�Ei;N�~8��w*��G�4�YB6��Zk3�t
�I~��-� ijy}��k�O�����Q�e��H�$>7��×�a�	_�wzE�\�!'j��%�%=���ԁ�L�>!Y&Vx���Jg�{,F��������$���m�؟�
�8���djo_Ni��k�`��i1U�Z���,�1����e�-�~�1B-�Φ��,��S0���%����@y�.$����;��*����H'aoP?�o�o���˽v~�I� �AE��G����3:��:gmC��҂�����Y���{m��b=t� !ȇ<dJ����	�J��@�b��f׫k �e@
Q�|a���T�(H
�xB�%�9���M
������y�Ehb��c�N=����#_a��R��K�����r�SzU�<ڼ���U�%����>@qG�I�&VR��C��yޯ��ýQ:h>1H�l_����#,=��W�|�zF�Τ�f�i	-����F��H]p�X��l��r����%�=|�̭��)MbujW�??�O?c�6����!���!@p^�;����ҿ¡��LW5�>=ϫ�n�
�~e�m�R�wok���}�䲬?�J�Ԏ��߯�Xf�
l2���ke'C0�X�T�k��	���n��JA$3L`ze�/� ;���+d�9�!�5Дd�,L���H��ڪ<����1���{0�@�-t��'~.�{ڣ.�Z~>1EB�nΘ��a-+���Qv/8����1����Jw&���A��/�J�XW�nT�9(��j�	�'�0��>�)M@�<0�[��1Fl�ƾt(J)�ԙk��E44��ij�~ʡ�2} ��*M
�w�q!�-�şA��S9+����'���X��z�z��	�W��{P[��Z�LY� Le[�?�ؼYJ5>�V$�(�"���$`���c�{�5E^~h��A��xC��;fb��$OUwE��#�#ؾ�OeĐƊ�ʷ����X��[c}�j�ܱQ"�.�E:?{���G`��;ʊ'�ўUy�K�����>�a��6���e��y#s���
ޖ�Y#�bF���c����;�	;�Dr��@�;g'p�k�����Ӈ�lD�{�v����G`z�u �<��B�>�EJu+�̧9~�34ꎃ���أ����F1V�a(�P�qF���{	���R�k����>�3?$�U��:���F"��s��?wY�J0�������V$-�m��g)C%֯R��8���តjĥ:wR �;B �'Pʇ�0C��B+�jz���2sR�	n��p�M%R��ʗ
_�g�D^7�ʬ�5�����n����Y[�F�t�I���B���YW���ӑ�)�/ݶ~�=^�l�2x�=%
�m�EjL��+�}���6��(�5�C���щ��)k0��+�@��S|�h�$&c\5���b��-,��yRwڊ�xD�
��'�:�1���:
C�pO{X���od&ExT���P,K�aZ���~B�h�D'K$r�l�E�6�R2Y{0	(!�~����΍9A�&oŉ�@��}Fx�?��)Bn�!y��R/��sm�p�% "?~JO8v�Кj2�\��Ne@�l�V6`�ї`����x�������o:6=G\�Y�m���d��C\VMB��$�{�/�9K�L��n����ih���I�6�n���n��d���j�FI�D�$"����e*�x���'Hk'6ty�|�87l����xn��/}G}Wwp`q�+Eψl3J;q2�g=�ʤ܁�qH��3�>����y�Կ���eKɻyY��b���*$%�b%�-���:+�3���BNp�ԛ[q�T�����U\Tt|�3�)��GY��'s��^H�m�܁@M��SQ~2
p���^���l�[����H;�p�Y�ө����j4�X�Ɉ���La�2ǤK���k�eY�S܂�B����@��4z�.�ˎ���憆zЪ�K��:��e���7G��K)�Z��F�u1�h�uy�D����!��w1hcTJ�N��Tj�@��<Sp�cI ��O��	�is��[��o���s�r�3�C߇"���tЗNJ��P$�蚫���$�Y�I����fp�L�pjR���[-/�?��������ũaX���������$rx"�'�K�⭛��w�e ���q�3�9 	�%��U�2�b��>~�d���9�:CN��:/c�1�`��G���X�'���NH��E�O� ��.����P�����鹃wUQy�ŭ�)�?��%��q{�����s,��a��<B�h��g�.m�L*�ֶ�s|i��{��M�VMD+�C7;@MQ�#nl/z�"Nb4�gs��1Ξ Qf�á�������?�]�+��ĽL��$��p�����i܆����$�<j�[�b�3�R ��U.�u;�7�u<���C���i�u�4v���+���7Nہ08mS⨎��{�p!@�A#�,Ι9���H��Q��c�%4�a�Գ�G�q�`�P�q��]�&�ջ�V�Ö�x��j�<w$(m :Q9J�!��ᔑ�B�ѷ��psh�mQx2�*�,=2b�P�Ln5�_�k������H��,��q�誄��7S���ӄqpb�����)fs�c��C�?�T�K�-�ᴒ�&t�d����f���|$e2E�8�n��<7vqW۝��A�E����P1��n*���+P����{Qr}䰤����[B�$�k���c	���	jm�S��ձ���B��S��|(����Bx�c?p:��B��P&I�� `-� �L�3TR��yy� _�#��+��@�h����o�����V(�f�\z�MC��j<'�Ls/
n�o1�������?��K0k`� �<+L7��c���C>�����OjU���Ε���/�7�^�k+v�.�#��tG<�:�U����VN�"ue�q�����������UxK�Y@`�~=SgI͞�����γך������S�T �t�R�/��oG�?�4�����V�D��{��<��*��}2�3���g����[9->~�~�&����{U�#��]@����aIiG�o��N[�>�wk��dtı���V�;�x:SL�b�?u��Q��9RU�y­S'I*V�B�D���QIK�Ԭ��WS惕z7�����8&���Ѡ� ��OvVк�G^�_Z�B ���6�n�A��p���������
i�O�C���6h}_#j�-��$�0r��aSWlv�ؒ�ch� Kwh���x���]�$�s^��Յ�;=�
�{����;{��9�G��L�q
��(��_��8p�،����c<8�t�]�*��2'<>5�7K�wC�e+����S	��X����8�O�"�P��X��d�M�>�i��l����#~��ѡ�C6i6[��s$� ���!$�W-m����Ϫ�h�BY0;E�W��d���M�y��L��O*m��[R�C0#���	d� �t<k�T��N�L�CUWk�Lv����Z�-o�5'(_�2��X�2�`CL��_�$\̆r�O�b˰��G�Ӑ&�o.�zg�7��?�;%�X�I�c,A�-�M��Âݫj�4n@;���u��5���$Z�"L zOD>x�ZEL	�%�nZ�;'/<���us�4�WW��~e�Ӊ���Y�b�YS;�//絼�5����2 Z��p4�5@V�o��e2�A��:�s
�
n$�uq��/�b��|8W��fW�5lP�EX�b:ysE|�Z��`��˷X�^}7���&��=����PGp��G����ܿ�����#�$-'x�aۃ�Y���g��:�F�V���&l�hS�&c~�L&����j���ySM�T��Q�B��jwU�x&����4��n�`E�"!��V��
�g��8>B�-y�n��߿C�7N��S����[�&Rr�������)��ԯ��2����P74�n"o@�C~�9>��c%��]Y�a`���y���:�^"�:Ew-t �j�,�B�R?Q��A��h�gk�HA�@c�d������8�v��a"��sZ$��҈9G%E����trwiӌ�+ǲ��e���W%4�����'����ۭ�5I?xG�Z���
��$�u�����C�=��@�͟�J[$��>I�
�Qv���J���~b�����$?�-�23H���=�1��[�2X���y��z�����1�Y���7���ok�JYJ�	�T	�hŌb%���9����VK9�ƷE��l<�L�#�?�͵]M�Ic�!��g��i�6���D�-���8�F�{��57¸~h,H.
΍ �yL�4aVA )O8����ܐ���0�Ikŀ��>�)�Ϝ.���t�:��׏�ќ����追'1���ܮ�vZR6s��N�-૭W�ѝ��;�����t�$Q��A�ЀK��j
����K���'��_���~R�-�tyry�����'g6�����rV�t�mņ�]G����^_��MXv�,�j1�6��$��������24u�v�{4�
۽:wj̨�r�g~���0��jc77M�|r-"<(�����
�`��Tw��2]+���8���[H��� 8��D�^��	�[��F${$��/w��	mBQR�c��D��,�k6�T�v�&�f�.8[��kZ�N|���2V\�Z
�꿄���綦:ky2ۈ�8!T%���bK���;�;�g��ز�ĝ��H�0�̧P��9�� pz�p������K|4�E����`��8E��Q��a�1,
u���c��~�d:�OS�L4R�m0s��߸t�Y��,�E��ִ�%������(8�o�D��އnty$��0�\��wEn���1���^	�;�6���B��Z��d��rs���}e�^���cp������O�Ȇ�tm�Ƥ��������J�e?1/�'t&{���(�B+ȹ��0U�D�����6�}�8��m��" O���DJ*ѕmш:-t�vh4�<�O��J;9��t �Ls��Ҧu�œ��H�����~*s9�:��&��K�p�G"D�&�S�34OR�3��ڧ�h��U&|�r�>C�����I>T�#a��K,�c��%8!*!^t���B�C�-�X}&�[[|�S�U�Cњ�Y�]P��N.L�< D��ynAu�% �� t�ufM�Gk [PU�l����Q��|��k���,@������ A�k�b9I�#��k��X�dMp&1��yɤ�}���!㻇{��V&�����$���nVWʄ"~˂��N�������7|�t�<��#K�Z�4�I������JmE@G��by��⤌���G�:�ᚮ�OV��V��i�g?� �	�_)PL�{�ʙ��E*+v���[g��O�x�h��[lNS�}��a�=�Km�iS�{�H�`2�JE�Ja�Q�5)pH�4�%S}코[+0h�nZN�J�E1�BW�͢�Qa�'=���Ϋ�|@�U���޿V��(X���j
��	�Ƒ�.�ϭm1�ܶ~#�N*1u��w�&^ƫ���/��(�.x�q�
c^=]J9fع��b<<_,�%�Gp��L�p0zA����
�*�y�1��ф�|g�I�_&y/�̰5:M�|F���%���J�H��h!SQ�곙xgx��;�=,�C��P�|D�r��ēnR�	�6?�����n��B^b��]��⋷�vq��.�)�L���w�%�Q6���z78�gR�B�:(�:��ͪ�\K��]�m�H� �|�v���D&?댇���"��h=ʟ�RC}�{J!~G���f�Y����OA�3����6����O� \��sO)����ǰ��Y��T�8�:�a"\����\R���Uw�A���G*p�R�Yj�MM���ƕ����������(�C�L;'�p{�4�/����ir�V���0&	� 6D3��觼ұo�E�ڗ+5�\�vJP��J�_�T.��_�90�c�y	,�,$˃r��E�@=[�;��g60����A���6�ˁ�e��$����f˛յ�����-��Ȳ�����,]���d ӌz�� 8���]=��ByU7�@�`=aJ�EH�y�~]s�=za���e�����
�ʱ.�q2vپ����ޚnO�]���������l��>��i���\���4����"�3��$��
u������c4�o�q�K̙�>�	�kז6�Я�D���E���ֻ��!s'K��'!f�[՝#U_`�-�j��?/ �此M�8�xYXD�ҺU�|p�}_^� ��:��wQ\\+���S�A���V5(K�o��.�M�?���qv�(fעa�k��U�7w��k�C�v����4�Uc���P�Yz�U.K��s8Tӎ�g��Ҥ�4?�7�m=�ߡ �bJ<K���y�N�Ti���)f����\��t��fƫʳJ�*�[�9��D�X��pT7���Sd�S�J�x��
�+�?5�6�,^r*�^���ݖq��0"��|P`�$��xn4�X��
��7s��)^i�Y������P7�;V�����Ry�7��`!��"��,cJuK�ʏ�7l칢�t�!Q6W
����_�;�������`�<)���f�ard��	z:�+���;2�S�G[ՄHy@��4 �m���(��N�£���arݬÒiU�Åh��P8�0,��G�<q̂���; ���e��d����� E
e�=+���aύbA6m���`趫8��� �]ƣ�-�*A��9�H�`�L���[�/�&_�6Q'DD`�.r��c��HM��n����4��\Ʈ���5d�?4k<�(@d��r����0�����T�kԄ9_��;D^JK��H�W+p�-7(������{�xhř��&)H��o���׊�b�hW�uHdp��׸������(q���acA5m�H&Zib5�lYy��ڃ�����9}ʥ
��1�L�y�r�2v.	����HX���ܡ^"-t�pJ�e��'�FF9�l¯��俫��k�5���tm3	����z���^=�YO�E��AE�,����Vv'N|�t1�����{t͊j"��]h�ؤ09�?��(�����>$4�������ca�5�C.-eHO��?�����@�.U�
k!̏�D�J4Y8�\����?��_0�����^L�!�73/��n�����J���&,	"�nj��`�B
@��(�)���b��i�3�g�o޳I_�>�A(+Q���dx��P���7@��i��a.�w���t��}�;$��eg���>�!�&���`����]wL�vfg����꞉Ѧ)��N�9\�Y�&��X�$P�R�Wo��2 B�;�>�{T��4 ~�IG0ݴl�ʚ�M~	n<p����$H�?�O���ѕ���<JG�xm=��9�z���Z�n���D���eSov���M]Ub��3����M��*y@�cGϒT�b!D)ݿ���o('�C?I3��W��2uA��1���D��|�8W_n��Dh����J}��n1��6��TQ��׸lH8t��]��ypF1�O-�&o�{l�w�V轐_�5�F�v��\ �K
��jتe�E�H�{������Fn`�W/�8Y_G~������nX*I8J�Y���Q\xIJN,�u%҇:������Ь�J�)�r��p�`��X�a�U��$�={"IɎ�[��yk��_K�uH�i1�i�] �p��jf�X}nj�ߐm�vBiJ��hd�7�'���2�Ѥ�0 �Uo`����Ic`@ �2N;rP[��I���wJ�7`j'�J�]�]�Q	��_��4����z6��ǡv","�g�����2��;B��~`c��T�����e��P�pH׀�����F�N���X��O��"��ۂ�Q�S�b-?�_�I9�}���8o眉a�T;�K����~�%+�E������/hX9�i\f�)��C��9
09,۩�P*��z�\TG��t}�`ݵ�I���pb>7���;�p�]�&���rΒ���6��7�H�u`�u*�T���'���s�,���5Ƃ �H���A���Ƶڐ�*׾1�NIr�h�_h�k���4��	������Po>�V>?LTsG�)�o�7rf�/Q���Mg�ή�Q��	����.`���G��N\�RQK䘮�����j�s�=���j��$g�_sy���A� /���gͫ��n�݌��[X��鮯�v���cQd��D���p=��e��m
��ʞ�@�r	թ
�>�<a� ^ɬ,�%��s�2��[������%k����6��>�9)��Ϸ2ll�����l@�ǰI�$Z0�W�ջ�;.9�I��q�5�xh2�Ё�����u� <��ers<@<,%ջ kԠu+h�G���?��$��A{��R&��#�i#�&3
�o�"-{���;yxC:��ZY<F�O��H���"a�ZQ#LΗF���ͷE
\�0�;1�I��w��N�����2h�NZxP}m�ԧ��]j�{�̠V
1/��8m�~Y?�M�E��J� d���g�_.;�,5;n�^��oDA	��%:��F�
�j|@D��h�#��rx��jOb�m��|��H8���� �)FM�
j�BV<�fr��/#��]Ba�g�N-sL^�k"?���縲�[�r��v������D[���:	b�)ȏ�o"Z��l�nm�8���� �P?�x>�;�R��³xJxe���U�X�|Hk�� ���@M�n���Q뇠}����/���ÏLX$�k�{H���-�A�;��T(�u��sI�B褧>T�=��1��OHd�SdO�̡��d������I_��=���kh7�lI|"�� i�i�IC5.e��H�.3��RIq���H�0�)�2�����N���%��n��e���[��2Q�u��VW@X��;��)2�����A�p�Vǧ=�:�9�� �@�V��D��M�L<�Jk-�z���H��
�{3��̀@e4į�Pr����Q^�:OG$RL��� \����ޕ����6A�[���qB4fqjA�>}�U��SZ����`SJ�Hv�Yf'��~�2^��
���W�������j�w�q� ��Y���|)3|M���"�Օ��B�,?��j_��]���uH�_�����Б�����pz2��9Z�l�NS�'R���t��25y���g�\U�Ξ(r�2Zd�Cf�r�D�F+�l�EL	���җ�S �0��I�rV�/T`乚>#�^�*�z�M��	�j%�l��S^��#a:�.j�iș`�m�]>���Z�Kt���Z�vtv+v1�	�nͻ��,<��p��6^F�ք`,����+b9�$E���*+��Pւ�΅��P�;qj�q�3-jK?�v���'�+���������>�O�:����<����WI�sZ1�+����;z'rGsH�@��N+�R�w��q�K�U~�
?=YDv����ZP�\C��JWyY���U�ڃ�N�����պ�րI�xd�O�~�����$-�*̝~(N0N�����HdS�F�����Ͼg�מ�{wqb�����΄��-���<�r�*���T�Ƈ��(�F�C���8^I�����[�yK���=��Ժ�����w������	��*����셪����KEeW�e8|��˃E#�e��W�[���FB8)/1���=�0�����G3o�F�)X)���q�Y7,��:n�������������%B��S/�LZ+��o���fڎUট?ڥ�Z���6��@�լo%�`��2
V�-3^�Ė����Y���v���ׇ'�G��S,?4-�	���U���T�����AS����oЩ)�lƅ@��"�>TB��7v�Y
�|g"�z�*�򑽭	2�U���ꗋ6	��z�0�;�HSR0Dh(v�7�������������b��d8q�挀���uz�˪d
5�],���'DG�-��1�hh�X�
��\PT˛��A�i��	�V�ڧb�{@F��K��^�e!5ҿ8 �ͫ2o��~�r_����'X�>���W�Wm���HƺW�o�x��"�G���A��j����ㄠHvi}�HN#i<lO��/��Z�3�9�KA{�IP_3��v�IⰨفHa�Aegq�ޑo��p:���11��I���ܲ��g�St�v�w�vu�O<��|�׽��)�^z_L2?��2�@"J�jo�@�>%`�����[a�B���ys�-I蟒ߍu��h��]�� �F�L�nl��z�墤7�G�7��z���~&��H��t��i,�Q#��<ʍK�w��{r��q�thh'��Q�	T����;�J�2��4����Z�4<7!Mț2���8�ž�����Z#�F�w�}1M+�0�E%���-�:{��]Q�/8G�k E]@e����(=����y���J��b��5�F���2��I[aI?Nܺ2zŸ�f� ��Z�z���o�y�M�z��k��q���2��z�a��榺�^�r���*[E���oؘ��m��m��x�{��R���a�#,����'������QԱض���bk�����Lɲ0¨��,L{���P����(��f��B��Ɏ
1����i��XK{U�ۮ���!1I�
>D�d���S`h�Z� ���5���(I�3�jvav��| \"�x�f��ۏY}��o��3BcR<f�mh/���F�,��@�KB,��t�����4��ġ�`A��<���I�l�d�ڧ�?M1t)���y6g���q@��	#ܳ0?'}�@l���j���)4��eW�6LO: y��Pؾ��sꐺz��� ��*�L�]���O�1��<ĬX��qp�ؕ�s77Lȍ_a�Dh@��ϸ��Ԧ��a�vG����qY:�L���;;$���c2̀`��zk��O|��co������道��7��p.~�AZc�^�6p�_����U\i�"٠y����?�x�s���t�0��63�G��7MN�7���b����Qk��
�������3`�oO�A�]z�!t۵5�sKʔ�M9��J�g_%@��������f���N����A�vk���r�Pmw��A���`���/�8��u�w���x��>�J�L�*Q�V90#u�m�ܛ������%�
;���/�I�ۜ�x�yaL:hfTX�Z������VGw�$>G��K��3��=|)��n��V&��SA'�f���#,�W����
��R<.ojC(A�M$ �0��1����7e��pyAIS{&��/�N@aPG���c�ɓ�N:w��r����΅]�w�0@,<��8�ָk�	;�?�"�r���%iR����>��CU�)�ݚXrO-��0��靉pw�����w�"����M���J�Oe�
�'9���t���fR��9���+�uC����ct���K%]�ekxe�� �Z߮f	+�TD�?�Ͳ�$:�+���?�W�E,���M�U��z����'����TH�^@9h��N�����m�ƥ�xD�ٳ��s��͂�5R"n��x�}��~X~�MY�G'�Y]�pC�[4q�+�<�c��v�����Z�<�o�EZ/�����h�x"I=L"�A� �]��%�C�����N�p��&xlo�E�E�}
.`�4�	�I����w�*�r������:�k (/����34]Bo��-+�&���K�0\2�<gL`Z0��+�
�.���8�	�U���Þ��m;{¸-S�4+}B��a#$�8�t�P�̊�}�����&� (d�����Σ��O9�!�gut�=�$��SR`N����8+G�~D.[���4d��7����J���*��q&�}<LW�?y� �M���(�3��nED��ӈ�lQ!��WU��#<������Bn�V��@�eXFpz3h�Wd�i���yH��8{qȯ
w�ϳ<=,����,������($�@�.�Z4� �`�t�9��m>>�O�rKF~<F�P�W��V���`�.+>�k�W�bW��to�t�{�e�؞�fVӋ?�����v�J6���53��l�읇��ү#Y���:�{K�0�b�Ԧ����>��ԫ U3��5q��1�1�;K.�q���\Բ������Ew3��i��|���pc��(���5�o?G����ut�FbQ�4h<G;>�\@g�G�� ���gϡ�i��i~����߀���'�)����ATQ��M0�*S@�CM�B�,ޘ˃z���Lk��?I-pE<R��ɫHW3 de�uGҦ�?�M5e��F��1�Lk��B��o���˘�A*�f��3�81�Ă���Ĩe��x��R����X���DFo�uo�{�]2e����䚚^����H@.W?��#x�
!�{5b@�� �Dl?��6���ndW3Cn�w�Ĝ���#B��{ !ҥ�b�w�3̐bǫ>�[Ȓ뭹��=��������_��EQ�E��^���k�8��r���Um_�kf�Q�!K\�W⥔���B�t:D����^SecGb'��L�k���4+�#^�qݥ
�Ĉ��U��k�X��)ў���b��G�L�8�,J��0� H>Uy�4�9�a;��SV�6�lB�:�N"��H�!e8�2~.�u�N���\�[@��L���q!{xUj�`ӗ��~ck�oV+'ˋD���w���?�ß	����X�ք�-9�)z$� �(��.����ݪ�����ԟv�p�����j���6��B�nT!���+&�y;�r��۸���!M�8U��� /�Wn�<!�}�0�T���k�;�t���3e�V^E)uT�*�UXT�Q9>�#��X?#�!Rx�@�LX�b\�"�x":�s4|��܋������l×�_a ���R��a�iG~�N�h�u������	�P`�������c�&[h�#Ѣ�����Y�H�������UC���T�4!+������
�wt�c:��5�?��P�P�u��l�W�R���I?��I�����[h	�AR��b4�Zh�g�Oƛ��k%��>�r���q#c�A��=���W"7T����=�ޓͥ����c�j�! ��J���(�zC4�V�ɢ�t��� Dȗ��Î!�@�׫9�]��Y>ܡR� l�W�n��;��O:�L<�<�����hޕ���f��&7���_�iO�-��`ӑ��ׇ>�W[1���S��O���e6��^�G�NK�A ���'��@�#�)���1�J<f�yR����&8��
xIq
t� o�\T0>�t�T���N3Q �C{ ��k�Rw����H}���D
0�s�mW��s�A^�_��4q��ͧ��{�6Ϝ87U:��x}��O(�i���D��k����c��ǨU�`�6���3�b�%qBv�ҌRP`��~�[��0'�n�h�i	(�K�`�-���,�*��m��\�a�'a��;-J�������M�6���J��w���_E�"�|���6'b��2�����WƠ��ߏ����,Ux���D�;	לhe�Y��Qw�t�����z[�L�=�'TP?P+�c�-�׃��.�y�ʪ;�֌ ���S�=R�7�����r3��(���l��^��f+t��&�ctҏ���K�}�m^-]U���Nv"ޡ�W�?ֲ�l�"���Nr>������H>z�ш�>�V&���(�m�}����852o��a��j�������(x#aR�1�6l�C2`1�C:Οj�_�>��D��z�Wo[��1�6���:?��1�E�@���F$�d�B�Z	P��ŷ��E�YEH��s��J��3x�kq[m�� �Y�ftq�C�$�	!����L���6^���W~O��kWq(����3Ú�N��̾7���|8�2�ה\ү��VF�j�5�u �]l��"+�U 6�%B�ן�x\ �*3�Є,7tf�0���gr4f\)е��T�Y{��,���<��ZH%Y|��7A��0�z5�ϡbx��N#"!UY0{���,�/��:	��yǽ�|���o1-@_Q��>�ƙ0$s��B�͊�Й�bٻ�"�HE��Ap�eO*�@=����$_p���B�,�c7�#�8��	y�a��O��=�^^�e�n�۵�|�����2! #u�p�.��N�
,�r�p���5F���M�UU�\�bd8O���b�,���R�P���I~Ќ��q�5����ϔ�Ԏ�2�p�°�'�
���Uv`1i=�*�JctkH�C	]��,���st�`�D�� �`�N�|��a�����$�v��M���x��'�{�ѡ!$�˺�j��N �p�͖���\�@��$��jG���F|[i��3^}<�y0�����+��G�r[1ݑp$�;�4����m�3��\��}�{˻R�#�Mk	q��ڜ30���&: �Kݜ^��w_����#�]�tL�+W��;�P݁g8y�j �Y��}�lꥀ��B,���,߂R&�"���~��Ҏ��E�v6��p� *{�t��SJgB��ǝ�-�I~�g޴bK"��`���*��cm�S�*L��V�WU�bE�H�I�P�� �V�E4�� �������g>���@�Fއ�߃]
!e�v�a��Z�w�x�H�4\��e�f.���$�3Q�떿�l�V=�!ZlV�)�{s� �5O|����V�N9���W�Ă̜�Յ��"�v�@�S'��w�G�'��m+��i�̓]LUw:|��`��.��@4|b�{_d�&��xMWp{���'kU6�����
C��A�<�y���W����Uoh���Xw�*��gS�;&U *�^����}��^�|U�t�q#�UO���xXL��ahI%С5�.�`�u����l�w��t�_�+C�Ds��hn��le@�ԓT�"��m��|�$WN�к�j�+�V\�\�K!��XF��!��z'�DK�hُ��@��E�Oi �>�ۉvѓ�=�|���R������}�=��.n���� ��6�$wXX7���� �^}���9~5�〩/V�� ��S��43&'{�hv������-�X��k�?��)�5��|>02���J�j����7"�ia��Eb��%OԖ/%�0b�՚�V�,q���59������n�X|�Ãk6�:R�'EQ�!�c>�e�+���� ����ʖ��Ɲ<,v_�������M�A,z�u��xx���Y�m�A�����[��\����4�c�&�!��2<��S���(�W�'��׫f�U��=r�8��Jve�70��B�e�G��<d�s�w���\7����?��G�,���.u����zdD9Ux��������gh�U)�����bM_�V���%?�K^,s�ԏ�v/[nV���`?��sƽ&�,�15�,y�үk��,1�W� ���	��(ט7��Ț`�����֫ٱ�d�5*|
w�+��:�%�"��T����A��`-�gG����'߈D$`��$���.�@����7�cI���u7�R"�}	�k�P�[-t��%����̩� �z�w�����X�������O;�Bh,|����;i(�ReQ:�v5�C���P�5� ��tk`�a�2m�:���ۀܦ��<:�ʶ"(=�Ti�W�HB���]&YeF��t�G�U�-��T�5���C�G�m��>����mC��iH5��Ӊ���?D៽]��p<Fl�+{�VM����~0Z�
�.���O����B�k2EE�Ӄ�� �S���)�q�N�x����$�Q�zI���E����DH�r������|�ƱR�����#5_�Fs��|�a����a���j��h�<�<��v9��W|���8ӈ5�I��0m��̓R�+p���
�0c�ϰg�ݮ`�L�+vt�ALyGȴ՚q
\�7i:-�z@hBX�.����	ԡ��8
ߟ�5��ǵ�����$�釫N(�f�ݿ�|(����Un�i���f}����<�bj\o�#� % ܓ���<��a-@Ti�j��� +-L��'��d����w�@���P~��%r|_�FF_Qy ?��6�D�Iv�٫�\'b��y�LV�	'Es^��\��"��d�����T/0q���sn)e���}��Lgb�SqT����zy�B�L���c��`�֝��I�q���H�O?�����Ƒ���^K"��l��J)ґ���D%dh����T8@�ħ�������}�{(�5���m�:)uQ���Hu��n&I؜������R�+��bX�b� ��V�t`O�P`P�����Ԇ�VA1�P�]<@���6�V3Z��E�
����0����e
�?6`E��
�C*�;���E��KG���5�a�)�Ǹ���y�!DsWG��W�v�����8#c�Z^�m��Z�YY!x�M�wC$��A��0�/���M�s�[��h#O{{\'V���xP��N��n^�Xp��j��("��eug��>�^�a]m�yZ}�c��EO�aB_���.=f�J��5	8]H_��q\��5=��g�z�X���l�M��l۶�2�$�����崟F5����Ŗ2*pn27oǪ��=#���F�.s��(�k|���.*��B��s@OT�R�,���(��|��s΃'�(_7�Cbd56��U�XWo2��mS�)~yl��Z-��P!���5��&�������K�0�[�5��\,Ȇ�\�p`�tk)Vފ�N��x��ŏQ�>��f���H�����^]�T���6KەFeR�/g����������镮Ū=�~�3{j��~X����C��`=�5)]?�p�c*�r0�V�X�:(u7�\�U2ׁ#"�vϲ��}g�~+�SM�R�%&��g����G��9r��~Ӂ����1ās��D�h�^����Z�%��^nف&4� �9W���V��ieM���Xr$jBA�,����hm��[j[�����!��ս�����"�䄊u�iM�+�
�kY�;S�|#���g����;��Q}~_��8�:�#��jR]re@�x
]���Acī��������2�[>���OR�U�*�9v�B�Jk�����6JU*,d��ᕁf��bF�]�a5!�q�7/��8`vy���Hf�rG��۶���WP��`�jv�:�i��:7vH����k&v%V&�1`~����FbXu%��/�s(e̋�֜����]_��t���=:6/�8*vhN�+�	�i\��Q<&�a�T˽�oֲ;���~��ք�.�]�n��B,��e�P�d��&���55撉V�H=oǉ���d�ƕ%��p�����a������j�X�ڸ���=i�
������~"xT���؀@�D��u�GI��S�Q�/��� �:�Oj�&�d�$��S
_���[�:+�WdJkY�I�s,��mx�zK�k1�= P	o��X�nY3�����93'�L�8L�\ri"��h
h��i<�ٺ`0k9zz#l��cg3�dy��k��xy;q���ӹm4{<����M�h��4��;�.��-sJV�n��X-�w%�(s���w���hh��8�D����<"�IILm��K�N�2���-sq�䡁��M��I5nO�O�uK_QP���(�XY[�����$���ā;�Ag؄����NF@hDQ^`�m|�e������M�������
���{|)3d ��n�cl��dM�R�x��i\tyJ:��lbԹ���<=���>q���<Nk����}��t���r�s�\��P�[�)h���i_�����0��G���J �譛#Gz=a�� ΒW�����b��m�����Ԫ�3�/�@P���s���Ta��!�v׫�$:/Ep/�`)-KV��$E&P@DO�����U���2P�"�c�ֺ]�bcP6����d�rU^D��/���Q�DPB\E�;��be����"���{�a�e���#��RtZ�������p� ��j�����-_Eu�b,�ʝd��p-�t�����~�+������tl;��V1�V@����\OI�L��헊Z�usFp��{�|�=�!���t�9)f�T��"G����ۅ[��F=�b1N��@�uE!Ay5�ooR4��zU� �/����y�����#�hu3�����ԯ�!?k�s��H�೒n �f0���Q@�l�M�b@(O�������f5J�XzVM��������Q�^l�l�N���p��v��S�W�׼g�oh�E�h�A����R�}������.��ӚmdU
4���!�ǫ�Q�2OC�Ӷax����(9��h�C��j_�����<��IK�=sb*~�8T���q�,�ā�=����.�4>�ܽ�7l�3본x;��C�3֋;���hP�p6�T}x�x�PEX�3(l��1l�� �)����\ i�����!��]��37%g�t���h���A�1�hS�W�א�6k�X�^����C1�z���8]��K.���~�R����l�foӞ�� �h*2N���lC�������������4�=�}��w�PC���-7�#�q��7�x�>�[�N.�J[E����v�62hh ��wcSх.?KU�<yr@!�EN8�y��s���}��9�3Cŏ�&3&!&g$�U������y�,��s����K�������٬����@m ȇW`D�A�|��~�?�V�J�*$[�J�q 2��4Zt��V�)#:7)�J��x���bmR)�f5ѕ1��������b��nc�����)g؂��������tNb=L��׋�81��Zgb�^��Ia��=2q��i4����c|���Ne���������`�6-ߏ�� ��f�7f�6S0����J;�Y[���"�ؾ�rQ�]^��$�/�3 O��Y!��1��&�0����n���j�L<W
��v��i)��W���o��m���2�Y�*�W�A;DSṭ�ra�: `(��r_�3�"�z�E��A,�j"�*���T�#K�)+��n?

8FQ�t�q���JC<lL�zO7�6�+s�$�U�b-T:�(؋�� K� s���}@���^�1_�TX<O7��k�~�ө	���:����.��U\��vU�'^M�cBe#��5/��rתB��Sgf	���3p�?/��e�Wd`88�4{���;�Kk�k�8��+BgA�V�ڏ�\��T����˒��8~k�M/:4.��@3����!��	��q�E�;v��p��4૰<m7�#�z�]� ܽ*(9%����0:��6]rA �튙R������{�b�F�>��.~�)�y�a��(�+�ׯif2���p�S�����A���ICsZА`��ٰu�׾٬e��Q�"�(����?��G���;��QPLD�`��c���u��H�z��4��i&)|�&�4���,��e`�����Ǿ�u�q�NR��k��(���y˥Ͽ��ci�6o*:ה��<<�W`V$�rO:��B�Y������6:6!���ܐ���h�ٳ]}Y�L֌�Eu��q�v�KNg�+2%��K=��;��^e$��Ϫ{}��\ ��uTɍ��uð	q��&�6jH�_x��N'o�a�~��ꇇS �E
;x���,���6>��Ϫ<1K��^r����_Kūe�����\tʦ��R�D+r}�"Z����$1ƙ�*��oPv�sz@VA6%ߵ�>y�����V[�P���+����xuiv�N&e!|�c~"d?�A	���U;/
w٣�3^�}ل1��?�7'�	)
�Ճ �p{,4.A�X`�z�0A�s���'�1�]	�
4�� �e�qK|�mb[����5]�����8Fe�9�	��c
�j��C�˿U�{?�3�>o�	,���f7��"[�G�ğ��`1��eT��f�j�ae��+��,���@����R\~���x�x���R3�1�����CO!F�P�����WW��2|3q��G�r:j-7t [��iJR?up��3:m1 P!J"rK��-`�@>X��?2���=B����*��/��"���Z�|π�����#�h%|"E:�/8)�	�i)^���^��� ���[^ɅϙPZ�)�B�\�u<
��@�K`��}��]RZwRE�'L�_����j�l�箅�1��c�|@�4�xG�V�� 6�䃇璽�P,������´��e=���kr?�c�mt����#2HS�(�k��(Kr!�9�^�[;�a�xQ\�XR�b)�w�Ƿ��>dcD��|
z�)O�J����|8�5^"����(Ӓ�8WAX���ԓ6�+aO��
�|A�@��}Mab�q�� ��-"�MgBM�ز��XM �*x>�x�����&fF(�I���KUpSM\}<��V!������ 交W��I�Q 8sRCh�Ka�*�/�崎6(h+�3��ഖ��]Q~*N;��E��5И��;a�������d@o�4� ��~� P��/�i�"�қ\�������"76M��ITI��#D�C��D*�z}��:��Y��[X��Z\��w���2ñ�`�6J�Vg/���Y��B��̈́$���B3!�)�_��|��j���y��E��\����X�a�W:)�H�f�d���I�VՠϠ	�qR�f�v��^᡼%�z�G�|`�n�~�9���j�
*&�G�ov���Z��Aο�q���K,���;_��Έ)�{��oXU��5�'����Y3=���<*���b��"B�o4���+E\��U����#���&���=d �w	y�O�s3G�����˟xv�`:�����C��&���2k�D����A6�ЉgQ��H�|��I䄖�7m,��v��Fa��
��Vp�H$}_��?�v�"��z�;	vl.>�|H 9׆v7��]o_lY��5�jKж;��@�#-�`����k�eD$�����Q�zW"P����P&����E���{��ɫ�;#ݾܔ�W��2�r�&*|��x�O�-i
|J�onj���!/}ע�Ӷ�J��5�'��v�U�~�/Ǥ��J��.t��i6�#��\�9���TaXB�<[Ӹ������nLK��!+\3�HO�$��|ß�bSX4�@gR�4�<�Q�쎕h71*)#�Nr-�7>b����I'e������*�Ȍ �b�m\g�k����x�H���ջ��6��E*bMh+65�F��d���Bb|?��G�LO��lj�ߜ՚����LO���S�@<�.��F;�Z&���_JR���Z4���sW��d��R��U�"`��/}����"� �q��B���OE��NX>߿����0��TA���:���k�ج��w�hw�5�Y��ɿ�vױB/�n_-��X��B��#4�I4���ZƦ%���Fj��xG���gΞWX�n��u��@o��)�g���>�o
�#9'���F#��`b�qHN~�ܤL�Bw�*A�)w!��)�<�h�G��w���o��/�p
_2�~�z��b���t�N1޵,�y���Wf��,���s��a��1Џ����`�o`]9*��~l�X���}<@����\$�3g߄�zD8���6߂٨q8`<�>�P����ϖ��7���;�O�vC�uz�{��\���E�f�_��(�&�['�>�D������m*�f�sG-����`Um�P�?N�T�֮�x���*͋&;6Ko���Õ��O9�4?�.m.X�ۚ�{M�.E�H9f� ��|,�UPm�5�����;Kpj�!m|t�[q�QS�06��c�{-� ������rH���R���D��6J����Z��%��M��~\�)��P�<�6��̫j�Sϼ�O�>m��ppn�����'#�2�q��f�{���έ��|~g�9 ���5.l� F<���
�V�fU
�
���a�s���|���X^�W��ف1K_L@�ID��!2�6m���ɥ����s�}2�j
�,���A�=�dT�Ē�a�l����r���Ύi~�U�:_޹IS����\�ؑ�%�򇅍���!��fpPmt3�vrx�	�����\*ՀW�4v�\6�\��VS��T̘���!��%B��zV�U�{�U���SS��mG����+�R��7<쌿;q�*�_h,_-N0-��%T�O3��I�����_����:|�`�̣.����vޏ~[�V97��sV��h���j�X���֔���~���i��(8��u���dQM-Q�s�K�Q�jp[����wzB�M�d��'��d�����5��u�a���MC�'����%C�x�X��[��*́��Um@9��
=f*�ԓ����Jq)w��g�"�����g���+��[��$.���~f����u�V��슕�Ƅ��b�Z���<	������+�/�K��H�E�>�YlL*�c�.����JB\��yO�<�S�f;5I�o��M�z��a�6�B��σc�]��>8�į� �DdliG�y��#:k3�Z<����v�R��-JaV����ӂDZΐnSc��Z�����:�����V�{+(\�瀵�'r��4Hn�f �w�%ی�(7�����e%�_l�kD��#�ڠ5��]+����-DV5᭤��F~�j@��,�x��6:Q'^l�0�Ԉ�������2��S�|VU^b;�vK@��.-�3�ޝZ!X��I��kC��ZHJ����'ԖҬ��j��C��5.�Y�H�����]g��H�9��x�hG��?���K`W���w6r-�_��C��-��%�Y�Kʪ��b��5r��\�w��>!P�SQ[�ڃ��b�lN��߯�����L��{A�(W3�w�Ə�ޥܝH1���{ԆA�������`*{�1��#C0�\�s�ɇ�`K���\��"7N�`��8֕��a���c��V�y�U��Q(��).�B�T��_E�U�\i��[w�.>��;¨k�g�m�҇�WV`�Hl�r�3�Ë��쫙�`��X�:M�p(2���rs7��E0��Hd��-��I�#��Yt���eڙ�V-�PP����v�c� i -���9o�]n��R�;@�O=�`�3L50�����=܉��C�^���a��N��㚀�o	~̍w���S|; ��7�`��P�4v��-m}R�r��?ygؒ<��tָJ�Evܰ��N�c�����R����e�g�"�z_ο�C����A�k�YŔBf�@Y�?�'�:�a�W��?D;�P��ӹ��פ�]�K����u�Rn��HFVֿ�u)Ԗ�\�.��)3�W�
ִ[�����o�ZD����c�}��?~~����4\�Jp�t,���r�uu��$��:���)L�����[����'��ss�B�4#�Ζe�L�%�Ecr�-P�=���ݮO����ߞr�8��(�����m{�>���b?ĲC+GX\)a�D��
5]��+=V�s=��k�PF��?�!�P�C(B�[�R��Ȣ��T�����PKlF'm����+-#�*���N d[e�(G4h�	�/E��^���7��ޤIy���C�)�i���<�X;FA���f��S�k�A���D�����E4��w^�:	��l��hx�"�Ok��-ҳ��"
4�ڨ�/�n-�,xH�����!�ې�d��*�UJ���	7��kH�������xXgQR�L��s���+�רʶ���:A�v��i�˄� )!�t*M	��Up�;�D���QGx�KrP�ް(����ц�MC5و��b��/���S۹Q8�P�Gx��vq'�w��Baoܩ��� !^0p��,��"AoE��y�mx7�Z��;�6R��B�����"x�RU�P+-�e���\W����ᅍ��Fl�}n�9�Ȏ����B��������a�$����%EV�,���V:�<c�|�!���>Y ��k�lN��Mu�_e���c.����V�P`�t�y*���E|M����2O��N6aI��6�?@�RƺIp=�H�Y���@/z�c�����a�aL���eE�p
7��k�ᶂ�E<�����\M�گ�����ŹΘ_�C��f��%�p�AL��:d;�
���z�E1�N�]��a��6�1�&��X����-�
�Z�0��c��)�U��ѩ���y͞>�����M�L�Sq�5^��"'�]z�W9P�Uʲ�F���DA�#��]ODiA��m,6��Bv�|\-v"�Op����4~n���wf�����ZA���_��J��ɬ�N6����2�0L��бv������`]�P�٨ͭ����,��}�*_T��ԽV&Ҕ��PLZ���)~�tm��G "J��[�jht�X��Z_�U{_�}ZU�b�	5��s�1�T�:@�˔�ν�E8��԰S�0�� �x{zR���������P���nW��F�5͕X��co�!�\��������ud'��
O�KS����'$}\��^�-{}zL�j����`��*!�\�VD��U����P�+=�Ř��/�/�O1��)s�����UM�Y/�1Yyf%8��t�|��b~K_x�	�,�V�+BW�S�
	�A�gu6�\Z������ñ>}W��S�F0�Y"����f�Z@�-zN�4�ˏ�x,FO�z)S�Yz�3ZG*\��{��r!�K�eX�Қ�<��ݹ&��^v �Z���SY<	����s�Ba~S�3�+��%e�.��2��)�1�M� �n��Ѵ�k4E[P�3�Lі索[e�%>���;�"�5~����KJQn�F�X�4{-��e��!���H��DC��	D�;Z���w�B �*�ѨV�J���S�Z�qA3`�t<�r1[��S�S������-�AD1a��.��I����J�Oߛ|F�*�PJ�H�J�<nH ��+�lU(�C<C:��<��x	L��g�!�r<#�*Xh]GzK�oO
�j~D�߷\;;�>C%;�b���L C��L���fo�H[<
�8�?<��!���9�Լ؉��Ǜ6Ț�$�1����j6d[�nU���L#��q���V�f@���;�"'��Tw1�[��6��c�DOG�J�-܈Q�I���<����=��=������B�<�O=�04�'?Jo�A+ee|�=������9�K��P]u"-�y������W�o6��!�N�q�>��!�d��o����7׃s�=� K�'�6�wx��U�D�1#�BG�}�|��^�:��fW��kcW��2L�+����i���;)��f�x�v���������N��T�0I���JT��J�3��8Q�3UF�X@��"(�։�H�RQ����?���Z$C���/]��1VwŢod ��S�m-<B�Y|�͍D�+�Ԁt�Ɇ�Q^4V&Q�!�9��j�d��J�U�Ȁ�2�H�|���[�ڔ�d��A����g�-G5hN�(ٜ��ſ�5�P:>�`T����عc���e�$����C�	w������z>��ӗ���.=Đ�Qy���xy�,��"�e�w����?�h 	���+�V\��u�<�������M�����N��sH�)��b�?RH��q���!�\���1�n�c�ϬKPw�u��,���G/���P����S2�~#V��)�6E`{A��{����(�+J���J�9�	���Ì�������i�-���j���HU���n
uW��#R��(YK u��JF�V���W�_b}w��`l�����:%(6��[�e'�S�w�KZ�9�/D,�'���]GIe���ix�>s�M\�9�j���UN�?  W((�{Y���SV٫e�?�BE7)p�s�(�T�8Z��l����Dś�qp8Q�Bz9�~��!'�-�U�{�rR1�P�V�g`��~���Ċ�B��ûE���WgB�^�$E���lX�)վ.I�O��a(�O�|!"�M��{^qj�+�	�7��U6��n�Ϯ�6��J�'Tp���aB柅 M�FR��T�i��X�˩͈��D�il��O*������xs6+z��� +iR�Et��9��<
ѣ�b��bc}�U�4ں;_�g�y�5C�W0��\�b�<��(���{O�io���Yl?��%`��95QS�J�yl=�?��QO���b��9U�&.)���<g���$��i���%&H^@��~�j��]�eW�"��Ĉ����ٌ�wnHW��!�>��0IM��l���`E� ��	T)F�9t��S¨�^��ZU����"�W��b"����ɂ�2���?<�	~��*��+���d!u�%�*����l���şѩ ���$���m��8H�|�����r�9�Fo�*�w���/�&�m��熊;R��N�ɴ\^[*����qf��:x♘������q�Z��[�,���M�i�DM����8U �"W`����+뼪�Ҕ0����qb�Z-(<8��*�*��Ș-�@�8�Wբ��& r����.�bA�ϳ��'�_m�� He����{�ܼ�_tɗg�� X`\�aͤ,j>�ĭ�Q,�̺�-T���b�l�O�cy�o�x��f����#�4߸	�ѡz���R��?�D�`iG߽Q�rq}rL�0XB3&�h�ẽ��uR��j�p���
W�xa��*�
������M�=��Ka�/��}�c8�6*���7ʗM����q߭�Z+�X���i\�j�r<ٲI���&�̟�#a���}�U�a@�L߲^�D����6��{y�����'�1�t�۟7���~��S��]� /�s�oe���#X���=��ahn�� ���Ҁ!p� �+Q�*U��:��O�H��-�-����Z
����@�C��]����p�F[�R�p�G�&�� z��\���R���ݙ3"8�O#i�5�yw:2d��$'�q�����c6�+�T+}��ή��ij1s�\�,�BYɬ��n��{]�[���cG+��c��g������_��
Tu�!&[�\�)7P�:	lN6�{D8�1�ot�������c�=�A�k��{A%v[��7������T�m5�����c����Z��sm��!(����;��M�?�E�Mճ�z!*-����J�����sm���͉!�f`0�s�X��������<�[kA?`�A%%x�ɡ�ʾ�&�y�c�&�)��8��J篞錨;X�@��im�u5
�Z�|�Z-�_2����gc	��E yp��E'��IupJF���^������~��;<��T�=ɍF�L����N��ǁ���O.��T��B_�½gr�T��Ѹ1��Ԍ�p�4��Y
� r�W��Ʈ�ͻ4*U�]=3g��>'E.t�+�������|z�9㐒��ي{�s�uG'iu���;�7��]:_��;�_Ys�r�10�`"��^�O�&� �(��x���ԝ;�/ٝI�et�^��Z,���{�h
Q��v�4�i���y]���gO6���(r��$�: 5���������~3,%����S; ��&�40��� ��@@uq����%,��?����X�%��$v���f�h �c��ђ5�cƧo��Y��1�	�ߏ�y�Ⱥ�����^��`2��X۱Hj�����{0J�Ԋ����7:o9�-E��[���l�ގ4Q/je_5*"z�~IfDт7�~a��c%�L1���.5�8�L�϶�S�ݶ�RG\���%F�O�[[�`�H��ǳ8�V	�ݎ�^c�&�A|� �Ԍ�v�(y8�NM�|�H���;��sp�	������u�p���%��up~�F(���p�	t�'$��}]��M�wҮF�o-��J #n~1tL|m���9�8�	[��\ �Փ�����j� �r�̳������;�Ae�	:	\<��w7ǂz�L�Wz��o3���B�PI:,c���6/!Fx��3>Q�]bq1`@���wݥ�@����S����ly�U`�F��:ɹe��}���se��i��k�[D�OJ��0(**<��չa��S(�]zÃoo�Q���T���}�;Z+0� "���G�]j����(5��p���8�`�Θ����r)$C�E�>޻�g��pX^�7p�{|�U�!]��P�8w[@y�z�f�
��1	���ӓ�^�|�c!��3�l�i�qkn���������h3m�9���*j������GV��p��Hqx��*�p��U�}r�[[JEFZ��d�R��ii�G���p�",�����D���83N{ͪIĉ)=�2^e��|·�N�uI��d�3����g1hG�w!��6t�qc�a (�<�}��Y�~w��8T����f���A�c~P��gs��xВcF�l?>�+��oF��J�5�$@�F��u��ڎ;��(��Lב0yEp�!Ci]T�6���^�ܡ�ijg>{��G|�~s\E�C�j}�٣,��0���}��p�{Lz�}������N����IƖ�T����"gQnߨig��u���|m���	Q��F�鲇��f�K��bٟin��a�YF�!�{2�t�$�CH�E9s��n"�;2pe9�꽟p�NI�#�u�f>���~��\g����]�5
��=��3v�^�ǫA�0%L��k,�p�o���a(����g�&�2�i��m��j5��R�$P�Xc y��&?����a�XUN�@i}%Z��b�h����m���~�j�vl��G�Y3��lU�,��~��	�k
W/��1^1:A%�r�;������x�wKS�I�����������ۑ��XC�ew�\<<&CaWLY%I�mt�}�ʏgy���L��*��8_�x,�q�!�BOKQ����{x�I�Fʎ���+M8P���cY1�[��%�kM�a�E+ޮ��ry퓪ɥ%����ȢQ�@��W�j����f+�+�~w��Nn�^Kk:ű�î���|����Ҭ*�\[>��_TOG�EԔ�������ǊQ�>��G���e�Ԃ�M=�G.��7�#��%���W�q-�D�0q��[x׫^=���y���Y�8^�o(�^�?I���A�ϐ.�}��2�gS�r�P�,Ġ���><���������hdy,Ȉ�X��W���s8����؏�{Q�����hN �I�f�ݘ��(]�X��y3�[H]�s��h�^��֯\,�6� 7�(����{����K���y�W3�RA#�鏎����8
��;Ϸ 
�]����KҋU0d�7��b��n���#��H���P��!����W��,
*�9�r�q���'ժ�(�B6J��e�/0Oc�̵�e�8o@ڀgF\��d�?+H�ڮ�&����*�s�p�h�g`��L�����Q�|�C�������s�:��iGD���Vq�/�̰��LYU��'��j#���9�(���f�%��	$�"R|gTE��Y�՘ڧ�2C`�]��K��4�-�_>l~����L[x\ �n�v�O5p@�+\K*�+��~-��S�E9<ՈO?�֩�}<O��р	�,y}4�-=�3��G;�Xv�Kr��B�[,�n1Y�_,����%�|�HI�rs�2t>��%9ųr��E:�L�(m[ı�B�((-Xp0��}���*� 6����!���� �dܭ���` rm�0�J��{�8��q/=�K3x����"zVܥR������<�y��,��g�N�24�zz�ԸnJz�ҟ
5��"�g����a�W! ����Yu�A �r�@���\��>|6=��ؙ��KRZ���]��	uϡ�umV�MH�st70�@xl6�͹��SKi�?-I`Pީ���w��t��?�U���v�j�00����jr�b���˷�����p�=cK�O���j%�
8\�]�
�����vD��;G�>5���rzKY�ݤvb�-��]5���Y��ߒ���V�7��*�$N�:Δ�;KwN�q�*�v�wX���M�w��i�9}�dY�v��ed�[���aؑ֫2�<R�}珞g�� ��Qz�D��q�8ҥ=H�"P
�@B�r�z�S�H�����v�<y����� >4Q�g���4��NQG�z�	�TOL5��Z�r.X7���f��8�}[/�~�@���.��}y'�r��!��BF��!��Y_oLP{�x)dgp'�C-��.�{���棾��Nv4����l�&��o�� ��=����X�r�g�ౄG0;���u���毾Į���Z:����ޞ�K��f ��,�W�D7���t�:d>H/q���ZJ�[ٸ/�u�S�:9�⽑fTO��o�Ǔ���娑)>���ړ0c��'Ǐia1L�P�f6��d�={Ŗ���'���[�hS�W+�r��Cv�k׳5��� ���7��(Eߧ1��: J� ]\״����)ߊ�go&�g3�Ѥ��T��U��_ʌI5����o#�1�SaIlj�X%�м�\�]^″+����v ��9�M���t/�)�Q�؆�
wU>�9䧭�q4>&����g��
8,�ҿ[�<�c�����Ĝ����=׈\���F����?"��R+EQ�*g��-N5�
fq�&C�\�C�6٨��67n��Ȓ{�^Mн����������-�!���_�t���l�ӨS�\���ѣ /��rx
y�V1��� �b��?�ly���6�gu��������;S�\j��c���o����Ê�M&��78�Qb�|:���Ќn۔$�PP�4���f�$�g�fY9�'�q�V@��:�v����?�x���� �I+47h�߁�|^��p�SN�y�:������]���F4U�������k��fA]�jȼ)y���jٿ�&b9����:?�[~��Z�^ɴZ@���	UT����HY'Z��S���(D�,-��u�Oުz��B҉bs�wơ�~W�icL<

=lj5�\��h��S�}��>;���/��[7����0�_a��� lP�fu�,�M�\�)�;��\�_�M/uS/��_T��F1\P���hӲ�$��S�1�UWп!�^��`�8�s����oe�)�Y;�qW"�"1�0[」g#���ur�Q��cRv��Sa$Ed.����5��J`=2�]c��o����A��YȨZɤ�zu����/z� �����D%%��&�7���i�ϮȂ9��VF�\�i*������p�`����h(Md��%���񘿂G0�wl���U\��|�3�Xs$��.[�{FiXH��v�ֹC/�=�hX�t�ik����!Yp���1�D:#��X���B���M�>��T#WV|��`i�d��FV٩��b3���V��c�(���5�K�q<�|�PX�+>S04�9ڷ��y��� q�eR�1���Fc:K��k��/{A��ᑞ��p�A?�JWM�z��wy,{M�jT"���9U���`�� �
�rii��ĲT��B��Z�ŉ�!�M���M�U!�R{�+�?�^�>"�~�2��#�(/�}=�_��wqv��
�@�s%�,l�'_���-_�l�� �����f�YVES���K�[�q{Ѷ�et���ǫo?H����c��l�1�u���,$n��:EIK+&����Z�5�̹�q�|�������d28 �-���a���=BX�V)�����?W���Ki��~e�(EU����Ԃݤ���|�3�h�-W=qgn.0��-���2��k���,�p��Ѡk�����sNR�ZG�\�Q]�`L�+cX�D|�.��&?P�D~�ax��w�d�{6� 7�T�9B(�&�]��X�m�7���G�UV��w��P����;�)���*�W>i�"��$(���^��Tli�(�Ks��\�	���Pl���v�=�!�����o�vvg3�[@�>e_tS�dX��ŉ�F_	���2���n&�<+��L��h:
��Ǔ3P��� �V� ��w'�Y��'�(��Î����/�H�Lc,�u�v�Oh|PUz��ZMk�ڻ��ub �������fy���c�/�Ž�4��]�0'�Re���f��*�s�0�i��fO��,�#�c�8�]'�G�}-d�x���6d/�����}%
���!�3��O�L���$$��O�h�tB��{AL�S�w�,�.�	�P�^�Y^Q�"�M��+��j�G��1��p1����rX�Pk&��W����C�����^3��l����;�
�]��Ҽ�����g����H���Q���z���=-�ă�X�o����ZIX�ƆW�n���(���@��{��{�V�������r\�t��*�"�>(��U�Y�/��^6�Ӛ�}{=�b�(�k�=�)h��[E#'�	����pҥ���fc���6Sò� ]n��(��莊��l�:<j��+x�__��S�%O� [@y)�� ��=��Tv��!*ā��W�DW哓���7'�c��)͕�!L���������ig3�fL���� �9��:s֬�y�ԕݓ�F�P�ʺ�=Kc1S؇�ѷ��a']�C�vp�wO�U�����/�w� ���Y��@F/
�`�c,��א|A�?��G�:���	T�������b�"��j������3��d�z�r�ym?�u��]& '��	Cd��(o�[�LåN:����,��&��0���jQW�Ɂ2�2i���]2��
ǣ�:kJ�cT
T��$�0t�ҋ���{��� ���\F�Vi�j`�c��,�DL7����gҜ[��p�IN����N�W/9Z}T��ً� 4A�
��칓�H�'���V �9r&`d�m���O�����Q"�tǯ�0���Y"R��>Wo2>�c��57U�P�f�Ii�Hk\ݯotloX��ʫ<������\�\O$, R|=��r�	|��R�*+��k�ԇ�櫓!�@����b�5�u`�Kb��x��?Q�����a�+��F]�XYΉ!W�TC�[�Rq��"�Xmq��
���p��t�Π�����gɈ�Emڶxw�[8� %��ƛ�oj�Pd���{�3�F���[��B����߅?E܇�J��P����̠��sͩaoh�ϛ:������U��;���ܩӫb��CZ���R��0d6`��ބ��u��u[�8��%A�LT����H���3�3Q�e�����I�k��xj��3^=p���@�G�o7��X������T�m����/�c��i�[m�9Fs~��clS^�.a#���U��@ð(��R��g�vvJ��`�/����:��e"���!ȤvS����Q�`�>��r�����=�p'F���9��gc���X5�,�0�t�����H"jq��Хo�6ל�ݮ���"�$��,�i8�=4��bQ$T����k��̣w���,�@<-N�y�5aߌo�?\d.��$�!��ķ5��	U���Rz5|��!#��&�9��=70ﱹ�>�w@ۤpcg���Z��Y�w�^]�^G{��_ ��Rm��x�����<�yoWG���@Ði�	v�|�V)���o� f��tU�.�6�s?�y���*�}=������,�sL�\�b�I�ӹ,���N�b�L���w���*iY�� Hfjז�z:Tz	#�27ƾm��'W�~�\����D�mg���ѫH�(���A�R�͆�:nU��mfM�@A C)�\�+Z�J��3=��z���kv�j���џLLat�3q�)IJ��[P��:��N,0�k월�;�"� r���f��j.x��qo%��"�Iv�l��� �t�H�ty�4�^�TZ$])1��
���~lg�@�18��
�~����C�/��#���M�!-��E
pm���G7pW�0u��SVwr���3����1�f��2c��G�����[{]�+���G�Q!V��.Z\y�ik
xX�
��H�i���n`���+���I�Q�V\=�K����	�N�T~�z��ɒ�?�d��W���`�y�0���l�V����xe$,�[�b�,,�;�8
;(�)��p��o��Xߨl��:�L�$��A7R� 9���U��O;����M77Dlǟ��f��z���9��E���g���4C8�j��e��m)$��� �9�m�|{C:�d�,s���L���7=�w*��v:��W��@[5>�=��C��ز��:w}�2"���{�{D��I1�x��2xat�4��l�a��
uش`��C�>C(��:X�^�>@�Sj�����M	 ���T�|#��L����@sh D>.Eg�)��m�I�Ó*�cGK���P��vGM�z5��Kb��3�ȵ����+�oh����ҋ���6���:�@z/Q[ڠ]~������~��\;���[T����W�Q �h�n1���
�]�(cZ�zQ�B
�krz{�D>�y�^>)�j	��Ҡ���H��bL���OF�#5F(�_�-.�����$�O.�S8���ARcj �a3���'@����lGch�[�
�<�1w]B�^z'��ͩx�
�� �w�%/�o������t����|#PGS����"�0=�bu�թ�y�"��E�"�:V�����e`���t�$%�#���"�|�(%�D/��ۥ��7�t#1g0�:ր�7K��4����񘬽B���jP�E�G�l��k�(�	�a�b%�\�:��c��8a��m��n}�E�6�|o��"��]�z��@,���:�ږB�^@��",�DdY�lx��Az�:[����V0}���(�(M���G�f&�#&������	��CM"��/���!,�M���-��.��*.�z�9�<�(�1~8ݏ�x{�=��q��7�~�˻�>w1��,B�s�A@c�G=�2�׻�p�(A��21W���#�O�Jkjx������X�����銳#��3pyG�l�kV��̌��˵7s���vԼ�i���!���H��g��(�+<!7hH��QAю �^`��f�"]��GQ@9-�m�WEi&c=vg�K{��B8.o<�N��
$�B�&�v� �W$���RfW�M����`��%�����m6ޠ��!o@Ȫgc���_���2l~|z���ԅjjc�Ɩ��)p]����H/�C��񐮦��a8_Z͜�b��f��4�B@��~����Ȭ�H��������Vy��`���9T�]G(�]�.]_���{h�@OH;v$��l�d�]�T�FS�%����{JS;} �O>�B�����d��-�L�ϛe�ᔂ�l��;x�+&�]hQ]������6���f ;��T7���s2�7=F��@�o��K$;�<sYM�;
���p5u'Yܦf%�!�g��SH&�ېE1�� ���F�7U'�e��J��~��z�gA�_���v�'��ϭA�)ɘq�<W�g���4��&�m9���m���&>?�L�`&��ߌ ~�I'���ʟ>#</0�4$�S�zS	���G$Ҟ�&P�*HqVuC�o��BNƼ�Ih.�(�N�Z�,���P(i_8Z�l���|[�X������lx�!QY^��T�B���%�$?vei�� z¿�977���:;]�E��~�F��w.Fѱ]9��A�%U/�-�K.��P"D����c�s�v�V��n��O��/�,ٯ�T%_V��ĴL�Ɠ	���	���z�|ڶ;"�Z��V��Ж^ �v=�����nF��y���'-G���f�=c���< ;��Ȼ���Y��0�<_W� epe�V6�!��"�*@�cxrr@��&��]noăQop�9�FE5���IQz�ŭr��K|��٨�A2�RK>��y���MmCL�Z�=��n�B���\�k����z����c���|�`i7�P��g�t��j#%��m��6��Ñ�7�a>��ʃˮڷ��š�b(�Ww�֧��6�-�`I���w�B�^3�E1,XoE��L��`+��73�D��P�����p3M,S�A7,����c	~a �.�i��9/ӡx�yv��Yȫ������mN��.�T���zk���nB��UK��[�����
�4����4d:��w�� �%}�B�D�~JM$�h��#��b�G���L��_��C'Ć9��l�Xs�j.1��{2������۲H�D���e���>Ca@�CM�z��ןF��ɔ$�ؐW���G�dG�����q T1l�ωe���Э�dK��joz_�Ǟyx-�sn�l/J�Z-�<+��*�������uM�,Zy6�����_��$�VG8���	� �/�;����L����Iz>,�g�Qe3��ag&������j��p�4��F^�s�͏z�G]�CM:�f�O���ǯ�oUH�ԉ��v�9YM<�.;��1'��>Z��~y��~C�e����}f�ym��\�5x�����R;����ޕ~�S��x@�>l��1�7�~**}�*��'��n��r&�f�L+D��ij�j�Wc��]3y[�"�ԯ�����й{h�	�+е?Q�36��9��[�Z�s�(���	�����Q�5�&�>ʸ?_fԠ.����x؆ ��"j�w!��[�?^�BW�){b�� �̢AQ�'R����E�&�Q ��O��=�S�����O��ʫ��0=/��w�om�)�ͼS�ZH���H�Y�d�`�X��e⦶����!�����g�WI�g��$e�{����:Ek�c!Q�W%�A/Sf�H�QJ�9�r�|8㧿7$//�gn�P��oRg_:�ׇ禯���@�����L��*J���"(#�}�R�����(��a��p���j�͘J�i"��YMώ�+@"B~筇xR�Y8k�a��hS��h�c����N��O �l�7x��R��������Bir���鴉�q�ȚS�
�(v �V�}9wK��:�������3�w�hqF�9��{/Q���C�����ݍ���P5�S����ܶM�6�qV���'X�3��܅ӗ[�=�ǻg��7=#_��e(|d�����Z�ԠN����QG&��'L�mP���qHg�X��5�AY�7��y�_v�IU��AtȔ$��|�����R�����*��Y�J9��:J�=#����l ����(��n˖���o{�C��z�t�8
C]k��H��	?�m(�a�%Ϊo[!�Ye4s�=��-F�+��ݧ�*xǲ�9��iX_H�r8��m�ωx���.��k��G�&�t���6�_og{��6-��+ݘ� \hciX����qݻ��V�r;�9c�B	-
��}�f�,��=��
��nϤ���rr��eHH��V��Ҧ�k%�07c�F:|D�V�,���7G�^��\����/qMe���|#�=�x~Eߜk+ݝq�3O��J���7-�Z�%'�}��}�H��PJh�����J��k�O�̠�?����~&Q,,� �lOo�kPX��Z���W���>!3uMͩU� ���Q��S�_�s�g�M=�O8g��rP-3[~��k����z�̵Y
/�*��
�$r��/l�E�ӊ̳���Wj�l�4#�q5i���Q�=b��?ɴ�Ϣ�s��>Ilґ�}}�Eu��X�#��t}���vԦ5c�._V��
(|x��!+��$���p�&�ݶj����]{�0g��-��TSʟu��OI����kL{��v�#��7��p��q��f�k����H�(ϵ�a����C���Y�HT���5���T}8�>��+hV�D[�WkZU��T����AD��~R�+�@IED|bn��G`)�R���5�M��4ed]I��>�����Q�9�*j@EhZ�l�^&���`�:
��S�>!��HF�;NʁΜ�"?���5�a�G����h�x����H���qI>8t�����6�Ksd�iù��/y��hs`�Ele�	Rm�}�[���H��n���*�@Z��.��}�c`m��[��y!�ZR��I8(I�pk�~�b&�<r�|hy�&�w1L����S3�2��7l�N ��lU� ��Nq�8��'�o�껉� `W��f�FQZ  3��_ �`I	���9�;�
��y6��r�Vԗ�׻C~����"�w��	`��%%y#�Ϲ��Q��{N���)d��"d3�
 ���B;���eR���_�rs.uS�$�����Ro���(玬��9�����ĝ���aR�S�h�����gmW��V0,%q*!�r	3f�(�$��IUvZr�=�w��~3��q��H����LQ��3a�Z��/i����T�ǹ�Dk����~��N�R"�Ь����4���K�EK�L���zP����څi"i�"�4$ǘ�T���d4���W�Uz���H��)?�?�^J���K�P�p0t�q�^�B����$^]��~��5�	�bF�S���V˹��Y[ ��V(�[\O\&W��?��_�E!o,���a6Hf�����%c���G�X�W�8#�q�6($O�Q�/C��[ý��Q�9z��w`��N����_�L�,��� ����H9�Yݗk`�|�˾�@L������p��	���_�P���HPf9Պ��,���z�8Q���@
�b:de�o��%7��e������
�S�"?�F����@�ˆ���g����:j+���l%H-�ܠy
z�D,�G����U��O$<Ki�L� �i�+���M��{蓻�=O�l���}�n��vmƒ�>#��G�z�p�����)�����x4�d�����nI6�!z�\�0HA*H��/ܥ�'IX�WJx�}L)�l�������@Ր2����{�6�&֏ᠴ��WEГ���^��&s�IY���W�/ a�\�Y?����E�M����浪٥�8L������=��l�����H�I~�W�������R���pB��V�1p�l��n����j��gϔ
�!C��I��}� �.Xx�'����[R�]��f�1�	Si��H��p�oǴ���u�ԥ��&�
���`�tdf�^P�Y�!<���o"�n��}��NN���{�po���)�0(������z]?i��':�Pw�Ā��:�,�(�p��c̃��[�vщ��ڳ�̞�3��Z:�ٝc렳̯D;������,������.C���6�H�,��v��T��j�Ben6�EӒv���9V�{)�|���}	��3 Z�8�H���r3":e�oJ���A�Z5V��N�j�^>G-}&`�Y�_m��t�,��61!w���}�1=�+� ����mX�~�����g5_��>j�K���p{D������ʆ�R�'��
H�ř��ay�璣��5O÷|:�H���J1#��"�雜�U��`'�� K� ����<���?/��>�@�WT*��Ĭ��j������3pӳT>*���X��5�V�#n���9Ω��JF���W�JxB�YUA1O���O��q��I���7@LI
�>h�<W�_j�s)��gm�Y;=`cqW���,
D8������A������O�<s%��b��t�*(*d*Q[�,t:���{��u�ު�ʜ�\���9�?��v�?�|��@ш�|�k�j�U�~����x�+�S�?#�\׻�T����
nؚ�ߖت�C�Bڼ#\61��c����6��&K���e��F�260�5-g�^P���M\������A��6g�Չ-�8�d*M*��	s��@H�}��D��:����&4��~%�N�����SЃWC�)�G�*�S���:n*�{��̉_�[��R��%�=K�t�:ێ�7�1(}CT^ާ����c�~���כtQ}���f����UԘ�.+�ܧӑ*he����dFH�Nm@BI��C޶�@Q���f�ca��(�Mġ�>P@5u[����9�b�=-h�x�[��i��P�3�7�i6�S��r��2a#�6])CI52҆)���SmJ��88nU�x6�*n�tuP�6����|k�e%'k�k�J�(b�gF�hƃܹgz��rncD���_�Ük�:ȝ˵ dji(��!�`P踥�}���<��eڳ��~�|�{�+0��� =�����ق��>�sz�=�3+=
,rJ~Oo�R����k�v�z�������?s�K�Y�������U�j�b ��]o��y��E��]
9F�}$t"5�@���C���d�f���ֽ,���wnݱ��,{h�yU�7;�R�1��i�syN��>O�q0�� e�\S�k#���}��/�r�����S���ݫp�oJ�c�ܹ�M�F\i��ٱ��d#��&�n�tT�qʨ��U�7�C�ջ3f��O�vfRۄ%���ji�z|��_6�טּ�k '.!��٬�& RF0�4��R��*�l�DN���2�ٜ5}|�>���Zz��T�4Ĩ0��s��\�����t��ƀޞ�>\��	ҫݧHz�$�_9[��[� ���Xp��֐��4$%����'(����w=��͇=��Z%�=u|J
N,H�{����r�K,��I]�<������#�#n�3��V-������`n����9y�g:f�S�d���Jm�v��K�υ\��Am]�0�%�fy���S"4�8}u���=8	�r����Ad=O�����	-���݊��)��uo�q�}�?fLב83�n��I�q�����v�~#y�i]:��(�^Ij�TLy�+{�D��?������.����?��%��E�y)�>���2�D���괣�z'��?�����N-x�n�R��N�+��ѱ���Bћ�6�0
܈@��m`H��}
f��Zy��]~�1��,���34?�0�e΀bS�ּ/S�il��.����֌P狙�N���^Ku.8�V��n^�J�=m�����%�6�V,��u7_�@Lb���炘{1e` o��F䶌ȱ"5��ݚ��l���C�` .,�&�F���?B�ΏՈ����uۚKoi>i�+��e���@�R{~0���6�⩚|�u+�R֤�Z�>w�Ung���G%6ho5Tl�|ט��֦B��Ϡw��{��"�`�\����4�����[Bmv�Od�Jú�A����H<2�9��E��*c(���/G��'H$~��!{w�����]�r��m��E��_��j��#X��}2AK魄�)��2�E-�O��/G3	�Ǫ� ��cv,c�ܕ�P�֭�� ���՜�u���G��*�S�!�y�ƒS�X���\����NiO�(=A�；��:w������˟O�-L��{��3Y`����}��1Z�]%�c�]���� ?'�|�9�3Y$pg�`7f���nr�--ua���@V_��}8&��{�7��������}fh&�iR��ɇ���<���/�}�z2r�����_;p69�u��������������8I�s����:�,n��R��MX�au��ŅN�`Q��g�m����8��a�ݼɈ�0�`)z������ט�,vj[fF�����

��������>C��v/��/���0��<�3�hsY�ܝ�8���|ՠ��<����/�HNO�88�`a�{nX7�^2f������O���*Ψ�e�JR�>����ȵ������5�9}Vj���:3��ؓ����@4�'K�f�m�ɘrc��H��m�I�g�Bk�m��^��al�(��y�2(�C	/��5�E��r>��Z�L�U0�7 ���KtUG<p������ �K�>'���U�췖"
�×+FxV0"��.�W�"3�2^᝗Y����x�*Ղ:��]�������ɔnDwH�\�"W�r��Y3+V���Ycs�ƅKOE��Eĉـ����t��߯��v��'L�\p��g'2εO��$&��m`�w�=����+J�"lX#]���0T��o1 |䎸�H�}�Ț�ݟ�;��w.���@;%���=`Q�^a����x���B���)2��`�S����H2��E$��0�@����N1�!������D�5d�j�w��;ς���^aDX꩒�a�����t�,-��TtNOU����(�3T�#�l���^7X��jaұ����$�"���/��ѥ��2#��m?Q3F�8��c�Jz�^�;����!��ѻ(p�#�"��+�bg:���
��9�TR��;�؎� �I���K�1�b��^{h,&ߠ��D�'�	����~������!}a��G�*A~�o��mn�f?"9������jη�FF�[k�<�o��\�E;�@�Õ��x�U=NÌCK0���&W(w{����Y�z�(.!�x�"��D��t;�4��3�UbJF��/� n�B?��<Q�,K���E7��Q�#�^u�'�׈t3ةg�G��QOq>�tj؍|���8W�0k.����Z|��"��&5�/�x���ۀʎ ���M��o^���~�P�41�qhj>z��ҍ�̵������hY&.!�dĺ�&
c䓊wޚA��'FOV=-w�
vP=Ld��� Z���5*�R�B�B�/x��ߦ?�n������E0?�w��	�T'�'ރ��D��p�X�� %�J`M�[���?�
g�S�&��� MWe��z�>��a_:\j�/FEw[&���|�
>���A�����Y���e�C�!��l�bH��B-6�o�݁f�����p�j�)�����ë���0�i��h@�~)'G��s5��t��e��v�>_.m������ǹ�LUi��M���yʦ/l�8���8���0�v�x��{dn{5�q�n|�;������� ��Śt/�CY�5���c?�E��2��uKξ����bB��¶����ar8����./��Lk\��8i���m�V�!��%����q����$�#އh�.�eG�����_H\_��TX�Ƥ���l�W�&����
��/�7R�V�"p������'�Aà�ߵA4Woq��+��>fl����h��Sy��HJ�iR�Q�\r
�g��S@��Hƾz�xR�ɞ�M��?�����P���j�ٟ��Y�T��Y5"r�#`�=��J�ss}���	����'�����\�;�hhh��C�n��l����[�n.�~Ͷ�)��aoȚs*3� �����;h@R�=�O2�=o�ʫ)���x=4WC�0���5-_�����w��.���{஗�T����U��I�>���6�ޣؓ*��4��9r���a�����c�^��Z���G ��T4��7s�0:�����_��*�ӃIv�@�8�d�a�>�b�W)�Z	ǈ"�Lz�d�J-=Y���g~z���H�im���Y�ڥ�����u/>�x��G������.$W��`IC��(���GVxP��S.1Љao͆>d����7r|͈����.��	�ס�86�ɥ����YU��aG2c{�2�Rw����8�EQ�;���Y'��P��H��-4�,�^�e��3=j7�3VDwe�>p��T�8I���7�Mu�p�<�3�'�V����:�3�,���l�\ڊ6lN�I��0�龼�V����տW:	���cM��䘴�T֩_ќ��d�ps�QS�
(�W}�5��!��A���9U���?ύ�k�]���aاWS��s�>}V���hE�e)��s}����+�}$4�DP����6H�H�_��X�/s��;sО�d�*��.8��(>j�=?�Km� j�c�Gάh,��%;�Хt��  -���aeO�h�Q�_�%�>ϲ�_!M7ͯyp#X�b\�KH5�NE�y��q�v1D��GL:~H���r۟ݵ�)��2&	ݒ*��׾I�9�.�ocԠL�AhF��*���>��Zk-�߭��X��֡�������G߽�F���mOd5C�	�E�V:�9�4�\]b����Hb"' ����ȪǤ�h�u���:�i���±���Cn��m �HUX�:)�Y0g��KqQ�]�%�O����j�Jqԯ��gHJN����p(b����H�p��J5�1�2 ~�P��c���^�YT?�f��M�F���ΰ���0i�a�� �tw?�V��� ���#���ɍf厁��zi��Ҍ �]_�B���^ۣ��,��^�tܐ��_�=o����R���ߐ��m�Ƌb���n�"|���-�s�{T���5���@�b� �?Sbe�~e>	U�.�:��I���	-U]
��N��O�O��i4�?v��u=���&���H�Uܘ)VTd�1cQˉ�c5��~���E�(����&!�wE�@ISVB��*S��`&J�����i&���yR1R�#�ǹ�}�D'�Tv���!����`���+w�]�J��1%}8��Ń���Q�:�+���k�}���]o��dU��� �$<�SwFh��S/����=��v�:�W��h2���y#���\:j���#�k�d�2�]^ݪ;�t��c\l�D1/d*�.TZ�M�; m��r���){�"�����t�n�E�WƢ�����ao���.UX�mbT��{es �
��(���}p�Hll���+�)A��l��<:���Sj�}�.U�b��10cJ޷	���r�;r�������~<ERת�����pʻB5�E�ĆXPE[�oo9%��c�����U�f<�튉s�=��2捻�9�6H�R*?�ͧo`������⎯Mn�j�e}\��yo�k�e�j��C���Bk&��LQ�`i���w;�q��ʅ���s��r�*�y��Ys�:���򏮅LoGD�����-�
��/!���7)���8�\��9��^� � �Ȧ�]o�+�}c��BY��V��(��&����1<�?�U?l�L�Hq{���������rB^��l��Y����\��m��*��$�W*s�)1�>��I�vR�$�L��\�Rp���r�X�*� �b�����T�E]�:-&���k�����u
�~��zc��BKX��zF&�ӟG���6˴�9cO�o�ɓ��W���"R��Y5i�_��=��j�wE���J�:=��;˼u-��T!�.�����<�&�
���f�2Rw%i�y���T|�K�Ru�;��B��sD�(>y8�4�}X��c��4���3Vn��K͙U�� y#���J��5D���	7�8��������E��/��R���
e��>�r�a��}�2'̈́`u�����L�bn9.vf��r|���*�d��[ �Zh����ʦ=�\�K��,׾��ը����x�<?�y��TJ�ӄ�v��<��w#T�!3��V��DN=�Y��>�pG�5�jxrf�@ug�T�s+�(��!iL#V�pjn��g"�xц�Z��:{�qL�~+��t�*��r	�-��<����q�_���([m��"mzi�q	Ф�`Ȳ4-��
��,̹�Ƌ��3|�~Oӂ=�(�%TA�f;F|��R3�7$T��F5c���1��8�k�m�Q�TT�y��L��b,�=��2Z)��h����c�J7<���-h��6�g!�2�z�l�C[x��S�X`��b5TŃ��2�6E��~@��PzG_ڋ3_��S/
i+�f"Ds�����/2R�4Ѓ�p��h؞Nq�S����Q��2��9m�����tY_B�ۮ40�l����ܶr.F�lM��ٻ�Z[%:��R�s��kԥ���ɽ�%�$�H-~�
��5Q�����ƷVxM���e�ne��&۹��Ԙ�$A��h7�CǝɆ�/={�r��J�L&�gaͯ�&�T� L!cѭhs_�������'Je~��
vi^�J\�Z��y���lG�bG���n�:���n���j�ax���UuU�8]v���
���3
����k�t��^�u�0�P�PqV��l�f�ծC�-~��t��}˕��E��\������p��0~�(�â�H}��^�>���l?���V��i�$Х��\����?��R�6ۖ�K�TDо���Aq�>��l��*�|��24����~��V!����s��� C�muC�Ro��}�.�d@�b��I�0��.�
'�&ƛ������mg������_�o�M?��'e����Z �U�R�Y�@��p�_qu v�U`sbB��u��H�҃������� DE��-�e@<�Nzv�k�c�L5�n��O�z�ZEW�����X�)�
Q媬����g�4W�@�v��Rd ��@�9Cr^3���W�);���f蔊"�b�F����1�4*�[U�U�ԡ�]*@��Ayf��nJ�2̍
x��*�z�@^��kRc���+�5ȿ\h�Д�G�𠲟Rꠓ��8�ī��R|��ȇ y�CO�0�� �w�xμL����>_N���M�UEٚ��X�E�����X���n$�`��
CA���Nv&*��3]�+~�7@-�����BbƑ��P �?��<�W�E�s�]E+�����j�k���J����O뀴���XG��V4{6���Í��T���v!�Ge������_��Q�i�粂Y��1\߻��F��O�l��d+O�[\e+jSzr�:c�^LLp_���T�o�RV�B�����S�̩�I�&����ƹڜ-��x����{�����'܅�_�S�imw�]x��*/
}���1V���'O�$Y��n��hB B�ލ���xbgG�����Y��Z,܁�1���tnA�?�҅5Q��W�]O|�Ư��4�H����+]����Q�R=��9%��4��㸬{��-IxŜ0|�v"0O��Z*�_I��
otm���5
ZPt9N(,�̚`�պ�J���*<���s8���ۿX(F�y�@S8?��#b.����a�TM�����_<Gg[�]����w@��d�Z%��+ܝgG�ݘ��f���jr:S��4��w@���r��b19E�Z����d����+;����M�����;�kY=і+�T'���'�>#>��?z��L�*� Q���T�^�r �^�w!�%7K����m�\s6�*��܉��X����0�ݙ'��X������"��� �6YJu����E�?*C�D�R#�������BJ�%Aw� c1�g ���F�'����zy&�o�O#^
N���rt֦~̈=|a���/ ��$�l�hޥ��	�(�5=���&sk_&�T�>���u��m�T�����݌�/���wHA1���9ٍ ��w
�ӯ4F]�b�m?ŷO�i�E��jFҵ�Kt"��v��k��C)+]���py�t�� �>u����U�6����]h�2 �JV�x�� r8rv(nΈD�����n���R[�t�y�_�����I���}�ž J�4p"�����1�f�}��9K_j�ϡ6�B�
_aY!4�lG����W)�VV���/�IT��gM'#ݦw�����1�
�3]�&��Gg�+Q�U�]�uh�D`�ۍ�㟝LڞL��Jm�ؒ㝙2��>��Ҧ�֗,���<�fg��m�S\s%�2�?i}t��E�#��Dűg�搅J�PQܪ�"d̦f5�U��� ��Є�ڗj���{Y[��J�oXG��/�RJ���7�an&2���"&w�������F�F�Aa���wDwq�nNV����G�f� Qvv+��,F���}�g��ن��8q�z\�G+N��[�/\ߎ/cLZ�`��q��%$�s{�r��b6���I��'�9�mF�a������_G���!�d7(5V�Ʊ�=�ߣ��7�@���6z�ͺ?J�ZL���9��QD�@���E3ɵ�dޯ�V��S�՘Fu�(�:K��2p�ʟf	 �6���Y��ǎ4F�:�"I'7�ܔjr&L�K�%M�^�VӃ`��]�?�Vޞ�x�"�f���w]��b�)�d���ҝ����\�V�
{1��x�_����!)�k��oe�}�1�X�L%��m1)��j���[#��y5�e���	������Q9�`/Ou��8UH�Y`Em*�Ev��X��!QE~��;no�'ѣ�!���X�&�Qwk�8�.'����wzc���X���b{���B`{aX�X38��4sf��q����p��~k�-�;�Y�?n�)��f�` ��<�&��T����z��b�'������2�S}9�	������>���;�'|�]�����k���n'�d<�pe�-�SkO5^[2���O�	K���k&�Jѫ��l�Z�����x#_�kmwB)#�\�~���~�e��,
�l�hyVe�(M���Xb��F�~�J���"��W?M�,>��6������P���7��l/8��9���"2�2(��-�ӈ�w��5��]�m�o�ى	�o�\��0��P/
�a� FiZ���	��[�Uw������?U��KW'�9;�"���l�3+�W[�co@� ���FrW��Y!����^�������Zb,�_J�AZ�8�F׃5t�D��������4�T��?x�׬�r�!���Cis�&�q�󨭮A��G�������ꏸFx\DN�L)oi%��E�j^�Az6�v�J����Gu��ps����0�O0 ��wH�}[�P(�#��=I5R�"\��W9�u㥏A��gc��v
�?[�Y����ƚ�.ȓ�i��x�Sj�z���M��m !2'�^�1�����]�h{�F+�>�Q����� X��@cv�8�8UC&�AW��쉆�[
l��jt�4z���s��~]T���x2���~�/������"�A�&����#����ז�[�PR*�q�j�U�c�.RB�*Mw��O�<�[�{�҂.��(�]�v|kՖ����@)л��_���a�@r��h$TE�1�A��IA�)��K���6, ִ;���V%���u�^�E�#�ˬ"m�m@���O�3��V�%�a��GR�g�f|��$�&���l�&�s�4��-�!S亸�O~��.�3���0��5�2��:�q��F�?��(M�>ӱ�J���o���,�Ss�h%�<q9�ػ�%�M�w�'|�ŞH{�ڗr�zr��ʌ~�!��h�c�5�%���2�5�Z��b�1X&��i_g��XS L<�m���8-�4V���E�v�'.:W����.��� _��s�@#|cW������QJ �r�z�$��hp����]�����BD];�{�V�������z��!�;�e%�>�f:#1�_��Z��H�pSV�jP���_��J1�S:��<u���[ٳƏl�M�f�u���+EeFx�qY��]]R�^1�dRX�]ķT�p��8?3��A���G�޲�O4i���ѕ�"�."�ԙ6s� e��y�����w:�2�!�=iiښ�\Vp�_��ʰ.�pO���
������T��A
_��.�2Fު�&���	G_,�Z̓����)����S�.:^e�`!Pzm��Tlb��������p$Oe'$�*
�:��)ɷ����I��t%��ޞ:$�u�f�K�^�AvM�T�o2~�U'* ѤN|%�|��ܖ�9_�BS�t��ָ{	���8��ߟ����+�������*��PQ�D���S���76���Q����l�Ke+�r?�9���-��pN<��_�������
 ��Q�Xte��H�@����@:Y.�8�u��	�0��;n<� cC��r|1i8_�Ҧh�ׂ��t�Of���~$)z"��3K����u���yz�.�6����%�#Xù�_� Z��kq5M��~o; ���`=�vsJ�JP=5s]���(��V8���m�9 �BZ�6ץ���0��q�a{��Ƃ��r��, C���R�y��<]_���"�����_�����TvvPB�
�x2��TB�e3r���h�ey�7�/:�i����Q!D�����J;\z�6�+1�MdAHs���M���08��h	���\�7����x�Sm铘�l��a���p�:��u�X���SU���9�������%�4�>rAu𣦱�|��N涨�^L]���6���Y��r�۳s�C�����M��G/����,?{ˢ#1�kL�pjW'`�_:�x67�+c���ѝ�ж���9�`w�����6NB�	>�$~ʐ!:�z�J�_�jɂ�l�t��x������kd�N�TJ�_�TRE�.����v=˖��8�Ļ΀�����n�Ç@�/|NK	r�/�R}��6g�7���Jl�F���!�1��e~�5\;�"�9m�񪏥4W�i;=L*��C|��h�&	d:S,,eNvbN�������"M�y����a�����j��r� ��!�Ϛ�888#�ыl_�&�?�u��~,�-���Vq�Q2���?(��}�6�Y�}|���\�ft���r���}��^��c����_' WF��,q)\(�Nq�e�5���bH�����q��,u�[��iRc�#�?k涣�:�g�|e��P��� �&2� [���Yd�m��y�atb󲲭��-[��×�do	{��_��Ȑ�_�(�;$4��	DϏ��3��H��'D�!^&/`��`���ZvQ�����h:F���'VH
]0T���U��Jh�6�@bvm"tM����8$�h!��Դ�[����Ǎm��RX9��
� +?�-���܄�(�Ⱦŕ���\������jDH��� zL�|1�*����yc#�� ��x�rp�7n�&jy��R��x�}�ΎV2�	WΆ�u-��iaM�J [;�[@�3��(I΢���$~W��^5B%I�S���<�]�U6�%�>dW�o˾1��qj��Z"4�Ϟ?�NI�gA��~���&�Q��*�ze��`qǦ���Ѿ���Rw��\z�UyY�fnv�:�e	gޚ�V�lH��f^H��5Z�w+x�P'�A�:��fu����#����'�ap��+�B0�Z���'z
'�(bس��a�uo��J��� �3�wQ�A�WV9n� Bl���ML��"w�dm������v��%�7��a��v�;q-{�o:�m��/����[�>[��z%���
����9{�4�Y�ͰO��ٗ�#�d���z�ܛ�p�
��p$�I�_ve�uny�|o7!����;_��=�V�n't`�LO����>���}��I|)~�Ԫ]ֆbM����)Eg�4�3����2��٤��4�1)Z�Ɍ��_U�Bd���x;7�H�C�O�F�-�ʆ֎��<�u�ڟ� W�yS�~��V̢�t�i�}����l��USMS
�����?���'9�VC8�Q�>��h^!�=�<�5d6P�Z0X��7 >e�9AK��[�{�� \�p���B�����&�f�VX3��w�|��� �?ۊ�2����X�x��/�Q"=�K�)w�*Y[1��>\��ID����ТL�����˛7�߼��Y�&.�g��w33#FLcCW����jfE���i��ã���
�&��PQ}�ʄL��<(@?������F¤?h�<�@��k���Y1��JWP��1�r}\�� N�L�@->#�B�ݳ��T���_ 1�{���PQc��e�8����ڤ|����!�����R!*\�N,�	Tfٰ���-�Wܒ�{���>��M�'t� �&�b�e����ŏ�V�fm�����G��߷ �t=C-�j��؉�|1��a݅�vN��]��[���8|��A���`҃��@ӄ���w�g�a�d`�E	Ƨ�Dt<}��F��ѱ��ʯ�r�S`�>�W+�2ôׄY�-:�oF<�w�X�w����s��Fuv�]��h��>v�(#<�����"0k̐9��V�@��}ѻ�v����he8���<?��C����ނ�8�������gz���m�k�ڑ�;�y�-�	�����Rf����ay�c'نq.2����@�_p'�#�t��^��kn�;+�G�	����lYڑ>bș�K���s�x�� �*4�Ք���� }ϕ�ЁZe�1w`�P�uf�w�d!%Ilz�����`���� 6�뷏|��-}*��T�{���Kp�:��ޏ�*�O�Hd'��_�GU�q���Ĉ����M�b���/�[^"}O��dz���*)0|W��Y(���o	���R�P�M��1��</[���]c��z8��ک�qF�S�|\ޮ���-~���I���ѷ��@)%1h�H���8���cȝ}v�c�6�nd�/�$܏$K�?� �;�E��U�3��Fv�GH}g��l���Q֏ͧ������ƕR�-�$�/s�P�fk�m.ε���F�7���M$tg.&�T�O�����@�G���6���U�8q�r>�g��pļ��.j|��$�d�����ɛ�0��r#���m�k�Z�Cp��z��MX��oV)T�r�ս�}�Ǭ�b���2����0����{�����hw�͑Fu��Gה��eX�F�;UmN�U�%��0�����^ K�>R>��%V�,�U�O��$kx1T+�=�s�U��<�n]M>8l�t�)���0'hۂi�ԓ�����	[Ӂ>��e	�@��$$"��I� :�)|�&7��M<�U*����($Y���.}�[+nA��8��L؉Ԕ�3?J��4�U;����5aߴ�0'����I�,�q_X�����;��
/U�����n�� FW)�tۣ��Us�+�x�p� �d������`��2A˝`J�P�]-��*6�����A_�gD]f����9K�\:UܳkԻ��F��E��q�����KD\(*Ĺ�����P��,*�=e���k�ټ����]��|�h�YU{�C�<�l<O�=�b2�⅟*!.<��	�?��&�k1�,r�M8���ў���������7_8�@�\5y���̎W_gy����iٮ�K��~�Gi��)/B�o��i��K��8L� �w̼�����\�5�� *��(�Jhܙ��s��x@z>� �<,��]D��=�3kK*�dy��/�2k��Xf��|CKX��\�3��Y������:��ݮR�ӌ'͉�r�:*T�~�5YK��O�@v��a��N��G7C�>��J07�Ƀa|&� �u��<�
�$��!���t>S�\��%���/�I�o91Y:RF�Jh��&c����m��+�Ќ5����j,�ɲź��,�s�����{��F̙T� ��؋�2�XL�ebOSa�j���E4G6�.�X��[�����9)�.z��q�u^���f�h���B�P5�k5;4n��9��E�X�3��|��Zg|�e������'O�>}���|/���ȑ�v�k���؍��y����np���۔�"����$�b$\r��Ť2�\�u,����'�W�����c����v��
*ì���q�����!?�TR�챉�R<!�����Iψc�C2/Z���1�����>�ȍ8?:�wns�oh��������\�jh�*�9���FA�M�~�T���؅�)�#(��
b�������b�v8����1��}p�(��l���r���ϧ���"2����^�P�L
!Q{��m�hC� -z���sߗ�޺�R�p���Lpٸ���QX�	[�&d`����!b\���9��F��82܈~@�N;����;�T&,:P�Ά�`������u�LXl�ҫ�rQ��#��5L�?,�V�W�w��}A̏}L����M��x��V��1������q�ǊI�A���� �`����@���P�}�T������x̺�y>4P<�7�C���\yȡ,������ک�Q*D�3�◗�H��S\�r��j*�����8`�Xe5��f���j+X񔤐�4,��v&�d5�m��C%�?['J��(�j�ڞ+�X���7i��Ŋ.n`������"�Ǹ9�ɞ��3
Sjq>#P��d\9�lX�"~?o} B	�}�C�*�6�#���[u���^�E�TJ�&%n��Q[�>�R����Ex��=����sn����N(�ϛ���C`�"����T����(���$�*n}��}D�a	)G��k~ԔgSJ6>n�~(9]�g�}V�"g�Y�Q?��cE���j��4��An�y
��7b]r3�*\�)��9��b}�\;rB��/�[�BDĮ~����,��ϐ���nG��Dj����QY�
��=Q@���Z(��}�} '��̯�h|�,��]�[P8J2]"Mҟe����Uʹ5j1'v�m��5͆�TY�9q��I�o���� ��iB/^f��R�@��4����IPF�ϓ�rE �G_�͊�`�'�`�(�#� �_��-��J#����n�,��������������
�&�Rv��i��O�O����jW>��bn+���CTE�@��>�����v*7��� ��B�h�E�yo^d߽M�O�Uq;B�r%b��w�E��r�qG���p"���#�C^�?��+�ט+*/so���FŬxE�
Ϝ���"{BT��kTԿ h�W"�2����6ZZw�T,
���xC�7��<n`bX
��+��{C��1�ʚf��(n��9}ew5�,����h�.�����U�`SZ�eWa�m�Q��MA�,z��僴cC1�3W���`yNIͺ�@��Wz0F-r��@�`�I� y�U��}L��4Փ^Z��r�z�*#!����*l"Ӱ)?�S�DW����D�,v�!�� R��#�&7�uo'+�n@M�̈׷�`^���K�%�N4a-,MK�����K�-_�Tܽ����J�O".Q"�SYa��l��9��X�aM����ݯ�=�<FY�cN
˛�p��N7��ɡNJ�@C��X,��1&c��J��S��.��#g���O�Z����(��`�!�#�ceM'"���Ƃ��7i������G@u²�I>���̏�i]/�6$o҄`�+�5��T�M��չ�a��d;ȜB�ܢj���:J���n��w_��Z����H.f�����j*�1�&ν:�׸b~H�=da�� ��|\Պ�dC{^T8��U�P�ȷa�Bb���_�'�Z�~\�B��C��f����X�\�Zd�'��恗@IY�&y�q} ��Ӊݵ�D�l�[)�1�����qp���Z��]����=��W��X#���%cL�gm5g	ƸU6�N!��Jd�B�NZ�s�ɪ �m��ŗ;��I�
��]��˺�C�0���m�&�ĴF�Lc��Й,Q�_S�b��ٙ�i�^�1¼�Hcʀ2�g������N��ŋZ[�����AZC[U�y	���=
�q��	���~7D<ԡl=óʘ$�k~��C�k<�ܞ�6|]���ؙ�ARZ|U��� �4��va�c���R<TNB�fOAx��S�����~uQ�$�&���l�{щ�.�W�"�fM$�ac�,{Ɣ<��c��/m.�a��;��"��¨\�W)t��Q��KwJ�$:w�D+���<�H��V͑�R($��D'V���3�!��[����4��fĺ����N�c�q!R����K��x:�扅��w���g�iwa߁�ȑG񮆽eO��D=)`j}�&*f��9SH�"K��&}L����,��@$��ٴ��߶�����f�?�S�WA�q~����L
��0���אp}o+ɮ?�A��<����Bo����<ѽ���EO&P�!��G�AZHu�z�YY*Ⱦ՛y�T�)������'"\@���:�3�� ��E����s�E
($X���a1@N�R�vx�|2��	7�U.�~��1��W�����kR$�yC�#���F���QY���<���v����)o�ϲ$����0t�x��I2�=�Rh�ݨQ ������i8Je)9(R#^M����&���dm�H�� :Js[�>/(̊���ʐoi�
�r��&��`v�V_ٝ,����)�?}����j(Zw��kGg�IYפ#.���h��e�nVBhȗ{+�0�����Y��LwL<돮���$����&ϸ�+�/�=���xS����[�A-��=×QYv� C�q��bL`����V<��էa�2�yi2.H���{yn4���l�MV��H@[�Y�lW
�������_�ɧu�A
�K]����HP8���|�}.�kĥ>ّ̇37�e�tR�!�KZS�KBzv���m��ui�ķ��;S�D�������
�_�6`�V[4^
I��;���,M����6���lQ���ED�M|1c\�A�7Q�������S5�ԉ\Nse�F�Ea0!ޥYNl�iN����%��3R�Q�T�E]t��iG��n�"�ެ�n&����^�z%YN{J1Q}�.�ą�)NF&������/��q�I2Y�C5�P��ê-z�o$���ay�����ڜ�L���Fme�gr#,KT�΂�$)���2����u'�0L0�JiE�D������h_탢�Z
^�,Wf�m�xl`��:��l+n�'
c�Uu��t^�g`k��D��3�.*��{䋘�oB���܉�Q�h�F��Z��z롏J*G��'�PP]v�BF��'@_#�@>��UP�8�dԀ���Ɨ�W�x:1Mq���/�N wh@�GV�?�۝=��9Ti�-��%Ol���a��I}�� �[�ǰHG������d Uc�|2�V#r�j���ҟ2%8[tR�sGx7Q$E+��DI�q�'>��Ԝz"$X��w)dg�i�[�f�0�ً�;��s�'j�&�w �?ѣ�V���/A��!C�цzd�@ԓ�S ;�(��n�<��TN�AX���Q�t�#�q�ϣ=q�س*e��A@�f;�@�Ϭ,l~�#Q&�&��K�As�
��2�j�W�w> �#[l5N��xy�<�PQf��ŐNpgZDHc(�<��s>�u��=�ݞ@F[<T)Al�g���~P����!���L��8�� ���~3^J$k5�kc�3,�)H4�%HÆ��a4�v���bѶ�9f��a�Z�o}x �.��,���:���L��|���>��̆'�{�HB��t�4ޱ\��FI�M1�b,5"�CQ�3�j���/��N?{�i��p�̈́�W�K�O�X�,X��LH7{)m3�)y�1����Ӂ�PN~LX4���L�7s�γDB��l!�X|X����h1�4��5�B�"�x˦TO���{i&H2K ]\;!k�KR_� M��@��b颣����:�PH악�(ӲX��Z>[����,�Ɇ\�
3ݔw9�l�C����-���Ƴ"�iC*��-�!\�3JT3�G����yݠ�� 0�q����Z�:�Ǌx�Dz]X[с�k<Cօ�US��G-^�2�"y�lrU���`����d�`��Љ������s	��d�g�}h���:*��M���K#`���]MB~���cjX�{�Q�9ׇ4>�����������X#�
�4jk	�ȍ.�R�.�:N$��Xk�l��������q%|�n��&gs��7TNtɯ�(old~�mޫ3Ej'��Ħ�;=˨j�2P4���#;�؋�)�j�/�W�܌��>��v/"����=٫҅�oF~'&Rk�47��_D��!��T�/|f%�&�j6�X��K_��zF�@�����%鍭]}W�̨�QTv��o��.a9�+�D�X��Ƶ�f{=Ω.�q�@���y��H�BZ����g�n��x���εI�nΏ��SH+q�9�%��D�&�v�;`�A�L+���t�,�6��qT5k��}�R$��?:W*���Q���$�|Xԉ*�Y����P��`FH�l�}^bڴ��M��!�s�Jao��j�Z�IV��U���� ����HN�^$'��=�b�o�y.�RX���I�&8,E�G����[�ӧ�H2n�D�>}�jLoԌ�W�� h���&��ڷ�M!�/��Je����́��%��IQ%d`��"����3W09���뫶C�^H�@Sd��ވ'aKN�Զ�koycZ�a܉� �Vk�����X��-��k�4�7�>����&1�S�+^�Gże\�YAA\��O{�i���y��k-���i�9�SYLh��6���(>�N$ө)����Ha�q@��I"n.�R�Ʃ�;В���^$s�w9��qc���{�ND��KD�� ���jW������<�h��p��`�ﱊ���D��,�`~"�=��O���U1��6p���4�s�HЄ�)��"��[kw�O¢0f�/5gI�;1� �tbP�e��O���k�,�� Q��.���b��3���>R�3A|^�Mw��?�et� 5�+��՟�@X>GYx�_�$��'ڽ�fK�jQx�i3�2j~u�5���9b�|nH�cG���L�e�4L�j� !z�#�P�6Z�V�ª�ٸ�w��t��Bq�����j" �1�;� ���!��1��B�%����k��̈́�Y�l��w���
ǩ�ym=~ۤd4��pc�8<ؼ��{��Voe���$K���j����w����,2�u)���2Sey����K�ĄM��h�Q�8�wܜԍ���ݞ��
����q���O����H~�.҈$��i�+0:�Ar� "�h22�P&��6�U%W$��7r��F�?T�M��/R��𽘶�э0�|�l$	��.��$ٕʳ�z�0U���Wgs#�'���^Cc���N���v���H�'BUx狒����t�i���W-D�	t�a�Q	���9�0���Lj�b�#��S�`l�P����tc��O���c��ɜ�����۩���tc��OFƣ�p�I�u��ǐ�gR��xyá���O�*�tO���.b_Xt�R_���,h���P\,�ߪ� ��#��Z�����X��*�d!��*�*���oʖͯ�����n����r���'8=�c'F5x�C�Yj�xu^"�z����p��_��ί����9Z���CNN"���������@�C��]� �n�ٻ�n��H&�ױ#M�V�¯=��cs��\��wTY�:��"��H;me�೘wT�}x����i.@�S��^\g��䍁���T����ԃ,�h;�|I^[y^�*�
��S?����vlk����qD�-$
�g�����_�N�W�~�媬��P���2y9s�Q���h�s�ho��M����x1}D�}?��T�S��\���^�!�#h�Lb���Ċ���D���|�ko;����"`�H�H}5���a�������G�3ۘ�i�Ej�p�,����vS�` ���)!F��?/ޕl
��_�a��&>!�c�+�j��@P�P�x��R˳�z�Ȉ��f��llM�v���_�ڬ&����;�8j�U�Q�_��~ H^��M0,p'�^��.j��q�Z|=3��Fh�}��N�/�QmQ�{З(�٪�V��Jxg��ǉ�@V��%ښ_7�,����jҔ�R�웖c��y���k��l_��M�T�����x���s�ӯ:����`���&���e��-�2���tB�w��Ɂ;�K��`O��ogìj�!�iΰ�h�C�Eb�~��L�Sy[	�N�W���Ry��~6X�+쇾څ��$c��<���6�i��y�)�e5�e˾{��,����/n��а�OcM�$�a2���i�E2eI�.q2L�.p/���IY���N�c8�u/�z??ӻ����'�%�"NP�Ocq����Mi�~@܃CM{��+�9�&��߻?:7dV.��%�t�5�4����E�����Y�aD��*�9irף��I=4�>�'�8���-$�Y�����V&����7�k
��oФ��/l��B۶����F��shOJ����h(X&�bH� ���.*�B6s�9t���_�ɗ�<<�su2=�?��gT�VA�I�Y��qsi�qc��K���aa���PqࠐMq���QhM��)#�R�h=h@�!u��+&p���u.�'�"���*W�\�k}���0�,��N[<Y���_Ϝ�sG�	��ܯ^���`����5Z��IςH�M��H!Z��e�Aܻ1!c\�$S�ue�j7\�x �Q�^m��O�+.ξa<�:�:N�s�/�상+2K<23�.A��vsb�L�q������W*���z�9��G�Q�*�(�Ҝ�ҋ���t笻��������7U������|������Vb�����ez�� �W2^b�ah��u�?��:r��[4M�#�C�mI���P{_*)����W�%S{�e�Jn v�9�z1�o��q?BJh��B�yk�o �=̎,�L�{r�W٨�׿�:�T��l���WNvҒ'+�6���\�Ի���{�oE�ժ��ǻB;�,!:	�{�����a*;���1jq2Hi�=9��#	�ro���-[LW�"Q^'��
�&wW�J�MaN/��F�Q����vgxަD�b����MF�o���ְ摵2�}�W���yf_�����h�ΐ�./>���S;�,qy!�a㋼��1a�*ی�bea�%�=�\C�a�ǋy0!�A�
^����<4r �ޘ,�tr�N܍�>�q'`���BXD6^e@ ��#�/�M���׾�@�>�����t���8V{�/E��O�8�-��Lc����Z�>8�p��,ql�9Y*z�D Nr�͍�qS�A�v����k:7Z�� M]L��DWb��Td�5	Uf�$4%���1V�@�3d�Z��\?Le���0|��׹����ӗ�۷ū���d������C�� [Ȼ�p�+T�/П�Y{��<��n���!K�[^ ���WӬP�oX(�=Y�V M�X���1^�6��9hd�0��/ӵFv������0۹-PԦ!.�tT�|�K���N�_Ѓ!FK>$c_m��y��\��g\��J�p�:��{�6�A��ٝ� �d� �;(`⹨dPD��4�R�)-�'2ti�Y�<c}K0����[4}O�RT�v�N��ȗ*áɎ\����H$8����!`�o�z��f����[z���(dZ�3���1���9��B�i�h5m2�*V��.���~�JT杝Dl	툶R��v~��qP�<b첣G�A74��� 	X<腨5P�jր*��'pcBpE��C��f\P�t�i�����&��y�2ncp���O�xڱf�k�-P�|b���e�������`�<m�K�,ܪ��.t<ܽ��
J� "�c���b2+po�����۵YC!�9ϣ{ˊT�H�ϵicF;��>߹�7M��o��b9m�Q�5�lO�6���!V�&eϐ����k�%�af�?�;���� ��h᣻>:A��>Q�b��.D�@��@�#�'#��A���r�y{*��ts�F��+lV#�k�(�p�!��PGI.�]I��@�q4��p��V�5&���P�Z��O|N�m�����-���������tqi#K�3~J��"�e��=��WQ�^ûb�jBw���s$Շ��x|�8� y^)��?���� �g�<��aK����>?�y~E���f�0R�#`?�a7�W|�tx���μ�����,S���Q.����C4r�oW��[��Po5������5Y���f΀�3J��-�)r���$c��
<�[��+Φ�B��*=q�����YF�s
s��Tu:J~��s#�u���Tʸ����~��n��|�Aǥ׉�j�C��4��1ϧ��x��[��m>k^1�i��TB�ާ�Q�@{�Ma*@�*�%�D��ݮU��YA)�l�Xv��ꗣ���^Z�q���OBg	�����+0����c�G�ꃎ/���)H�ܟ���R=Ԡ���3t�	�|���O��Q&Z��'6a�A��R�6�#aB�w�b3��^P=�F��h�||���q(�� ��Ok��K�oD�;�2#K4�*<?�z1Q��|9r��i0o_�}Zo��9)�+Q8.�:�5��s��	��S`s �A
j�{=�t��k)���r���fF��8�)�'�+�4)K�r�tf$~���X��
e�+q�	��'6/{"_��S}��1����)	}����^��;/�<�y=��m�Tz�$u�ʫ�A�Ĩ����hVef��\�b��TC��֑��:���H�3}C����������v���s�?/�H|Fߐ8iW/5l'J]$TOY+�B�K �xD��Hf.ۡw}I�S��
(z�����1 7�>�����ķ$4_����� �|���4J'�b�����PJ�x�M�bBgo��˯�?�� ��_��i)�T��z��t �`k�@MRG��swh6�%�͹���������D%����w`���ϻ���#�ꠒ�k��tٌ��TE#߅�'��}�����ٜ�*�����T��4GE�$�&CL5��>|� SW��\��]_Y|M:�i�В�Y.='%��^�M���p�Le���к�&�w�M7r���?ܾ�Z���V1�e� �����%1�/4*µeLb|_�Ad/�,�s9�@���6�fȡ�椐(!>!�w�$̄���~b7�@j���3��E��|��i�[��؅9{�'�;e�\"�󏖜l͕�	�� ��_T�<�����h����̹	�},�n�A��!�m{�EHy�f�&I�no�5���դyf7T��Xf~>�ƧX�'�����=��0 �tNCG]SA����<K����r@Ԕ/qr6��.�+�x"� !w�^�~u��g�-[�	���\�BWnj �s��������)���Ye)����]	�F�y/� �F���t�Pd���
���p.n��H�զ=�D����46U���:}wI1��p7�ˀ�����^�Fzy�&��� �h4JM�&�/����좽�'������~Cm�>w���d��I�'�6���ޘuT~���1���8� ��=!n�������C��)�׮M��>�?i}o���P*�f?��̱��}0��Y�w^i�q�g5d? ��Q'Ɣ]�_9�u��r��x��?[��0����}�uw�/���A���5�?.D^��`�������ߚw�f���%5ˇ_H�%E�յ�hC��d/Œ]T>��#���)�
{�+'��Hp�F�/����g��^��ٞ&��pRS׀�oz�	RXI5�a�z�;̹)Ġ=�Һ��܄�%��h�hϺ7�=F������'>0�]D�ɪ�yBQv����a�GS���τ��@�=	�:�����7O	�{^��Om��顺37�e
/�&�0m�F�q�,��������N;��^w�Ế��xFx$ �_3����p�X��|zC��
ml$8�#յV��������������X��!��USSz8"ō���KF��;���¹��������U��]Y���{�t�\>��Oگ�'O�TA��+[�v���^`��.�o� ��\)�G���D�6}��~����3u7�W�&؁N�C+x샲3�n�O�}�<?�X�o�lB�b��lp����&m��< )��֛x�n�U����/��$�Y�36��$�T�vf����_�K��� �p+y1#)rr�**�/�+d6m�����N�Aб[aV_�t9�Α��9R��F��,i��F}� ��O�Cc�t�ф�WRG�Gh�Y�6�HW͉�2xӞ��WUE/R��&�P|��n���"�{X��bc�9]/x_�Z�4�ܓ]���~E�n��vi!���H��� �K�%�3j����W\�2s���pZ��Tb�X��gV�N�8��&��7�kVZ̦A:OJ��ar�<4����(�,h$��""�^#����v�l%��,'��f|�U(墠df�QI&@�*�@�艓_�T�<���b��ˊ���u�q�(����lPE��8W+����ul�8}�Z�"�����/���,YK���M��c.�3@Y���3���.�4y�� �TZ]=0@���U<�9���Ɗgg%8��d�:v���m����?��2�J�7�9�o����<���*���I�,�@��aq$�O���B������Dy��xZ�X7 esu�4i:z	E�b��/b�`��z_�,|�N��p�wḊ�-TD{�,�2 .�9���}`�q�]ʾ�K���?�#���I:]�	;YX�� ��D�l<1=�V=v���)D�<ш.��ĩk�q�Fe��D1�'�.@�^M!2���l���Jk���=�7��H%�ͷ?,�P(/�]��@�T��D '�3�;qa�Z����������{��]�N��L�y-$`�t�`I�Ji�k��;j�^;o�8�%,�������-��1`��l��;��n����4�k� ���w0�5��h�a���p�̈�&RE)j�Ս&�TTLod>5=��s-	[�{&/�yT_8��	T(�D�(���ڝ��8y*�$:�o�?�:�m-��0��ދ��G�J
�������J��N�òT��)m�.γ�Z�C/޼�x��e03g�P~G^���.  ��)Lw�R��m���	�扢=~�2��KA;W���3���0�i�>y��"���tbߖ��A2 � X�!���S��ۉ[�hm1q'1�0`� ӿa����KP�̛��ncF�E�OS��S��%�7!��>����7�ۦ��V�˹coy��g�j.^������s�)j9��*3pX�?� �|<0�h�E�l*���db(�2�K}�wf��E)��*���f��t�ZbP��W�����4i�{�����,܇�j���6m��[��)�}Mw$�_~OF���1�C����(԰�v1	�ӑ�[w}��.K�DjВ4�0�0��52w����\�TBw��XOo����, =��L,�`���hƛɡ�<''�]3�(��Hv�Ȅ�7��X0'������5�T�}s��Ʉ�� ��sy]�up�+���I�+SubZzL<�yain�Z�aޏƺ}a���E��o�7��f�� ���1A叠���^�;��˙�ޢ,֑�����b�#���'մm!_��q�ؗɞ��ٌ�B��]�����G��R��{��u»���F=0�f��RS��;,�ۡ��E�4�`a�p3��!�S�L���y��-���çL|�4(��^��T�f��wi��bOs��z7	{&�ȣˆL�璣Q���v�r���G'��v�Jr0��c��왓��E���ff`5�z���#QDY7��˓�qd�h��RQ�7)�P�65Y���2�Zh|�EƦ�\H�x��)r�r�mk��u��<Z߈Ү�����g\��7�XF�X0�.���S5w�!��5�^��d�"����e�>�ji��Ȑ�W(�olMd��C�9h��҂G���!Iiv�EY<�k]W{.��kJa-��\#<:��hzb~���d2�ћѴ;]��gߞƷ�/�"�o-�X�ߕF�$�"����}6�9�V��^�^�Ȣ��l��W�PHJD��ʙX������oa�X�N:<��V"k.�<�{�;ǎYE��X� �>�$A
Ǔ������Θȸ3��Q�jM�S�w��\��ں���$5ָ.d�g�\���u:1�{�,��s=�x�+��=�.dU���a�@Gr�2ƃ�þEM����z4�=����T;��]j�e�q�,�T�Y|r�D���B�A�ۍ�'��Y��f�b�c%��� �k��K?��5�V�bȣCVF���#˨)<�TB	�Y�N"4�UiP�� q���2���ZӹF��Z����jwt6�,מ��(:_y���B��a���I�.�S����'��>:��;��#�Ms�p߀^0X�!}�h�	-gĂ~����uS��Z�|�BBǥD��B��|��n�5Q�TF��+?�ʆĕ�k���Ǭl�}>(t�+PÞ����=�"���老
.�'�s�
�a+f�h�n��.R�D��>�0�=�B��q\����q��[=�!��,K�ΐ7�9�\Yq�e��vgwV��Q�T�F^�����WŜ�]v��sF�W��L�#��/h�&��Q	%�����␁0�g62�/0�򩨓��8��Y"/������_��|#�����r�&������[�S�l�9@dD��A- �`��<)�K!a�l0�FvcKҞ���oH��dI^��!����*���/�9�9����܏�σ��f-����_�-��0�p��\@Z�ԧw��R�}	���Lа�l2�(=N�ؿ��
��R�������N5�;>	j�<I����m����VCцfFy�Pr�uY���a#2S�*I���:j����Y�/`e����<�$��$ĒPB��"ǩN���%'�I���a�@r���f�$�$|jC�D�n���8��{���h��4��q�P���醙�/�G�q	�kы���>�SI��|��v���#ae�]?�'k�Q�#czS[�g��q;
~���,u�d�  �=�����$�F��`��Zc�Vg���ޔQIW�+7�4�Iͯ!:|r�!^;D�h�� ��T�{�L4F��rՌV����"
�ʉ4�Bik�;g(I:_�3/UPш��_]�t1�����K�p修�
?���}��ޙ>�R�Je.�Uj��3��bBy(�2$�V�HЬb�J���Ĝ�� �e��TK�ȝ����b��̌���/T�lm���?m �#@��y4��se;��C�x����� !�,�g�o��m8֚��v
�/����R}=��!�e��E�{��Z���L�8���N�Ƽ�r���A(���́���qo==W
����=#�N�9Z1Py��0��K�4�Jc�c-uD@?c\�-��a�H�M,��
�*�UЅ��A%[s��O����Y�rk��#�T�Xa�1�%�����elu4d�����lS4��]
��҇��D�f��[�&�Q�0۬[D�'5�w��u������m�O�?�f����ЊU�0L3�&s�����芝�>�?¯ů��/6�6@	f����d�W�H�~U�d��RV�%_���lr�� ������1WбVpt��#qւ3��agw�n�ã�M�Zl7E~�T&����Uֹ�^�e�r &��)���|��q?�k����`f��屗g�RCh(�"��EA��KA�B���6�C��j;��VL���U*lGΪ�j�Ҋ�}H%ňK�	������,�S�-&����ohƊ·�+�ց�zԺ� �ei�xU�QB�u�r"�V��#��G@�L]�fA�k�h�Ɲ��n����%��b��}Wz���>��R7�9l��P�>ӑ9kKʬ��P+wP���H�A(S�a,z��X�� �%e�KXn�p�}|�^5R�㩉AȽ�dj�Zo".j�!����,+VsL��4���8�����60u�iz�~x�1t��?��Xv��RKf�z��_��2
�
_���"����u��>�
��U��}���lw_�4�O~�=�O1L�;�I��2�����F�gH	^%	ϛ��e���oIո��ue���a��ތ��7�BaϺDj��I��HH��!����?^�i����z�+Vp�I&�T���<����%�@���C_1�}�/;𢑎`%+�h�֓�c�T���>e�g�v�<������ޕ�QO]A,)	j o�'�S���xw��@�`����x{�XYtӯ���P���#�5p~emr�q���Cbͭ��Q�A.�WƐ[��K*0�Ֆ�Σ).��������ʈ�YEO7!�(��D/���xΠ�E*��cZ��l�I`�x [�y>Q3��4 �_a���?p��J!�P_��Y�5���#�D���c`�GQ��-�[� Vt��v�Y�O��
2
�ځWz�I�����`q��X~�l!SKIF^�^grl<����:�E���b�l$�2f�f�o���*���V��k�.SM!��,�����$�22�
�YFJ�"�?�F+��`��|�M����
�삡]̮��W5�M*8Eދ~��\�x~�R���.ݷ3���Ȕ��%f2�]`����������NZn`���=������D)iS���ã�~7M2DJ] �߿1
�|�x��e��'7֦�W>�d���lъ���+\������ψW
 ���IM!i�X��S)�Vgl|;7�fC>�\�/ k���~�h���q,(����r�zd4 �J��R�ŰVQ��w�q]�<�X��͆@?�\���*�l^�=#�ٵ�_��H�?\/]��osS�������
l^�+u_�-��1�>����p2@>����%2�iѬ�u��e�'pY��'��x�?�u_�Ze=�Gu�1R$!�u>ٌȯ[�+$c=2�B0[�xD_��~ك���6>����H�6M^�J���l�.u���Y��Q������6D_���m2p����%��5�����������2w�ʍS9�i��;	\����2�W��� y������(C�
E�ؕ�?�-�E�~:l� ��̬~�aG�je�����ҏ�����E��ٚ�X���k�q	���Jf�Q�@��4ɢ@��e����o&8' �b�(�ɨ���p��"kd<���8O�z"��^�UH��jL��(�#{^���>$9�u�K�AP������"�rU'%��'�C��w��\���Nb��PmdI��Up��Q�.ZT|�b���9��^h:^5q8��,:_y��>~ga͏�^p�d�����v��$�Dn6�s;�����(�m�[��#pP�FӒ"e��p-��P�{ V
+"�x��.��CB�Ѿ�4�":1��N �(����RD`�b�@��ahț������Wb��ü�+1�U3�R6��D�j�祂2jk��+ �A� ��L���Ǎ�0vO�t�qr��_�7R�a�kx��w"�/��g��[����]�����4lY �j3u�f���蹋�Lk�15���Q�4,W�"�s O��a13�-%��Uo �]5)Qpq(ֹx6M��r�G���[�'Wԙ�=�V!V]��Z�K���}�O���>Jc'UB!�6�4qd����3Q6�etG��<�"1�3�I�)v�v%�iIuU/�@�<�.�/F���Bd������T��u}���S
I:DL����ԐI����e����A�\)N�������'>fz��[��u�O�����Vq�D�Եo�ߪ��;a4`S5j��myhM�b~P�+��n��^�nyY���zB�f �����q�x�ks/9����5��d?� V�p�����j��V���@ހ9�
{��jxdQ�q�SE-�F�mh�o�5�pqr�t���~��V]P4�"�|R�j�ǅ�,sԊ�8��-��[�x�F��_]g���q�%����+���y8��e����s�*��6#c�Q"�i�%ɷ<Nڤdi�膃����d��H��-�@���[K��L;����:�Ȫ�xkkl+yiM����F��;�%|�������n����N�}Bi�ü4N�֞����dx�1�N,ԆY����O.(��&H�i譬�&�����Ol|���1�E�/+����t�Q��v�Y��XEn4�Nw�5/��A�B��4�KxPj3��F�5�0����k�Nn���Y�/�=��8�j�_� SZ��F� g[4su&r辧��86�1�K�as�e�a�^;�nc��2ŗ�9�A��k��[(����j�.�n_l�m+��?�����Fjh��t�;f���r��P{���
.�Z��X��K�"�����$��O���M�0��<O`Q�ɔ�F=G֪�v|�-Sw�*�(�!��y#i�-�|��m��K��[e�c��)�F~\=T\Y����m�q��e�ȫ��!B�}�Ǔ�lAk�\HU����4�J���>L�n��o/#�y�#�T��Ӿi#��B�����W�=�`YS�����P�/���|��#T����AL����R�,I�ۧ� �G܉���Q8.��H�P8��C��v�(�f!��03NA\�]�\%����`BZ�a��0�OO��.�>���N�V����lo�R�(ZA��ڗ	��W���'�TD��z�Y�<��a�l}FoI/7<�K�G�qd[O�럈�_�����2�~�V�y�;��$�=�v�	�.���pkd�|��5�#�ĺ����H�t!~(�\��K�ˑ�z������^U��ժ���,��Ḟ��cJQ�S[���(��u<vkIK�P��X����;?�X�۔���U�:db��ػ�O� �"�7Mt��c��>��ɡ5��qL���g��YJ�����1���=��
.uч��b݉'�+`70}/�4���M/�,���v���o�7v��9]�)���R��|~�����B˨h�8@�8���1�����VG��'�Y-���m��nA�/wR��[�9{Et->(�z����e?J���ɛ&�\��za+`�V^���z�CF����͛�����[����k�f0y��-��Y��,���abȟ�Nb�n�����'�G�uҭ��Z(��H�X�M�<?`$�z���=��ll�Q䐎M���{��U�E#+ �m�o�g������~k�`���e��#��O��8�#��g�����b~��*�y�����`�����h�{!��y�I*`�PN�
3u���H�Hr	��-8v�qQ)aV#IN��;�xt���h{�$�<��Gס�]�'���9IJ?��쇪���y�3����d�H�u|�>' ݚ� �`{'F~�V.�	 �x�Eӌ���(�L���I٨�����h�
� 	�Mi�I5��ufO��	w7L\K�R��M9�5���o��rz	�@�!��CB�/t;��bQy�b�j^�JK7��G��$�Eo�p�?,>$2e}ަs	�ck!k��s����
�p�v�p�\ �J���&�m"fd�M��F$�M�5�g��	�[�ή��_(�F .���7Nr��/�1ء*��G���`�ksE���nrJ���������dG!��.g�z�X&�E2��V�~���QG;�p�`�f$፰x'>�w@F#[:��&��{�ǆ�cΔ{fk�g͔��Dq����Ǡ�g�8n�Lg.���Ձh!�3�]H��Y��T�R y�5�dH0H�>wQ+W���ߏ�{!gp�9afO�<W���V�e)$¬N���Z8W�Ov�,�R?���M�&�r�N���A��\{����׀���M~�΅]�R� `>�^hU~uX�^?U��3����L��,f��\�o�;(G���ôqGVgɹ��(�5�DR���axmj��C���?��@��F��3ك%=Ғ�}�D`�'U�n=!����ț �-����Ta����[�*��%+��H5�m��҅����d�#y�z�oɜ"Ψ�h��� {�P]S��߂f�`'��%Jo��lU|��	g��"�pIKݩ����/"s�������q X6�$��b���S�q�� =��-Z�X���:_����یJ��Yr{�E)������♤�<2R�>��~W���m�9IL㠢�QB���On�w����2�L)��[��Vuz3�*��}����v�r� Z���)cT.Ń��ug`S�O$������Z1�>9�б_��}��w��?^����vJ/�w�NǑӱ$�,-�,���� �]�/���̻�s�{��zՆ*;��c*n�ë����{-��!�cu�[8vǘ�u�o���Μ6nT�RѣC��4љdͳ�o:���+R�+}?��5)TPK�]�k;������D�3F,>vY���)]�|l����(k��'ˉ�&�aC�;�q~���.T㍬�� )�r>�^�ԥe��I���ٮRa�~S�^}�2�@��N��u�����]Ww�,�E���e楳�~ē�ihi�q�;"'����^�!L`ahrd
��M7��CnZ�>dB��	蟜�ֵd�xf���ƃ]�h�Y>皐�D�E(6H[o�l[�E�=+�.�;H�XЛ~c��K��>HX�8��^����nѿ]��?�9�Ϙ-z��Z���/fx;���#U���Ĥ�Yj��i[��>cϖ4�nh�[�{����E��+�d�$�ߩny��Lka+}��Z�((��\�Bg���ǋ`��5��L�Q�q���*�⾣�f�՝�ͭ�P�@&ߠ*��6cTcc/,��,a�VG�x�Ę�O�YI8#�&*Ǐ�P�&c�z�g��lҙNn��0+����]:h�2=D�f�+#E�:����ƛGD��� ��H�Fj1�XdH���H�n�k�q��ȇ=�s�Hni�����'Z��
�]lN<��#�C(S��,-���#|�eƏ�OWNJ����L)yɰ��.jQBO�y7^ܡ-"53ۮd���_����8k,�	o҇}�e�M�	��yUhO��G�ā� �z(����h�7wF�~y��0K�J�X;�Ec����d2Ul�|u�h�1]Z��F�g��I�Е�`6Q\����6�T�eyzK�MmN�T�[�d�<7.�7D��I~��T6��0(�dc�V؁,l�++��.kq�^��vY��v#V�_��P@��0�U��F1��O���F�)���c����WWe(y1�����0��]��㷊Γ��ª�c��]��x�`�F�
�B�N����H�lT���[�Ai<�(���QO����疛iI���&L����0ؒ���dt�PH�X�3<E4QNz�t�P8w��wۙ��Ys��}#��R�ȪP��q&�a�L.4�Kl�%�|H����n(ͩ�-~����l�<I]Af� n�;��'3Qa��mΣ=_lKm�� �z��,��Z�2�p�f^U�sߞ^��:�7�n9��@��i��kޯ5|�a@�
��W񂑕�C2��S��KEq�d�_�s��3�����,s��>)�j3��[�,b�8�0_qDm��S�,�ͩ�J5���XU(�V,�-'���-fe�o��?�ݴ�XW�[��%o�FOR��-a����M4"gu�1m�|*�4��2"���eb0ry�R7���b�ց�H�
���cG�V&V9�`q�/ZH)��a�۔�-|$�h�Ƌ�
k�ؙ��¼���{��=����+#S����PG��m�* �)�H��wbu��Iq(����"ʌ4oCt �l��G�I���(�$�$��I�	��U��α�I�ӓ�d��`�L�ܵ�9���8���P��lu*1��My��i6�Gu�*
W|��֛�x�j;bB�!��ݪH�6�F��>l�6��*�XJ���M�f�u�/C�s���9��E�$���]oM�ىtf�'��sE��@sz��|�@�4|)�t��W��;�-�;�P�h/���mv]]���e&�������.R�iQ�/h�j��+v2��ɓP��ٮY�F��/�O�H�eЇ�}�V��\�h��|ǤC�}�գ����g��b���ץ��#�U��� �/Q���x�ī`�&�=�s/Y��Ǳ/aҗ-~\�mKY��� xr��]�>���o`~c�,�K��C�� �<=��R�
�8�I<��쎍6��$ڇ�w3§��4ӷ�Xsn��V&R+┠�̄�@��Ke��f$b���ud��b6��g�P�Ff��b�͈�楌Q
F銑h.7�o���Oz�� �����
��Z�؄��)� ��t�����|����+^��d���tS	>�<����H,�踁<�LZ/l9��Lյy;`eFx��(.�j�ץ#�i�C;�ә�H��n�Z>���R1��F�t�������@����
y���lQ3_v����YsK\�l�}�Åb���n�@M��}=�����}0/�إR����H������m�R�S����N�!���lӎk@�,�n����� /VeqC4�̏�`����(6Fn��j)�ﮒ����l��b$$"�(���3\���ݽc:� �a�p�Q�i�]�t���DA�Q��.�6�2_�˝B���������~^��N�/�e�ʕY9W͢�G1��M���:�t�,:��PE��.=��PrZ0��1�����:<q��Q�	�-���r�^l��FS-�S���O!�G3$����װ�#"A�yoa����"E�-�޹P#(
ʄ�':���"�V���!��
�Ӄ2ۍ!$���+�����pPn@<@�0:����z��u�2<�9U;ʕ��ԅ��`����z���>��O\9�R"%`V����� jU���OmX���#Ȫ��6�ʭ�Z��(g쨠���*�]8��1k�Ç���{��Y�����hd�Z�H�{�[<ƅ`���F��%HZ
�M�MY)#��R��v>p�s~A.
6��9��x�Ѓ,�i��W���[�y(<*!��!���<��6	%�7��&e��s3��r�������*7���K4K[0��L_yi0$��jb�8KaV��]p��]4vnѹް�߿f��EǆP� ��X���\÷:�}P�0F�|��æ�0��#t�T��2#W�����v]0�Q̢�-j�U~"/�K���UǪ,'���a�{Ҿ������t����� �0"q_^��qb����'�{\YLC
 ��m�m��#�ڇ�ׄkXRG�u�U���h���*��gL{4]g��s��t�j�t! w!�k��� &s��l�&��,N1gAsa�G�)�uc�|�d���
.^Q�P����}l��D8@>��i\ �m���	�w(�N8;�*��DB�
�S�i����I鋿�~�FĘ�����V�1�.�|�r�E
�pz"�?��Yu�HJV��\�6t3kEc�W����~U|4��w����.���r��(�O#��}'�3�?���뚩��\�P�w4V�k��f���e �㗖�[�:�I�jh�����W��4��3�9��9��n�23>H*t:(�}��s���!<�{�j�+)� ��?|�3��/\z��+l�?�r7+f�Q��Ğ�zm���}.����"i���NN��-�~��Խ�#G�/c�4�q�ʃ�a�7w�c��c?��OV�q�t�,7Ձ~��S?#'@�|�p����\�=�2/��MS۫�e��>�b(�I��h�G2\�GPi$�LI^��!�[�[�ϱ-(SZ7V���XO����y`��?c�}���$���g�e'MƦ�R_t�|ιᨮ�T:z�pe1ڷ��^�y�t�y)��8kn9pS���?G��s���h	9�׷߉��3X�%�は �TK�T9-~��t��͐�'���4�m�zè����zV��#p]t����r�o�v����-�7E����م	�*wB�6����"2 �#<\��K���χ.��)Ѐ��0�{�^�l�4���ؔ՞-)iL�oI$� nQ}-O��)@#� У?n�} h���j-xj���lV��d��9[�p�l7���� ����~��������ǔ��Y����v\|���I>�����
t�O֟Vڤ���H�[8���Ö����,�eɧ�����5���ƴ4�D�P��"�����-��r���>]f�0�����-,j��j���SF��1�M�@��4K==�|���\|3�e:>]ԵR�m�:$KOMe��{���T���[9�\���k�'���O��e�>v��A�//��f
}i���9�^��e��
��n�u�\t�?-�f	9]z3m�������r�G�IL&--���0���'�J��~�еxaL��1�Vy��^ܽK&��5#�I���rA._��F����*�� Y�^��R]cLyd��n�� -[K'Gc�|�(��������-haaR����|��XB<�� �c�	�j�gC����c�<��ɹ��� �5�~l���i^?�_��j�a�z�T�J4�Ejk��|�-o���3�H+�P�(�lE�ÍX�L�mE���_5��#���Tָpp++k@H�7]J��k $-���>'�f��(3���	}b���DTAu�Y��U�r �=����T=K3 ML1 ���E� R�_�F���2*�-��<��/�B��ǔթ�+�J��Un�Ϊ$gT�������D�zZځ��
��ѡ�^q�j�V@�-V�g��Rƻ��L��{;�#	�
ŝ���.8�	ܜ:���n��ᷘЖ�,v�@�:o����oJ*Qb*̅r�˩|�N�x��>g��)��V�O���\g|e�\V������*�A���턪n�����M%n��'��U�0�j`Ge�����hچ�����ֿ�V�^�Wq?���ˮ��c���:�&�+`�]�u�=��]�C⯜��bj�.���Z���[Q_4֊�� �O�q�����p|E����ɺ�� }�	zN:�y0=G�V�Ys(�!l�'�5*�;��\9)��kBX_N̄��m߄`F�?�ŀk�Ǻ�5u��1b�h��kV�~H��`�qْ�Yi�K'd����gr�z+x
���|�k��&y:�GD��0j\Ghh^R��	�O�'���T����e�=$�r����o�u��EQ��ͺ��2��·���L��RWz�� {�}�e�.����4�2�_��`>x�$�
��ۢ��܄�t�Jo���c���M
��P����ɘp�EX��,���Q��J���k`8��=ܰ���e�)��i� %�ŗ�_�g�e�.x�ttC��̗�hJ����^1�6����R�*#��i�!���vZ��:{�����p��I\�>ƥ����Y���u_���=���Y���xؿg��ޔ��O�58쬡VU�zB�`�!�@��C�m��&%i.�ͤNY�H�o������V�x�-G���<��Oڰ������Q���}?�f(�R4����F��������h�Bas������}J`̙y��c9�\§��Ȋ����%X1N!jKـ��n���S�n2��ہ���e���qnQܞQ�K�è����~�9� �H8����KWX�� ���{�-y���fF��|�t�-�)� {�7�e�)5�{�@Z��OHl���۝!�	� $�֫9SkC�T+\ܢ�����%.Ɠ��
��}��+��^å���r޸/�mnB��ⴘ��"rϺk �`���yv��y�ƪ����8�6��`�!k���.;��pqq��i�j��L�m�s�r$��,�Y�%����D2��[ގ�Q����FT��.��YU�Q�d
YV_a�(�Wv�j�G]ΟI�x�z�|��� ʺk5@v�mr&��-����e����r�=h��W���V#���}
~��޼�����a<��H�YR��}~�z�2���xl���29?jL;'��Ԅ��1�E����^���ւ�VR�)�~��H}��7� ʟ;�n�Rp��؂i�b�3*7������>��BGG�`h�����3�>P�F�����Q�zz��'�Hn<�W|�Q,ch>�#�5�H��e��%�>�m%V���#{!�~�Z���]��'�G
T]%X��j�+����ߝ��-H�Þj�(�����R;�/E�6��J[�����q���[n����م�R�y��\J�R&���~�@o}<�����K%�cYb���3|��J��_�ߕI/��<����ޮ�>��{�<Rr��_9����ȼ�52vW��&�ԡ�f���ե�E����9����J�� �_s~��D��b���z��蕶p�NVY+��~DC��R���c��5�2@�n�V/�pB��%L%�����<y�<�9%��0���ל�p&ds���a��KB�����;a�U0ָܽ&����Zu�VI#6�-�7���	���§�p��\@���d-=28�o�B��γ�O*+$��í%�H���V��k�t\����@�LۿPĦ��7�{�/�gA�3��5�����H���f��l'SmG����T�����Y���$}3j��YՆM<!~�S�(U;������S��5��6*�d%�^n��;G�L��2�F�Q���IC)�Y�sH:�8�e�4�Zg�WրCȒ�:41H�w��?�;�(�1l�Su��P}����x�E?M4Z��#�Y�?,jkc�{�j-`�|���$� 0 l��������#�	l��P�ݟ��Rx��k+�&�7����(���LU�\O��κ��X�P�.�B[�Fᦲ;��^������Iit�+V���S�JW'���șs_�9��2�H]��s�zP�K���!���d@9a�ކC���6�*ڭ����ǂ� Q~�%��m�_��Isʨn�h���۹����{$}01M�9�m��¹/��f9��]�z���[/J<�-j�N)�i�=�3��2���:4#��1��l�ms�m�W��xY��1����	<��`)�G��!�~lVNT���wV\K��H�r���w��v��E������J��%�5��OV�>ʩ�~<�m�H|ʋ��ky��8���GFrk�Z�Y���q�u	��Y�J.jM[ԏ?5�c�3���f���@m!(Ɠ7c\V�k_��Q��XS �?L������d�W��	�N�~v5��?��R�m�ct�+cd�[^#2�vI��p�= ~hN����}�B�;��P�.�$�0E���8�:��
R:V���?�-*h���P�ʍ,�2I.�V����Roi{����V�	��7�?z�Hђ^h�c��{4��/|r�xR��OF`��(ۥ��?=*��;<�������G!��U�l�bpo�gQ����[�L��K��t���T�n�}��1�=���Fϰjm�I��<&ʧ�`��bΣ�c|F��}e����5�e��Bz ���p�Dv�s��1�]E3�xUm����������:�P�xz���������Q�Y���?k`}t����0�d��x�����	�q�Xꭿ�{o��IU"�6���+_���l00Vn������kA?!�b��Q�6یN�,3�UƮ�I�X�t����|CV��m����W7���(��eD����ƪ�C��5����G�m]��� �o<g�"o�z�Z�"�e���%��=�<J�Ɂ$���}�v4f�h��s����N��)�+�~Ӽu/:^"�s�"F,!-Y@�]-��`���zki�q��-[V�!y��S���$[Z�Y&ϩ�3;��)�����A�v��g����
�;�0;�&�U��fK�E�K�n��tEʈ�d����4�'��Ģ���J�-�����c��bH�a�� �$�����
�� �fK󀑶*g"��o V�a�W������r �������ҫ2��V��N:�+g�����~�E�0��_��ׄ�}4t:?�W��N�:7����0�if`:K=���p��F��غ�*k�P�xȾ�h�K�q� �x�UX	�~,X�se'�6!u���KJ�,k��6��^�@,��G�m��#%��� us�j�*�X��f
��{!I��:̑�uԑ��hE%;V��#��N��NF��T��*
C��HFOtR[u�Ȼe�S�R&2!$���j�"�=�=�=��Tϐ3c�m-k+�ի��tS!m��|Yz|�i�c2a"��?T����> ~p���,g@�5��Ή��pE�1QWWS^��p�����v�sO��y��XUQ�MY��{�s˃��W���C��_� u�
�/�6+���nY������.�k�߱�;���D�<�D틣2:��p��P+ �x�*ceqv���ڣ~ng��P||t�T�جl��z�[�*.���f������W��d�[�������ɿ�E��/.� �����Ȑ/�[?a=�Ў�a2q)�j�n�\H������_������c�f�_Q�e�3&�(k���B���뉶�([棨"�� BZ�q�@v/���LN]�{���M��yܜ0�M��)F&�����;ڪ�SD�����xZ`���#��МF�"8	M|TVu2����-��^�>m�G�+f�{2�\�7t�q���ky!��ٮ|����F ��Q�Qm�_^��?�e��b����)��-Wh:u�����Vo��yK�1w�DX�`���'T��c�x0b>��T�`5�&�ڱ��9{y��x-�ǃ�-1m�`�K�"���@ug�
m�w���a>4?�sd�ֽ�pN�0*�v�T���
(��u���i�w*S�J�SƖ�Xy$���*
��W���+M��1��xgk���T!�h��W�c��U�E�G��{��`�4c��\rx��L�V;��f��8C��������f�bM��T��[�1�y�
V �e���	���w�ƭ����SM[t�Qϳ%.���5�5,֐J)?�� {��+To
�\�[���Ϡ�CJ3��[�U����N��2��ZF2:�$X�;^��+�4j�Ow\�|�������U7�0�L�*��V��'v^�`H�������)��dMM�'V�j�5��H�X����l�+�!�8�GYZ:���  ��%�#j���+��^E�/�dR�ɸ�����N�����oE5���d.ݗ������mzY��{
'7$K�	G.j� ����0��� n���03T�d��ؗ�+|2ӓ�l�:���s��eE	���m�b����M�e��oN�FS��Fas_�/3��ʧ/��H@�x���V ��O��`��FO�Nq���w�+� ׭���]��RZ���/�ѷ����C>��w���4�g�V}DP��D4����?:�H/~�5����7���$��2"M�~~�ک+V��K��mݢ�E75��~[�$���$��d0쑋��~<���jl����i��bTS����NƁׅ#�B��8�y�.��+ox˘�5_��0�PEb��Ďc��ȉ<�VM��EښhY��K���q��`Sw�����g�.�A�#��ċ��!���*7�����>eܣ7s<����ÿ�7���Ky�c+'�<
�����Q�B@ �g�)��ű3�:�n�w3.� ɯ�����P��^�����|�m�$��w?�[�"enⱋ�NADp���Y�����R4��K4%��r�&^���!q4�����^���q(�g��Hh�{�G�pUi��?�ǀ�x�"c����3O��7i�ж�j��-.�7�v>���L+��9��߯̏`�b�W��6��G�HJ��T6E��4e�g�
6P���z�E����?����s���j��Gd�K�$���Ky�|�PH_�^�]g�
W⒇�\��1��[k}��]����B���,��>N4�5���^����F��ʲ/�i�|�CD\$	<�+����?o4n7]Ѝ�G���:D/t�`dƁp�<���-$��7���C�7k�c��쭌uN���TH��-zA-��Y� ~ԇtGk���N��@��&x	X�(�� (.t��RXm�Sp抐�Ep�节����[�[Қ阹��&ѷ��G^8�R��A �%��W��B��:M�]�0�����Au��@x�M˄,�VL"΍$�I���(BF��Z�E��HV�oz���)�Z�<b:t�j�\�3qq���ۇ4���*�(?�\��Y���~^R�	�/^���'�Y��+�`u�Si�i��N��_^i~�B�w��Jb-wer6b�wNz�ﰲ�S��ѽ��pUho��u�b��\d�a��Mq�e����R�uS�����5S��B��Sf�z�S���6��#�7>��ӊ@M��J���dx?#�}�Zw��?+��6P�������#�a��Aϯڧa�v%�,[q0���H�u ���RΟ�EKV�B�!E_�~v���*0�j�����D5j vm�^?��TԽ�:=�|�5������9c�3�.s$����f�����W�X~�0�_�)i�ȿQ�/?���zѥ��m��r�V�T��C#p�j�!�2$��r�:�������Ms(�Mh��+�ߵ��ܶ�k�@ԫh6�w�z�}ĭJ&EJ���u���y@x��GѪ壼��7���U!M�c��k��o�ѝ��(cA���ޭh�t�/��k���
r���tf�[Qz�۝��h
ݻ���z+�͎׻�)tL� ��t��M� +�����iu�s!�����߷�Pq������jss��9���k���Ջ��������7(�m�7\cV����/T��4�h��E�^��	���f�ua*'YF���%��SO5� Zj�3;2�Z]������Xp-��6�5�Ĳ�B�ȝ2�����?���s���}Y�u�O�n��z�cf�8��y�#N)*"���b��;��,�'��e���>��m{!"��{�sz~:����!�U��	��<�J�v&�5=���JsM�X6ƞ5���������o!TO���%F�f�D��ڒ]!�[}��:�	9U�!��HIݍ�� ���ag��\:r�
�N�5��cZW3=�Uұ�P�
��.��#�û��HH��S������p�d�m"YBM8�(s�9):G�=r���>����,�bs͠�����7 K%�+����@׫�L0^��o�	�FK�[m��{V8��3 I�L������m�S\H��]ژ���$���/I��"9_�CC�Wh���rf�o^u,��I��`&�L=42�i��Az��[�Tq�O�.L��d*'3^?N��|�$���ZnYC���B����s����g����p��h���Zo��rx�Fg�u��+����b910r�yG�D\m�-/I��DP��Z��~�b���!�������Q��y�r��#Yl	��� �,J�>��n�!X�5̎��Y	�B��Z�_��3B�'�)?����?G��E�o�l��aC'z�e�:B��,�Y�W&c�=B�,H�E�}�Y�.u�8$����wm���X��=�v���n��s���$��n8�;�Y�@����b�1n�A�%o�Î�!I?� J�K'M��߾?c_����[��G�'����?
�rJR
�8�.�Ϩ�q�}������zA呣CHQ�l��޲Gq�GƇ2e�냭�Gݚy� �C~��;c���I!�3�7Fw�R��V�kr���� B�z��A�ӥ��=��#�5�˿<y��g{�����v����[�-�����Z�$O`5zM��H���REud-j�<�N/}b��zB�y���l�cr�m���?�s��5�U�4�����B���w^q��I�|���Y�b���_�j�����ձ�!ob��i;��:�E�oiW^��`�������\���y�o[o�(2��|�1�鶎Rx�|�De��:�c�l�k�uw+^�"��f�@� +�QY���B*�ި@�~.��l8�"Tr�m�5�!`WY�f����w[ij�8�}D�^�R^BNd��n�"�F�]vP��n�aÍ�np�:	-�uLl�X+:=�Gs9(�[�g�]ְ
k`�����&���4�Ұr�DMs��z���b�\�d��ة�7S;�\O����)�[N"�U�j�Wf��a�ɑ3��{X�2���s;�G�Tԙz��{��Q9�%>N����D!~(Y����Wt��d��j��
W�f"Iwm�`�D�6���5�����RR�/��3^���W�+��{��4��z�R�BӠ9���y��Q2� ���-�|��󢳜����l�]-^����59b& �M����JgM,�j5�H�ފ��|(�����gw��
**pG��3�J�~8́��-�x:Q-]d�<��l�yx�'yj���{���� F�����e�a[���r�����m<�b/�U\�R���R`�4i]S{!RDJ��z���lq���;.<)�'W-lM��銫�e�RIҷ��#|�������Y�+��⦐�T�)c�F����/ަ�qPx]uK�[g���� �_���1�Wԇ+sF�ʤ+��hm 9+�!~�<_>)Vq���j+LLBҁ�g�mem-�0��S�	�.�1Э� �19�r3%�?÷3��D�X'� ����H�sMlLqi�X�]�4��Hkw��uΚ�=�21���}��uq�U*�)l��)j#��Fn�>��g�P�}��,W��,��ȯFc��!vg�ѩ*r͐�o�����Y��ՠ�Ϛ�>{���	!e_^��(kn߉7g�H� )M�o�O5����F�L�@��A�$
!t�xj��l��t�y�U<q��@i������J(�!B���Y�*�,fv�cg�4����T��+Q��Ww�7Y
y��ǅ�.-�����:�H�8�bK�X�A��#�S��lZ�vQ����҄sޣ`�z�G�M��(1+� ��w1����ݱn	�N��ʍ[�D/|��=�����Y#���f�P����X�.Ż�O5p�����f��E��q�B(g� ����>��M̒�Q��2�ܥFn��)�A!��_Ȇ��!����M�-"$�f%ȪT�5�Y���&o�ټ�ڃܧ	SW,�\�M�&��:"4��6'�b�<὚�����y]e��d���q�lh\�%�0�"�=�5�v'ĕ�^�d
�.��BYg@�@�& �Z��v��C�%���櫬,j���7w�a�ҩi��|r�JLz�a<?�	�M�4W�p�EˊYC��jB��`�L&��H�&�3���iek�>N@��R*
~ޡ����a���؈�y��#��^�Rw"?��O*j��_:�<Vw��.�������m��O1�QwzV�o�1�l%�N�����$Z�S�� bpG�G~BE׌�`�:K�_(�
b1:P{�P��v�'[����}��%��>^ݜ0�=�'j	��z}�
�Hn�G^��ŏG��f��͐
o���ۥ�^Xl���|�{ds���
A�M�/>t��ܳ��@d��^�I1�B�]�k�u�x}���P����2o��5C�z�=aA�IDv6�J���������Jj�G�h�_+;�$��:o��i�[W��c�8Z�M^~!/j����@A��K�g��n�;��ߓ��Ew\C��`��s�E��
 Y T���&ˇ�wڐ��v���<5AB��o�#I�>��!ù���F
S�f0�ү;�]G�����\��pq��"�}v���6�ue�4�@c�&���Z��QU��
.���O���[�.5g�ƟɗT�pw/N��9ҝ���05r��ֵ����p���!��X�^�V~�5+�z���F���qڲV�9��ل���lIMC�J[�T��Ԕl�0U��ďa2��s������8����� Ԫ-|�-�EQ�^�S~��9��z'1-h��+���'�P�zg(V�|&����=�;�[��s�����ݒL�����88�-��;�r�<hy3-{�I����E	����7.u��
ę�'��M5�Q �#�
�%h���!�Pe5�_\�Da��՗�����h�>�}<�@��Cي�g��t1��S���񥾞�Q�[p 
M#G�Dը!����E����8�V�5.��{D����9��Y�탋L�N�2����S����:��B��-�P^���+_��瀓�ߩ�
�r���;:��8�n�������o��rq����Q�mb�.��m��x|�j��ұi��p�^�"Z.���d���I�Ќ��v+=��#=�:���p�Ȍ�u�L&w��zf���wX�ay����Wt�Iy:�V�$�.�yR>�_'�G
�������g�PcJ����FƊ�{x�;�? ,��ՠ�e:WZ�Ӵ��'��D�M�A�V�� T�q��*���n�/z�J�����+��J�}X��ܸj$=�j祧`W��%�C� ������~c��U�d�ᵆ{��*>͆�|�ϗ��H�`�b'@��x�PN`�ɻ�ޯ>�u�G�n�N��)�C�Crc��J�������)}/�`j��;ظ1aQ��ZJի���/4���7����������@{i
����~���ℋG3+�<�	��Q>��DQ��/1�p��k��Fn5wv�!Ԓȴ]��/�'>1�
޴E��� `�����P[.�b�#dD���x�@�z��f�X����ĉ�����Qa&�m� 7MW�$*w�{�X̑�;Ԟ����ed�mD0�2d�;"��ZC-���p6�\�^�Z��|��8�Fى�/:�ٌQ�,��4�,����R$� �c��eV~FX��o%D��������d�)��@ɂM�;�喈�!�V�.)J�I�ˤ��+h&�}lS���;%�=�uɴ|
{X�`C껴\/�O��V����|t=[s/%<_��[_�Ք��_�8�]�d�y%��r3k�:��sQ!eۡ7� f3w������
Z���Υ���.����q�d~���lè���� ^J�6�V��6݆yɟc�	@������z�n�)���7�hN�޲.�Zb�bsZkӺ��-��PkM[xg��t��^3w=#>q���RQL~O���IAQ0��fa�M29�[��г Љ�H^��Ö��)n�jEI�~7���r��%%|:�F"��ib@���%�%|���̺�*�`��-�5K	��䯤�=�ԗ��9A��|�c�-۬ZU�F���޸�XK��h�]�I�uI��M�ɷh�r�YV�䓒]Kܾ~�_����B%��S6�͟Oxz�1cv��r��"?r:(��{P�bB���e��=&�H/����-���A|]����n4p���}߄Z����[����v=��s�hjT�l[(�lhh�a2x������@>脈K`��Mo�=N�+���{�dFM�5$�`�":�?;���J,�� �*F��|�p^�+�8#@P�Q���kj��e>HϏ�G�8:]��;\2����.�l��+La�y&�����Q'A�Ȕ����i����iv^s^���۩�6��C��0��BxV#�V6��U�	��h��0�����e��	�4a<�%� �_Զs��jΒlӚ�ǲ��Z��BɁ1m���^�@rA�5)[��`T�F�5�0��f��U���P�CYD�G��y�A�y�[�=
t�"HX_?��ޘ)US�D���b~��R�*x�j3!� ����b�
�齡�+rH ��y��߫��'���R"�oeQ�a��Ҍ+S�h�x�6H�/���l�
�E m�; �6�Ti����>�9�u��gg�y�����ad�a߈�Z�n|$�P�p�7��K,�\��\8Ī�����7�u��b}?���7{��ؒ��tڛ��1��bv�O(,��b�Rgz��T��W�#-2-(���K�����C5��[s5DѠ���Q};�akCk��NF����[g�Ec��b�U���v�jc���`�r�f��]�u���ٳ�� �������+g�x�(mx�_LryP�M���=���mt�_KǗ�;�:�׍�	��*;����阕��t�&{L�[��������[��oC�yY�0��G2�ޚ�v6�Z��qI1O#��}>q.#(A~߬_�+�x�	k��L�͙:s�(=��ΎD�c"��	��sYV8��f�ME��1ޥ8w��|�ϫ��C!؝�|��w��_�Г>Lm�Qw�^��i�a<]z�@"☠�M��Y��C��<a	Q�}��#!���>�N3h�7
!�3{D'�t̃:/-����1;@?�c��۳�?�O���2/ĒӢ~��D��0�z�������F����/鮔
`�pӮ(t��W*/���QJ���ٷϫ�Em���[�����H�)B9�Zi�

[%�$��e�ɭޛ^:�~��7+tc�����fI���}7.���fN�jc�����R�D��J�i}>��=#�����J,��맀ڄ�5��Y)�#����^A�ǈ���JZ�(5P�ܻi�;�NT���w�b���{g���GO������x�t˼�P��d�{X����B��W�׬��Sm�w�I��Y������7��IH�+�(�e��P(�iC.f �:���C�4��-.s6 �֭:w��ϭ<�;NӃ|ю�P1�Ц���8B�����'~��������0[��ǰ6<@ۄWn��J�|n����7�x;jC�Y(�:��}���B6�����y�u�7*��!������5�G=GUf>�#.���t������Ѕ��do!*�A��b�r�N��Ho>8��4Aj�3�l��C�PG>�)��T>��,(�[9:��9T{h��mE��uIɚb0[۬ɏ��,(��"P4t��	 ��J?��rt��O��l��D�Y`��f"��>�ܰ�b�"���W�IF�єbum�����lѢp����;_e�3(hw�?H��:h�+�����d3m) d��r{�d�8�^ԕ�	5��zy�Z#ٝ��Q�zsmYc���u����6����g�E�l�1�Al�l�\��!���V�± �N�+��H�L��#xB��5��Iy�O5�⿩Ȝ
�}�~�쥅ԅy�% �|"Ysq-DR$�j��r�E�`%Ep��]�����ʅj� 1���n"}�˷��zD���j���n�jzh뜏����� /g>H�vBE5���.��Ub-����]ϤK�L-�lf��r��DXL����T#��Ǯ�����>/���`��F%��S���|ćc�Rgn�����E�E�!��C6�ò!3�ȡ3AS1E�hYޝ�������=�r���%@�^p�N3@�=���:��\x�B�Qk8RP{�HX>���v��Ҡ�n�f@��G�o�u�y�hf�=����o��=6�o6���&֕�C�r��壵+FĻ
"d�������O!K�^��q���������4]�:h�edb{�O���C�
�:��N7��̦� ���7�W����=��%�J=��c#�H8��|pQB�[[���&w�n-�+Yb����t0he�7���n<	b"�e|ZEuG�*=�7���
��f�.)i}�]��1��.���x�Գu�Y�W�e�>����ݗO�T�Y�<��>6`��<!���󲭜��9\�!�=+�7�6��up�[S��*�*�gf������@�8hU	#�6 ��1,^���{b +;��-� ��-=�G����SE
!�v	6T�z���%��H1�������+90nS�c�a�~@���m�#�GO[l]{�6О�}��r���'f�8����PhϽhO�a� ؓ)�/�׻C��u��mRj���#�P��t�P�U
jї�<	�~�Ki,�B�3�4����BW]�rw�$b��ש�j�!��m�Lw��xá1��{0�"Mu�����U��LXf�1�QQuWP$O�?kZ/CC��UT��.t��L����^J�+�U�@v�R�����?�B���o�T��Z���ix���8�|j)ܬ�1��+�t��I݃_��@���%�L�#vZÉmJ`N���`������+ ��^*�/�@�r��$6�0�����s��͒���1��ߛ|(؉����Y%�(��D
�3R����N��8�S@����X�BM)"�M�~��JhþX���@q�3qiN�Cbҿt�osay���X*���8䆦d'RO}l���BV��um�[�W��=J.�*��� �E
�)w{e��a-��zd�Iș�M���·oM*�ѻ���~� ��;x��\gQB{�$H��qa�Cˡ������=�=T�v��m7¾6\*�2��
vDA���ԬV�PW��I3N�d��c�i���.�
t+���v��OS@*(-�~v^�|U o�\�|U`�雒@&�(���_�!����ۯ[T �r�+u�8j�=�j_�{�
E�۱��tT���h 6g�a����s'�D�s�h�F�R�^ٷ�f���$	|~3X������`�\m �lގ�*<�\I,�;�{��S��t���~�Z  ���l�O� �w}~t�ei{Hg&�w���`��S�����xa���fa����N�R!S1��ՙ2�uǀr��������DkHŴQ]��G� mw�B��>�yUZwJs��Ȅ[�	3��� 5�jY_��MC�56X��%��8�<vY"'y�Y<ip���-����L�(�HO����Z��N��?hdA���X5��m��J�1o��6:YcG{�b�-/�َ��b\`��e��
fo��\�\s(:L��B1�$AeV�����!��+�5h��a2�;4�b�G�����q~V���폡G�28�9u�������ұ���~�z^SBAgoX�����J#P*��Ћ�i]~Am���t�Ћ�={����ϥ#'F��I���F���)�4�K�lg���jqp�o�̘%yǩG���q-�k����9�=c���N) 8�G��"6 2`��*��6v���Ź+�a���c36�~����һVL|���W�����*��Q�XV!(�k���qf��e׿��oPWu�9�2(�f��;�q[sp�$X_q)hWNR!�3�Pg���Ie$�g\��
��!�e�y�_I݊��s�H�������WW�`��݆�u ��\��EH���jV�j-�R<��F[��9E�����N������P{�T�\�����M����ˈS��3����R�8���9�N��#Mu �GjhexbL�kذ ���	v	Y���HHa���cp����3���}m��Q��v�L��	��E�`���� -P�����l�j���2|Щ��H�k�R��_�x�H*�#;\�7 J�eV�\����6E�Amdr<w��UӶ�6�|�����t;�ЬEc�����5`f^�ZĐu��-W3����s���M�G՟_����a5�'����F�� 6��%J���B*O��|��I],����N)�/sW-�&
Q=���a.�-D����� ��8��{�yb�AM���u��f��T��hإ(Ĺ��U�;�+�I�(��+]z�5V0��p)��cZg/�}��j����n�($�b�?u@OD�x�L!4%-����[Y��Tة�>�}7:p���t���$d����A�����>�Ҏ{˕a:� [w�	B����E�<ТӃ�[)���M���Ih�䥂惮옂�7��@r�+�Z�fP���Y���![6�e��˦����;J)�0A����}ҙ�f �b� Me|Nt���m��M�}��4^��/�`Y�7j
���]����-�tN���j�.�Ϯ���8�z��}�ݏ���m�%*��S����hCt'䘓�Ȉ�v�����ɖT�9���c9|�L/Se���Q��p@�,��W�_��K�9�䱎8@� MU2��le��QË�V�S��s=�G�̅N���u+ʆhEX�Լ7�]�5��`:��VE���������x���RV����lE�7��>�#j4�C�yѾ�vN�8(�L���W�[M/X�{�������ME/L�M�9-�n�PP��N�˳�}Xb�Y����@Ǎ�[�Y�W�3�/=�nM �i�'lG�P��$� SZ&![��+A&��n�m��EN��"Q�pO�j
�*_�'��'��������Ħ��e=�6��|��`!�A�7���h�l���r�����Yz��EaҸD>��L@��-}��c#;�ʵ�ֈ{�2I���;U�Ab{D�:��J��c[��c�ln��X	C~M�.���fN�8��G���\jY?�(���v�T�,Dꃁ�9,�k�� #Fg���s�e�Q��,b5���qٕ7�����D�Ү$�,���q+�+����E���WŎF��B�z��6)|�;�j�)ل�<�1̐*l�ll�S�oػ\�}#Ӌ��uF�|��Z������eˊ�^њ���-8�_*�<�*�Fج�jȀ�x�EB�kf��pkV�!�~y��U�:$`����̳"̠W�no���
,�n�_D���Z�Z41ǉEQCm zU��u4XH�!��!��/rs����I�Q:nW�`�1���;���A6,l���;�X`�300��go���f�V"�ex�kR�n��t5%�C��'��#���&.���B|:���ui,j4����;��SG2�^�\�Z��}-�&�����H����b�(*��n阺���IP�/[��z��9�M�r��a��˞$b��lIpQ��K�L�M���:���+[F����
AL��q~V�A���W�@b��g��!7eoPd߭Sߌ�(F; ݾ<Nd�`�P⫃�FZ��v��
���C�P,��u�颔���MX֑.�����';�Z�bT	\�V��ߢ%-ȨLv{��d�J��3ˠ�s+�׌z��&�:��	�O:�Zop�tKͣh�7 Y����a���aV��R788+s�bw*Bs|䝔:��M|�x���\���Hr���&�-��?�o����z��C���-ܟ��