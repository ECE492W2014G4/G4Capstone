��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P��v�"<ߞ��&'��k%P碶�R�ӣ�sĞ������FY&-揍�2˗/٦��l�=V%~p<rɸ:���f�^^X+�� �I�k�<r�o�*�qՁ:\5W�o9y c��A����Ǒ!�Vl��-b�I�}��Ew����=*�������I���\K��c�ț�,}\��1^1��d��DQ�Z�����{�cCunm׋j�iSG�3���X�3
�?Ld��0�g�wC:��^ ?��s�8�P��mZW2�P�D��X�x��b|�x�ؚ��@��t�\8�|I�Ӏ�^do�k�n������CEN{�[���n4_)�Վ"mB���5�-�.�Rբz�!\5Iو�	M�	�oSh�o�����%��r;�T�?%�>H��%Ya�X�׀o��j����m�@�۸z)��L�m�,51Q������5��:�$�5w��uw�B���]��R7����q�k�%��������)uV�ʦto[ڄ��t
EN�������u t���|�Ѿ~{�L!M�*���m'��i�F/��j��Pe��%:��~y[�-�5%Jѝ��La>�{Cĉ��e��P��	;�ιj�<Bl�|>n/G�
f�������������'k��g␊Kf��Ί�t����Ֆ�}I�P��f�m/'�4�}�^"�t-/����%U|�z��dMO,�w��|d�Z3�3����7�ڶnr4�}��A�1a_1t)�\b����n�����@|P�c*ʐcA8����`@���6�{Ơu�V�H�jG&Ŏ?%1C[RŠR[٦��o��Ԅ�����Q;�/���`:��?���`!�`&aP�,3�J�*�#хŰ��s��&��
9�����R�y�P������:$�G5ZҦ��QV�D�:^�}(�f('��w
�A*I�*� ��ɧC����=���(����X��4�{{����-��/��m�%��R��W�����lN����@1>�W9NP���#R��\=�n)+7�:�ё���]��5�i8g@\M�FW('$F�p��z�!Th[����i�?	��Z��Jc�{d�}���N뢫�i(3JX�qŪ�h7�Pf��ӈPΨ,'JQ���.x�W·cYG�MS��9����$������mJ�؃�D=��#OosN^}�Z�x���:��.�5.���b�(Y �/zZ���]�d�yBl#�y��M��"5i����$�N(ӟj��M��6�/*�O��YD��$K�q�oĎ���EH��L� E�b�S$q�k�5�}�&�V_
D�Rx�O܅x��RZˣ+����B�R@���o)�3�-��m2��6�-Q~\I�6b����'@Ơ|:/(����:�Қ:$)��G�s|�N���67{�b*M���ߟ�p�������y�[�'o��l*7��aBƷ�vzbJ��a8�����~O �Vw{,x4��%6U����w1Ph����Y��/���X��O�R{$O����&t�?�<��DL�52�J�'Q��J�b����wLE����D,0m+ҭ�^69�}\n�ԑ�|����шQX~!(;py9Ҵ~Ϳ��\Zo�t���I�l����Je���7aP ��-���f���%_3P���'�-�`�9Ū���Zw��i�Y�R	 `���ʴ���2��z?8S��9s}���9nAp��2�o���e�8�g>R8��U�3�%V�{�af��S8�'��J�L�Տ��(��Q��t�b}EhBHT��G͓��Q��&��Nw��0E<>�0KǄMzN�}�[�kC��#/�}��ӂ�{)pyr��w���Wr��O㿆c|2�D�*R4���mΌ]G���N&S��{]�j<&.� �HXA�!��6�#tĥG�&Is�\�}C��t�*8���^q�.?�Q�%��s;~DL��>пÇ�>
�P荌j��z���z�^݅����܂����ފܜ���jӒ������/�E
P$_28�a�e��k=Y��4pZ�:�M�v�I�0�q�R�(0����^�8�%'h*���9.���� ���8��#��P6�&��Oh\G�u���ȋ�u�v��rŅ��Z�����4?��f�l�<,$Z���:��]b%��[Xg�͍)Q�>wUlSɜ r4ъmt�fĔ.̫��Kz��QSӶ�ք�N7R��=��MT*A3sYo�#��6<�ȧ�F�����%��)$E�5�HкyH`2�9#lx`*������v�������O.����Y��m���i��6]f7.Jt.'���rÎ�:��^Ee2t��k�G�F�S4"j����%Fl`�38T(u�2l�i5,��`�� ^�Z���)�Eu��a{��Uj� � ��x^y��RSW��J�#F�-�Z�䫤"�BI���-��1(Ǩ}@���Mw9�jq�UT�k8Ҹ̾�Y�L��(���P^D�l�!�\#v7���YxX�a��,��XO�-�x9П�_VT�HVח�ի�����#Z2e.�RG�e�Q� ����'X��6*U3p��ܒ\V0����>rt����ތKEqo��� ���{L'Y�+k_W9X{��A�-`Y/��(�f|;$�]#� O��_���W�&��`��%dC�Ў��\��3D^)Ǉu��|�`P���o.�e�f��+y��'�Fr|��v���g��xq�JV��"�XPT�	r��&ƋA'Z�%>�^�	�g$Jޙ�P	��h�o�жe���#��+�JV��V�~Gbwn05|�#a�yA�6�38���~qh�ĸ4M���|��nQ�߲�M|��Lʵ��Fu�˒��9��h������� �@�kF�Įҩ�/�]�x����\p�O�Њ�=�j����]-�$Q���>���h��{la��jM�=�2��{�.�U�'�3�A2j?���r�_�ax���5�aw�!խ��/;Tv�3���[%����"�C=�����M%�'4!GP4�zX��o��ȕ�x�M��-�^�����<�����]~y#Zn�U���NftW}6�k����@md�����י�$�(o���H�ދ�̯�2��L�~�,}1Ϥ3l�4gK:\�i�P�_a�>l��Y��Q#�6��NRh���"�cVj�4�+�'���g���X��W�)�o����ū�0��ƃ�;v��L�Ӓ:>��N�_���_qnU�j�!��5�B
z�8F�lj�#�F*#���i���'/�s �����b��?����b:'L��k*
e�������y=�ǈ����c�B�1�,�dD�ˋ945�Bv;R�\���'< ��ۄ��4~�S���"!SwL��r��p�u~#z:ӿ�Op"�0���ԋ�����)��`�B<�<u���q��]���T;��v�t$4��^+���X"-�Ņ�&�A�s �ṟ�D哰Y����i{�E�ݢ�l�DY�1���O3�ϰ@��O��2��Ǆ���1K�c�h�m��m���BӮ����kM���_L%�
�%|�>?�[��t�AR���Y��4���������$@��#�5��AF�+�e{�q��}�Ɔ�ʑc�g	�N��T|��=l����� ���<����7#�i�)��zQ��'[�6N�ts������^&�/��2wD��V��v�l���ֱ��4������ZkD�cQ�鴦،@������J0��ų))�B���z����]?����o��UŸ�|�t,��E��;��u!d8B1�D�M|#���^��x�%/�0�p�}����x�����D��D#P[�{�Z��]���Y�P8ͅژ&Guk�X��STc/\8u=(�>̣�B�z[���h��(U�;�l;sW�����޶+PpW�A�Ft���Ԇ�!�8f��{�������)�N��e�5@&����D��N���D��ը�UO��V����ܶ�y�� ���wP�L�Q�]��כc5���YA˷��;�)}�]�ߜ��Q��R[ޡ�%�!A^Y1:�O�q1{C�l��F�KȏO3m��G
 �u�Lp�	K:�'9��>��pe�/{��XD��	�Sj ��eFgZ�pa��I��Lb<���:w|��(�|����|Էh�����ٰ���@��U���#��d4( c���T����nKv��E�Z{2.�q ��Z	c	L���kĨ�5��\܈v8���*�BN�J��u��`aZ�&VEp�+Is!�}t�܏��Q-�>߿�C��oT���y9�e�M��?��¯�g�]�&X´���YgY=�7s<��/$o~�9G�I3�Q�Wj���V������E�{Ca!TOB�ńlf��䭔�Z���=M��Rm�t�6~��bҹ�0���$ݖ��@�*���J���dz����w�,|-��1����ߚݸ�����r̎�|D�*\*�s"�����6�{<Fn\�W���+����A=�Mϻ$���F{5>Xգ�e�}��}b��om�1���jw��q�k)B����HF�k����kz��O�S�T���	DJ�'PwG��4�#���^=Q����C�����_2f/��;���XY��,�u�%X�8)�%���a�I�ɿծ,*���+^*P�8�p���BIO���AA�
G} #���=ds�[HQ,��~`!'��tR+���y)v���w��x�D�b�b���fq�e	,g�M:GM>��Cі�'H�� �������4g0: