��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�"��F9s�`&���a�oq���F�g�O�]�<ݲ����eCL��D���{�5��8̝DFI��Zp\m|Q��
�}�6C���UnF:<�jΈ�2�����<����sf�k��,jڙ�����2��X��Ss�HL��	�������+g?���N�Ż�����|�v7�{M��VNB
��Rs�゙�Ld\��X�'��R :�J���^�����kMkx�Q���3!P}�e���Z�Y?.�U{�RP	�)��lI{tI(S
7ZFӯ�?�"c�=��x���J���t@��{Й�?U�Ցp�õ��֖-Ƅ�p���@>�=�?����5X�U�{a�ٷ`J���/��ۜ?3N��֪w�P$O	���D�
��kx�;¼�KN����V�fR-ոA�ng�z�#��d3>i�+�֫�`���vcs��H�e�벑�G�0��A;?�����7�.�U��~F���v��{%V�{�t�6�	��t�w?�	�p&򽟈u�i�ɾ�
��w���#�������^u��kf�x:xE�l}$bӃ�1�Ґ�@�����-|�<ф5mF����p�i��5��4w���N�������A7\��~c��j��v��:>w��M�.��cq_�,)�(���8��`�H�s0�Q5jqQI���^��vИ���EHV�j����<Hf�8�ϊ��k�"B���	 ��p��>�dl86a�I��c���m�Y��Wi썜K3���17՚�ѫb3lR\-% ��.��ԅ�|��Z����h=_���l���â ��@���t\i%9�&���>J�:�U�P�+'g�|B_F�-�ꣀ =��͟Y�1�Ro�wt�HAZn
<C��C����i�]o�����#��ا��T?�6�&�N�s9Q ������X/E�sw#{	$,�ʏtzn��a��^���Kܷm�|�?��ډ��Ώl[V(O�Krr��%g�����;��,�C�
V���O\1_� ヿI)P�=�6��ϷJ�td�&�Y?j��{&q80HA�U��.2� y�T+ɽsh�|%����?�C�ι�^���(��BAC@7��_��gp�B:�����([V���E�#4�d���'��3��B�C�:V�c�GU��b�8�a��r�P<���P�8�:��֘���HZ5�m�*��x#7"'���9{�k _"tS���d05ۘ�����Sc�̴\��>jEsOÓ����2$9���{�(�8h3Sc�����a�W�v9�%��|ݿ	Ue��Y���(| ��Wr:�����V�KA��HF4�� �+S}'�֫�!g��_x�ޖn�9�-��`�S�t}؄yAH�k�"|T�%�/7}b�8����\:q�$A�����d��6.��SN�b0vE�׏'������Vo�n2k+��Bm�8tq9�����+n�ťK�y�!�T���Z��!}���Eni�~����E�	��i%i}�A�,����a�}Jo�x�=P�h�;��^�=���A ��XE���#���r�*��k[/3ŇN8ۄ�_�/��5;��{���P헢#���T��D��n�r|���|f#qi���
 �4�뾁��o�M�6�ʆ�#x��Ѯ���&{�1
1�2�~ xL��A�b*�xQ��qUo�d�Pv?��y��y��e'7ֲQ�4͛�5^{^?pk!hDf͛=�^���}n9}ZKl~�S����<�|$�VD�x�~�	�Ɂ�z�%�������{���=1P�����t� J�#m[9-�|��˥C&~%ءӂ�9 n1�@��(be�,o˂�u��_Wz^>���l��{ʉ�OvG�T>�U���A.���i��?@!�&�b��D�f~�K��ί��1ߥ����tj!��Ȥ"E	<�!�E��(�k���[��{Zl2�=Ӈӭ�c�k���|��-�t�Y@;�	�.��
3�eAcP�h��ʢ(���;������"�o �k�.�+k7��r`+�h���1�t]
#Z�$V��W���`d�L��~"K(?��B�&}ɢ�Hί�vO��Z�s��~u�����T�b`���1P{k>a��t�z,A�!u���!�
����A.��P��[C�FL�2:���7���v�$�������f��כ&b����ro�$~i��hr�]���x�p8��cu f�)g�����/V�yq<
� �AynV��Xh�gޠ�'�M>��0�!����0&��p��M�`�^ӄ=>C��D����s��UfH�(jG�e�+��[�#��4���"U
����bB�$L�$�(. �� i�̌�N�m����)��+�6�m��7ev���q��U�?j�U�<��6S}�G�	�,�K%R���ih��Z���>>)V1��'O�}ؑ��!$�f�����U�+�<WCx}a�Bn�Vts�?v�}�"MJ��&h�,�e��m��=�@x���ıʶ�񁬝*��8��,x�>+���Vw�����@/�+	�rw,4�+Y�X!'�a!�OK��r��uu�܀~�1��q�Q�(�8P\�IE����#Г0w�`й�r���Cu�Ml�H��yvq}�7���$3 ~aM�,U�`�-�(�J��� �Y�GS�/�Y��.l ���� |��՝Z��4�7�_��e�
Y0M�֍�(�qf'��q��!�CR�M����/d��S�fF	��� �.D7r~�'-�٨�M�tQ'>�K6ʎ����������\t���w_����1����g���y�R]���u����;��Ic��*��y�u�d':�h�^]f�J�ܫ�G�K�N����i�q�n�yt�!���ު�&��ۧ|�܌G�x�)�Pv�yi
I�������-щ\�U9)xPw�o��϶�]�V���9��.`V�k��lH�*�e:
x��Ð|`�����$������c36��ѝN�.��^��:e�_X@b����w-�*���{Xɺ�z˾��E�E�cRB7si�OH���Pm�H�k���vl5fB=�}ߋ��.^�)#�V��i�Ԃ��Oigk	=�q�[Z]m��<B\�
��:����c#�Ff��8Q��[�'�!V�Ǽ殇��:��U�ϰ��s�(e��	�2�SQ[�X�R����Ϛ�lp�i��_I��{��ɁN�����DgE�Ug����uFI7W��Da�H�ϥ�g�i�b��y]�$��x�,[Yx����3��m�)��a�n���-q!Yc$wH�Bgl���b^~����������U�a��$�B�l�������YzJ�k@����w��}=���1��(����1=\���.J}�o�t�<�5z������9H�m���Ár����󅈲�	� �,�:0I���_������!�/m����sl�-�`Kʑ~=��W}T���t��ј��ĕ�B��{��4e��,jp�Cv4�-�����>�O��c��>��<nl�f;�<	I��@hv��s�;b�Ӎl��s�����+p0G#C�v^��g��-�ډ�S�r�_�ɼ ��!�џ�(I$^��g�0��x��_V^�C�K�K!��Z띄-n|�k��`܎��I4��*G;&�roq��+�{�>KPȁk��X��>��Bs٫���%
� ̡�gw���p6��@�d����D8}9+��1`��,~M(�aS@r��/	b�����*mp9�����b�A�F:�`��&i�}pvw��cw� ���kt�kE���V� ��O�����Pq
^�(�Zi0����\��O�_�l��E��^��>�𡜂p����p+�M�NS��j�U��5�XΞ/H��M�P��%z���%i�.!üO��A������@nΙU���0x	�-��^�Q2�,a=���ѧE�	}w]8_(Fwt���Ecz�8��,���ρpM�f+�:��Ş�j$�C�T�A�^lj5�*�|�F�V]�(͔6��&���(�<��v�&&��@Oc*�8�S��b4� |�ۯ;k����� �� �@G�����\f3N�+!\ι������Y���(ֽv���a��z���K�8ìp	��8%E�"Zy�+���蝜�+5��"!��d��z./�0��.��ֺ���w*�E�kVʑ/:�j�Y���1�tlsa�fՙ���Q{����o)kҘp|5R��
�<ĕ�4F2})�BP��>��b��o%�`]L��!(��IZ�2��;���{Ǵ�gqU
�w���S���\n����4V���}xc��T"�{�y�����ky�.��#�~a�n;q���o�pE$m\٤��{��곍Lq�׮5؋���������nR��&���c�ؘ$�0����j��c�+�.�����Tp�w@'x�e�F��X����7�2H:�g�N��)o>F��Z�V�e�+?��,�,	��T����J�kV[9p�_�Լ}���.�;St6�
���Ҟ^Lp��e,v]�#k�h��i�ЌR�O�Or��J(D,��e�n�7�����TQtYNh��Tk<�,ߌx5Vy�7�ޯ�"O�;������H�|�ޖ��xgt�aa��$�c �h�oհ�ˡP��lpԇ���8�Kͣ�U���#5���;�o�=�����\��&���+�79mhI�����)�mo������F<C�w'E��α�o�eB�m�c+
̟��}�(���UzNW��C/�3MG�#����oW�$�ϱ��%Hf�b�8�=���W�}���g�ˇ_�} �-}�$eX�G�'��u+V����v��I�'���^\��N�<��Ot��a]�̴t�Z��Z¨��R����.-�=8��Ģ<��Bf�����&��ۖ6k�U�L���7ǠS�M�t���h[�:[�6�9 ������"�/#�%e�r�mq�z����cl$x�~���T�Ͱj���s������G��𪹖2�B�*��q���0ٟ1�}�P`e/6���:J6����F���?��s`�1@6�ũ���A-��lY������f�X����4�b���0��!��`-1P�����-�-��Bs������)o��f��2��0ޘ�&��$`^�]]'R�D�x��~.G�>���C�ޮ-�y��	Z)�|������c���pΡ��Rq��qm~�]��0��<j����q���~P�QC�;f#<1>�omǘn��傧Ei��(����0�0w_��5�kP'j��&$����)������[y9�r0V����5=Oq� L��W[f��..��lt�]ȫҞ"��}=�l���t>&v�"V'�v��y��h�*����qcȐ�_u	�3MX7�[����Na�1[��	4�������a  ��n�BSK��RI5�Xj�ٶ��K;�i�D.�@r,W(���8E��4�E�mmГr�#$g�?�D�M��~�M�~��*2>�x�]J �b�t9��jW�9\�Bf�M@��n�]�tAZ�6C�N�Q�K��V�����
��^�J�GC�*I{�	�]�%��+�S� ��]rP[D�8y&)~y@�`Y�Nj�ݿ���=��'�M�*�
�A�#���4�6��?F����$�'8�[��#�Z&m�4�D����NZٿ�ϙw�S*,3	�}�X�͟�x�<ؘq���wa8�y<{/��y�P��9f��ܰZP�}�E��5����T�HW~��ĸ�wd@�yK�ڔ�8ԟ��V;��ȡ�z�Ψo�Mm\��B�;�:ׁJ�\���|6c��%�����Тe���
+�V=��pnJK Z	�B.��R^����SrN��L?����l��U�5Cm���C��p�[�N>�w�a�*����	��/��R�z)��	��)��x��ɖ9A���!�-�ۓS��<�l��n�ck�p�[j��=����9V�Sm�j�>��럗��J����0^��w�],�U��G7��+%6��]�L���,l��_���hD]�LN<��[fSE:�9;�iO��сM=۞BX`e>bZ��P'>��59k|������|Rڒ��So���%�
����k��j���l������Tg*��;#�0�-w���1]`�- �
;���dHn��p ��3;!՘.�I��C��Y.��\����9����H�n��T�]yv1�5շ	>N�e���s�g����#l|N�.�
��U�ݎ�d�yAr\�9�WdH��j��"�6v�H�V��Oq\�V�g(aH���!b���$c��FyGI~h�,�6�I��e ~��>��,��8�8N���[�95B5xg��2�S����Z(E��ڭ�C}iG"0�1��ݹ�Ɵ:��bh?F�lW$���,ִ�I4�&P�Y٭	����l���7U1�p��T�d�<���	_5-��Nk%
Ե��&j5��aB˗+J@���",h�q�/D8��BO�P���E`1ѭ/@�ܺ�q=>�������SЭ��~��ݵ�w��ٟ�]��|r��׷o�������H�(�"����U�ի_Ɇ�0fR�H,0���)������/�	���o�FY*����~�,�^�^Ý[����I���H�S��1V��l��p	�LI61|��˗���GB.Aܠ�(���o��L��ǅQ����<�Q�~�+�[����SD��ţl.��P�4��-0�d�J��(G��A}t����ט�+R��J����?�O���ЀN���u~"�{�X�d:;LE� Ϭ��C�] ��mt�6��ޢbwR0nĖQ���ܕt���Ģ�d�y�����7YI~޺藂f�}m���B7�+��1Dދ&jj[�0����t1���K�G#�_�:����o%� i���ǩ'sI�B��d^�g6j^Oq���;I��\��I;�D��i�@T���Զ)TE�_��n80�Yt���Z�_6�S�
z���{�9�].듕���@@�����[O2�m�h�-r0>����瀅�Y*9*	�|�bp��#i�<���O?�\N(�1�t*x�B2�9F{�o�\?�*���_�1w�}|�APbl���m4�8扨{r�s�䧚�v�[���}�)�*��ECi;Dw�N���F؆+�6����S?�uib���Gm�PT��J��c�]A�=��y��bX���xC���A}��4�xT�֬��(�S]��F��Ӹ����Njg찱���<E��;��aFv���9xnN�H��; �N	�e7�=�!zݬ�p���g�a� �S&��z՘��~��=o��R riX7M����RLm�z�!L��Kǽo���1hԛ��|&b���T�uR!�&Q�7G�24���TC���k���2���żLa�4�'�[��z��X~���32(6"���~�`���!5���ME����`o���{~ѣ\ғ�D����R�������f�V��=vr
��5�ޝ�/ɿ���Q���_l��gwKm�lU����o9��bb�zr⦧���TV��r!�G�{�A�Ԃ�V{�Lq̜n�FK����?I_ʳ���n�p�gc_�t44��Y�3��A;V�|E��e6ab�0�Bj(U�����,��2���>0���]?*�z�ڭ���b��M`B��o�AD0���Z��Wx�Gk�i=6-b��2� �A��X4���=�j	6�n�,�d��:狡�G�~g}���-n�\:u,���)�1��q�������E���xM�t��[a�/���Fm���������&����[���W���9!�T��&OY⦂!�ި���B�G�TF.��>L��Ʒc�����r�W�{��T`¨��¿�Nb�'�]�&,OZ���f�u%�0�O�2��iPŒl���M���!���%�!On����`x�ia���X��5��;��1_F�^>��em֦��C�O�k��
�����[H�v/wR-��M߶s��1��4��7�a���H�����S�;p�V�*���Aoq���C|,���G���-�>xw\���� k�*k�}ߪѩ#�Gc�)�Z(�a��fe���ʴLЫVl9�A'�(�%�F�+:P�w��G�fܽ���#���:���*Iz��.0��(����W��*KN+�%BJ��\%�\o	��E�o���L�pn~��ӷ��N�$r 	#|��086+�_f�,�sՐiV	�~{��z�w���@(�M���m/�Zi������R8�m4Oj�>A'��U���d|�ȃ�j�������L��͈�d�S�u� �O���ԭ6ݍ6�هJ��(t�ʧ}u3-��^:uD� ��Ǵ��`�*8������d�9��W���G��=��*�@)4�q��둵+k����Q�&�u��XU�
j�NHT�o^|�9�o&X8@�ī,q�,l+��s� ��iM�bw�]5˻=1����Є'VCƁo7|��Tg�oU[m-*�ǧp�����zç�]����^��ؑ�����o���^�d̯s��
EM<R�w���	�,�3���{���M;õ�GW��˭��OJ���ɦw��q-@q^�w'+ߌ�d,�����e���4�jb�~���Wo!�*0�0�!�y����ARI���5f*EKU�	�#���&C��[���s��x4kN��>ojt��ޚ�h���\�0��'a���4�Ve��NzE>��	�LÁ��S��u��D�F�A�z/
$���u_%�k��)"����#�I��Z��0��|�|P=9iz���^��)�����A�a6�-TJ���,k=�L�T�L
���	�{�z�	�x����]e�n�(�X��b���*oH��Yx�m}btr�m#f��_�p���/��{d!���P=�m�C��R��g�� n�q%�C�E������XΟ���2�!m�F�=�.�0J�����CH��Q���,ǿ�1Qp����?���NzL�,�������C	�ʾ'0Z��^.7�+8���
lj�� `�(��1h��!�!Ձ&���H�0%����v��ף�wҧ��~�/�i��r���k��)����z��'�����IoJ;̹f�i3F��&-mbaX��a��d��b�wҲ�vs7;���!�B��%Y��C���fZ+YK�o�r��jAB�m�pc
 ���V�>����[�e����h̛w�}� �舯��M�v>h�g�I����F`���y�TQ5�1���k��m��*����j��v�w/���^�	�"�"��c;F�H�j>p���if����wl������Ջ����4D�:_l�HJ0�x�T��&��j���4=�7���@����n�x������e�8�/L�΄�)0��S�5t�
{EXɚ��z����hLy��[E�.����4��cT�p8���+pu���)>�D,$c=��eՓr=slH��"ڔ��43�2ƣ�e<��3����,}��$3j�:�1�h	�f~|���b�^w0����*�9V�M-!<E���3�._��!��j�IcPF	���S<9IA]$@�\.'D{x;5���Y%�l�wih��ȓ����{-5��6-�lH����蝟9"ݮH���WH�M
^��2,EV��
��­���fi�����R�c�)��~. ��m�ތ�~c&ȏ
�C:w��t�e�s�/�!?B��ԅ[
�@�O�f~}M�	͘KCé�eE�!�����1A��"}���Q�VTQ'3�QQM�xm;�mo5Xxu�bX�?��V=?0���[��:��:�	J�R��00�!��?@{�{�R�S��#FД��&%á�Ra�S7f$��p4c��˔�ڠGؽ12:�!@$�Y�+�Q�ٟ�B=��긆��\l!���׵k!�Sj�n�QU�Y���,@j���z�(�H����$4y�6f�����
�%-��:yM*zn�۾T�F}`���#*���~�b�W�K��4�nf�;������_!�O�^��}&��ln���R�OK~��`��NvԚG�G`7(��|`�'���i�vT�����Y���t���]yyM���1?iбvk����r^v�y�;�O�F>�N��[�� ���Xfi{{Q�f����%_8��K,�ø�_���@u�g`R8疾�T�z���3Xi�Hhh�lBی��0��vO��>�Mƚ��0L��B����T��ǽ֏"�x1ƭqXqW�R"�aj�^�YI�9�M
OG�&m�%�Bj����,�Ȫ]:���}w:�w����F9���
�hn K.��.I����X��w�5���Gm��W�׷4��Tc�c4V������4� ��G�����kGH� +�P�b!�ئ�`�;�k�s���R�mC(�{#Fc@p������T="b>��<$����	~E5oE�x��(*��U���N]�'�WI����>�*{�Pȇ��/�\��mMi�;�m ���
�
M	�j�E-dH��8���un�~�r;~��;����}'��5���(p��{tK��ld$
�E�߉�G�G��0��=P��-=�*������+�f�q`	�7&<1+p�yQ� }wg_��G��H�~� ��Seӄ�W���7�ǭ��I��S4�K��ތ@��DO�b���t{���2�K��=t>��նγ?e��s���j|���i��4�g�d�^x7�.V��}
'3)	6ɞ���	��ՍJ`0,G��[T���_�CU@DT0*ս�:�e�D��>$ǷD��F�=�{�C�f��5}�E|8�k�&����<$e�A���\�2��c6��K'��;�A��o�Z�Ԥ�1L&�as���\�������QG!������5�s�	��࿼���Ҧk�+�蔳���賲_%V�1��d�8��k�Ypyl6�5*�y�"�=�y�"Z���b����4��H8����'xx���Y��p�ʶ|�{`�{�`y�Q?�b��_���7����)��]毟�J ��T�NyG+/�[٫��	�[��b���@*]ϦZ/����]7�p�w�.�`�Y������Z��E	��t�?�*�S��%z�o�ښ<I;�*��ɧ�n{�(����!�x^�놩2:���{Z�T;U$���G'�����E�XM��ks&ؙ.۹f�p�}]��ja7�nj��6��*�%f;�,��U:��P�9Gf+�S�o�٘���=��5K5H۔���c��/J
DuRZ��p	�M<S�'Y�oS�(Q]�v�;�%h�O���V3�ᜃ(�T���1�Rq����z''
�f����D�hĄ�9֑Ƥ�z�~��dg� 5�p̀�y�$gݛY��Z|��:Ujl�ZR�%�/�y%�=!p��d,���'?fpv� p�dW�d�C:�@0�+�t�˯�w�`����q���tݝw��w��BĐ��8>�Ŷ+����B�$ƀ�(�v�|���3�(rJ��qI�J�/��B��Dn��:h《G�������ICZ�:?A�U_��>�*����22p#�C�}!���]�:u���{�ͧY��zl}z���Qz�����!� �8����	��2/%9��b��䠣)�z޿t�f���U�M���{9��A��K:�[q�0C2Nr��M���8��.���Q�yٕơ��I"�����΢_ �}���L��W����(xB�AI�<����{�^(�	��
���ڄsS�p�_'��c������	R��:��XŞ��j���ԁ��,:L���,�K��C,e�ޣ6ՓŁrez���uATn���P�to��؄�^K�"�)������?�l�[ֆPW=�Jq���f'������5Ű�|"_8�B��r#x������E�ʞc�J���Y�9#E����3�����7��W�v>B-g�K��������pW�e�I�B��(X����X�ǗI2��Ta%�	'���B���mھe��T�SSS����ъa��e�4[<%��	=}#v���۲��6���ja�fx, ]R8t����Sj�I�H�V'��`�}�Tbl���i��vr�
�>J�����,��vD^�"���%$+k�7!�Ȉ3��ŋ/]�lt�?�0��+�o˛r&,p�]�}�;�.�䧸���I�`��ǜp�8� ����D�4C6���GS�\a6���9�D��Ѻ�+�~Fx!���J�usK�C$߁)&vx�*�?�z�1 �A7`זr+-�T���a�s�����t?8�������.'�>�`�sxZ�$L��L��>����,�d/��ƌ�0���ұ���9��ow�л�w	$�K�.����0�D���%�!$xY�I��ibQ>�zTۜ���D}���h'��7�� ���c�}��b�\ktf/�7k�9勫��������B�OA�7T~�@?;ܯ�'i�O����u��h~� ��A��RC�;�U���)�G[�^����7R�#NA��"S��س�_FC|5d����{@]S�(�C��^;棧�q��:H�H#��;��H�|-���&���뷇p���?�@���"^����}��٦��Q��W��e�b� ��*�����M�j�w�1�Q�A�8�I�r5�q��8�����acd:k��^�C�_\�'�TOOO�)�Gd�Y��JʈIGZ/���m|D	�!7n@m& �5T���"8C��@����`�8?U�������P̭LQ�Ϗ�,~Tzq�Y���^�Gi�^��8�Py�Z[������8c"��xS#B�JX����Y�"T�w)H�����gb7���ÕR����0����P_�n(M���ňm��*%p���	t�<z�
��*�i�h S�I!�����U����>�א�>
�	�|L�~I�6�7p��Fdɲ:չ��!��^�`�#�?�2
��&�$14�G0߀��	_��<��!jK�c rakP��4�E�!��s��!H�p�Il�N�A�$�iY�P�m<OE���ǻs�.hc !�V�ҙ�U`W��8���:�'����UxPU�Zi�Ϭ��
޻��R���>�i���#<|�]h�|Ɉ
�G;�'@2���s_�f�}"w♖��xp�9�{]�zm�L������j�V�G�Ī\|� �߸�4 �>|��h�,��Mh~�/{�;���f�l
��(x�� c�L�aC��b���8v[�.�dB5�.xxqf��!�G��zv�CNW��-�����O��¾`Z��$p���p��F�Xš�]ie��ϸ��#���>'��X�/,�(���.� `��.zr�a��џ@�;H:j*D�>�Ϸ���C��΅�k�W^!��De[�-|��U8��+P�G��e2ڪ�ȕ������g��Q{_q�� ���{x�t*�"�9H��"P-آ�7H�7^���DC/�#v�]�%~8��ȟ���^su���F�l�Q��դ�(�	��@�`�����6i1}߫{�w���h���@V� ��k�cd,iyh��������;L !�r9CY��h/t֛
��PK=�0���HF�/�$���������l��J�����c�������}�Q�?��g�-��	�$�0!F5#"�z��
� �(�8��̳�2�[��^{6�^n��b������-8N���M�~M8��U��L�E�ƛg�ř��O��^��T����ɇ�����v9	G���d������� `*F9Y�r�
ap�،���,���WgȞ�J��"\N���i��$�nv���-�7�*�j\\�H�'Q��%��Z��P��"��R>���_�����jqX�,6|�ըՏ)���dԕ�7��~R�ɦ۔�,��M���Ʃ����8�]�9�:!�v�I�� ,����{&$�J�P�f2;ln{ym�G,%���b�%*\�A��5��0��н���Psީ�W��#@�]�e<@����\e����Y�sGN��gH8rh<���ɽ��'�>p���q��7�!��g�K.4�"�����*��6w�,y	��1�E�w�w��
�C�(�-ψ��x ����uW|�?�<@*2��ê(��>�g�u}p�$�����S���?�x؂��2bNZ�H$�I����M��h����սG�rU��)�y�]N(�W�c)(��<xgJi�2�3�xc.ͦ}�t�-�>{�:,��x�9)�	���]�tB���&��-�����7�g�Ȏ4fj����K���MėA1��䉒�KhA��Lķs�q�����w�1�A�L��a��i�7Jx���E�xx�c7s�0�*�|4y;��L��'iko�q�×a5�j�/��>^ ���w�aF��,�th�֮}j�#v���c�<S�ɼ��!%��sI¦�뇯6���Ҍo"۹
��s֗a�_�Y�J�g�t�n
��3$��:b���z�#����Zf�4�\_Q��)D�j����'�E�X7䰠/;N�NA�p���X��Rj��*ƣe�p��F>:0q]Ji���#��k���� i�s���}�����¸`�삆��S�&D8�n(2��/�YOٚ.������<c%
��R�C�|�=*J�.�}f��q��i-�3ߊ��z���1�{NvLXܠ,�P���/��XF�>��7���7J6�2J v"�W�YK�Î
�j�:�r�s��If��1%��9��� .|p���߲9�+�%@9�j�}^Đ1Ϛ��kt=]n���]yw$����e�J�W����y^�9S�"��y�����ᇝb�v-�f�������&l*>f�$ނ�m#�u�=���L.P���;��#��*R����� ������v�e 8F�nhZ���n�����o�����
�v�t�G�g�����3�W�%���X;���c��L7G��*(��C��ӻ[|Ⱦg�����g�C� WN]㔇�QSh�{
Yy�/�Ǝ�?|�y1��fy2�v�2�*��jn�P2fY���S�H��*4��3O�EO�0,��p�4Z���_j�;�����=F�����0�>GF�7�+��l)_�u�=��\G�0�w�o��4�)�����d��y�T�d���[b]�h����q�(�  �>~��<���B�M���`��X�L�΋jU�O?~'ܙ�5VW�o ���u�gĸ����U�>��n]��rY�V�E�g�o��(�U��wI��.!�����n����p$d�f	-j	�3��A��H�xmQ׸�凮����ꖞ 7~l�V�E
^OL����+t�H{��B�X��p����O^��گ���7�HTo�T�`�k���a,8VРb�!WHr���+ˇF���`��j#��ֆl5s0@_��s��z��
��_AWw���A�_�L��G���Be��
��W��^Gvsa��X��U��lX0`����~,p�������i4���Y�D�X��_�!m{��:(�ո�����x���!�6$!������RC8Ν#�B!�`T?OT�)�P��\E�*[��
:0r5�b�EzZTg�.�y��Z%\żP|~ڂ��!�	٧$���5K&Y����C~�*RGs�D0�6�����DI6�уҳw �%р�\K�4eʓ��-^;a���(��l�:�N��Pi�m�Nx��&��@ؕ��)�o�Q����s ��}� Е��7�vc��኿�Q	cp�~��B��X��[h?�R�9�k��B}��z{��[1�Y` Z�>�@GO�H�b�,1�o6�������d�#ԡ�G7�}�!�q�6ǐ�/M���z^�V��ܧ�Xn���:�9�s]��r���6���R�C�P4�	0VUE��]�3}D�I�,u{A�T�����F��_Ud�5��|�h]�xƆ7���4���(9r׌ג_n33vF�9qT�d�z�PSe�\�:Dza�$���+��f;��m#������Skco��W�*����P��P޴)��a%�����g��0��tR�����6op�Q..%�Й�qt�is�cc~�Z!t���E;]����r��G�P|O��C/�.7�n��
H�M��8�
c�g6��L��Ic�
���}�A���ҟ��,{̓�|a0\�E�1#�5�m���D	����8^��7_����GY��*~�9l#��I�Iq����Po�۟Ga��5+َ�n��z���OaH��ew 8�C\����*,p�w ���h2M$?X�Ę=w��ͱa�=�D��#�HT�H���������� �$�u�q}Dd��!�1l���ȑH�=&q��l�በC�a0�M�Gع-���)޳n�k��<7Rt���>��˯і����ze�G�-��B��8�1n�����h�ʴ�'���>��S}8�9l�a�H*�7/�ɏ��1����fʍP9�v�s?q��A2��w�d��*(�㈹Ѥ̔��������N�w�IAa� ���p5��a��z�8Ro[|�xY��u�4.� ��t�E�|��
�蛪-��d�0�#�rK����OC����1��	��������\�NE�5X�><��_JzU̬�y�W�ј(�(8�pD�[2M�Ai�+R�p�Li�>x�΋~fY�E��t#�p�B;��y��T$.+h.�\���:8s��p�����␾��e�0Xu� 2�{А�u9�}���IZ|bRӎFQ�w��M��uq�.[|�Hx�Y��Yo��	+yɬY�9v���ɉ�1;��{�L��g�c����ٯǽ��l7�!��O�*S~�$����9U�\�-�@�!�����؇�7�s>������F���{��^�h*��;���t�|�e0��Wg���Bd`$J�X�Ĉ��]���t_�u��[�u�Q���q.�I�nt3��1��E_HN�<���Q
r_]D~v}BT�����u��q)�}2If�L�ƭ.�E_��d՚a�VW9Az�	�U��>v0%n�n�<h&T1�ܓumt?W�c���/#�g���h�X�5����3��ʂ�p]���.cuU�r�ٲ�>+H�`���J`:�8�c#�O�2vA��r:�i6��N��<��lԇ�҅���`�Y�D����9�+��Ӏ����Hτ?Ŭ�&�F8�빳�8o�%WI��2-C�������o�\d���KR=�IN)�������Ց�z�f/�0�Ll�b�����S�X�}�o�jQ��a����|��=q����%��旡��.U�.����x��n"7�+ʂ�W0a0�D:�ф�w���|��(���Vb�ul�V�xxi0�-箨x���I���\{�I�ӟg3��ǘ�3�1+�ne쯊���I鈟��l�t�� ń������炨�%_�˲��\���9���?p�뼤����#^�7� ����,�n�Xu:֭%7�6��5���n\T��m3!]��|��`J���Z�X�X��"EǊ{�r��ͭ�g�x�c)M�M.�6�Pf��V��!�՘�d�I=���"B�5�le��_��+������t�n;�l|'
D��1��z�a �m��Τ ����a�i�&�l
��/��j��y9�c$�S�m tJ|�7�P/����ԤX����tTG/�?5�!(@G����.�a�W��Ot+�:�r[U.�b�vZX���0��<��~��uk���~�J&~� �e��0��M��sUm�LM�-̪9�s���~>�!Ϸ�c)��,�a�r���2�G� kL�`�QQ�oZ���Ч���:{�X���!=�)j�F�N{
�ԯ�jD����;��m�����V�ѡ�ի���J7�5$CBZ�^�<,E<���{��\j]�X�@s-=U��y�\*������3:��jO80���K�D0;��8�Z�}g�f�;�&�������۠c�0��cD�K�h' ��;0bw�fJ�~ý�(�#���QI���7ď�,X�aT��qf�%�.��ݼ8��i*����y3��ZO5��W�!2�/���v���'r�(��f�~}0�3���旗
EܰT�y{O�m�m��/��N\�jl����n�G8i�G�g[�����J=�XC�q��[h�q��C�!�hy�p�(��~b�ȋa8��.��5Z�=��H�8�R�=��ه��1�խp�#�˿���ie�k	mt���ĳ�e8BA����Us�V]� ���U7�&l�����u�0�Up��Ӛ�Dc)�,5*�_�[�����9�ʿ8�L#�Km��]T�������6E˶��+�o6wv6�ct���&kW�"�3�sk�<2��i��"Huѽk�rH���Ѩ͙I�w}�FhA}����7����G��2��gUS��1��b�"j�*��{O��4�9n�Z������Ջ�8���_���w-�	��	1��o�[��]͵l'�F[G @{y�t�O�l�;�`ob=�D����6�%%uA��O�XS�tI���0u9k�C����&0�m|�єԔ�rɸ�	*��mHG��!�Z�K����J���Op;��GS�0�{����v�)FV+����G9�@�u`�����Ud/���Ea����.�lY��6�c�T�^~�R���"Z��r/xd���ts�ko~@����D�\�0�k�Q-|6����.�#�����cZNd �KY��_�a�pއV\�aH��Iw!�O��$<��9t.�{�	�{iRQ�D�+�1�o4eM��ӓ�G9`���
�2��e�h�{���u���w�K��.!���E��g���7T7R:�$�3��l.gB��J�ĩ35��!xojt4�;����\��g�S���f��͚��}Ikp	[ˍ�wB'?�)A@�O�Lq�(ۄ�n)���#כ�tB�tx�T'oLl���?oA��[�2�O��_���ټ*`����:˃�F˧�I1^(%�@P�ý���������NXJİ���W$�vjx^�6��Vh�K3��F8W!�'�N?�("r��R�(g�M��#�&�`�1����$v0�3)b�AL��̏l�l7r��Vр2;3���g�(��hr���'S�{	E���cf�y[Vk�r�)���Iw�e�rГE��x��|r��&5�Y-[�u`�_�Y�(���f���&�G��|�
q�o�i�ppTL`�=�:�����4��k��ٲv9���t]S�y�s���'�t!3���W�ji��S�G���>%����3||�H�V�hB�h�*�]=�FtT�j����l�V��L�T���R���f*�}����#�8���-�o��7Q\=���ɱV9;)1��fL���N�O�o�P�:�=�!h�|�89��=s_�|+DVM���X�����d���Z�e������J�C��5ԣ�]���{�m/��;���.�zV��`��q껦�)��-:����۶����sX�EWc������4(�J��IjN���)�u��;x����>Z�����p���!|�����Y�U��`Ǌm@��i�1������:�Ov�*�ߟ\i�ݙxn����5��ʆV$p~פ2;�Y��r��Z3{c�`Sy�U�3}�Wo��:H�O~)�ð*�V���*�^�]q��+ð(?ւ������T��:?��c$C�roH���0|g��i*��9h*����x�=�Q=��� �`h��t�E��y��]��Wi�����[V-&�,N�b��j��*�Z��Q��ˡ�X&WH{�O�i|Z5oz'��
]+��f���������:1�O������M��^ˆHQ�춣/� �R��q�I�c�bи�"�v�}Ӣ��>
g�ki��WU�!Z�T�,�mwH�_iP��W��/���$��k;�,�D\���8������@�n��@1��f�F�������߷jm���i��4D�h����y��C���yl*� �c�[^K[`�Mm`%5��D��-be������K�����}�U�# �b�$$\��D�9�xy�Q��n�����OBb�����%�t���f�}{4��>�� d�%X�OtK��q�ڶ[�őpT.��e�R�Ri��Az5eK���e�k�@�\[�3�8=l����L�����-�@,����zQ�3C�0G��fj�=�8�cV_q㶗g�ؖ�L-ڌ�{by���'C]<��h[!�h�:��6�I���6fRp�B��Ju@F�=	 ;�J>"/ow'a)$��B'F%�hѳȢ��ⷠ��De�zc��m�_n	�Sn�&J�M����]��b��u'����j� b�.���@u��	�f]�TH'(��ź1�	
�ck��O^����/m�5kY��Z��I[�=s�d7������[ܟ���TI�>p<B����6}zq!+�2r�˻f?̌��Y="�0�M�LG ��j�&�+D��L�|Ӑ�{	�U�x���h�n��߈�X$3����b�< �kG.�4�������Ed,�'
X�75�En3|qMH�!�D�k�Bɵc�6t�6K��{��	�,so���0P���L�<��S�]BD�f ��3 �uOcջ�H�4�/U����h��e�K���j7"���B��Bֱ8xr�mk�� �i<�4��U�'�ސ;0�V����+��V�*�ߝbT���+��Vv�H�X�9��"T=B9�*J>o��ҥ�pȺ��l���@-;�-4��O�� l8�jg$��ny��ޙ��bn�gNB��Zu�K!R*'�l�b�܊���>guZ+nY����P�UVy�)��2���x��h�g@�;ىF�0�x^!~�䈂��I��P;�L�n Zg��t��3ۮb%�0F�|�Ԙ�r�u����ɹ��±R������3i]	D�(�Y�m4�<im����o���D��$P�ı=Y�����!�3!�}�Q���U�7H��yV��~����z~n���I�mW��j~��uW��,�ڳ�h��󪢦��[HH%�"q�i�����PaMѝQ������Q��|�,�<�*FD,6b;�Q�k���2��E�YO����?�����A��7�o*�e�QU��T�(���j�-k�����6�`�`1�,{{��@/��#i��Y��Az��?�F@�ʒ�Q��iK���LzX���Kt���NO�J��"O�д���p�b���Ĺ�c����Xm�}�����X8|�ͨXhf�V|��V�i;��0<�j�٬$G�n}z7���z�&�W/�-�˅�@E�زd-�h�h���|�t��RI<V�B��@/��}�1�?�͊2e�RZ�B�8�໛C����ÎzI�ţ����0/Òlկ��a��$�]+�����������=��n@ON��"#�"JV�{ M[m+�#Z� TF5 Vq���5(UW?jt��sG�i7ȖF4p���\�:�i�/���4�PuG�a#x���X<��~�:T9:h,/o
��D1	u���[t�fej��o;.OFK�,=�Ɛ�)#P7~���Ygu|Lx��D����B�fZˍ.�1��vX����o]���z�:r{f����Q��dF�Օ�K��	e�j~��H,�g���\�n�|�;��+�	��`�ô�@U���|~&�ԋP$�̟z�����L��Cw;G~��|2�|��B�o�/}:�6�>I�!E47����m�lbK�E\��D���Si�X֤�W�nq�#M��|����J�h@��
�J�T�q1��N�	l�����I5Ja+g%��}�Y?K'��0qD����>5e��p΂����0���:-�l����r�7��!�m9�D ����|j��뺸X&{���J]�Š��!�����:ymi1-�U7����6g���MD�RrOr@��\;֮!�� �ՠ����PsX�߼3�M�E���x\���Ἅ\��uH=�%'Bo�t��:�y���J]0�? S.t�>d �_����,z�y������[
�aP���8U8��笱U(u�u�E&��/�=W�`�'%3��0�c�ÙPY�����۶�ѵSf'��I�nYޠlnqs�
����	����S8'���l�}�K�r ��O����	�=�f�N�]!N���9���-,�a*�q8���G�UDJjs�4�N��:N�Xv��x��g�̀$����4��i���!]ܒ8뤅~�{�����)@�<�h��:G�¿��b}=�8�5��[^�<݄�[�z�"���Υ��Q���� ڐ|��ݽ�����X���� ��B	�5�㉯"ɘ�яx?�������1+��xqxA3����cF�&�Hn��asZl%�$#�o+���[�e��_�ݹ�����5�Oi�	vx�"�����]P�L��<1�NV��!�m�߀�����g�$��ԇа��ؾ���%�g��£ǉl�SgO�l2������A�S�'c`	9��Hk��N�B����2�_�܃BF���g�F��u���X�i�>�,��d� �'%K��G~}�ߤ�e&M�<�y��L`��T��P�xPv�st! �?M����P�P��}���n��G��@(�^�ɢ�'�>nT��6�{�a�An�X�����hskB���&g�,���F��Hs�0�Ld]%H~�6�4/���p����6m���}s�����%����8�N�eY�M��qb�w@�����@��$�=�`��|Lh���-��haE�m�"`yz��A���n{s���4��6��u*LAl.�/��52�K����A���۝�P���BW�ɑ>P-{���b� ��`��������T�cEy����tޣ�q��|=��������+p���ٺ_��p