��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P��v�"<ߞ��&'��k%P碶�R�ӣ�sĞ������FY&{R�edo�Mml��t���C$�i�h�v�����A�JG�
��w+���w��_3�&��Rw6��*9\%�';�٣E�a��l��1��`U(Β<��'�^�O��KC��bP���٠���RН�m��+�4Z�3�&����sFp��&�0��0Y�'-��pw
� �6R=#f�M���OB��QW���QAu�U�`�22Ǚ'�w-���6�Jt/��j�|~@ԅf{�h��P����Qi�ڼ�83�_�F�
&�Bͬk�Nr�EH�V�%���@��X9T����:ϱt*���-[F������u�f��A;�������F�O��nXsF��L������%#u�*����*�5FG(m��et 2�OA+�9�Tɍp�&��$�?
�/��T��2p?g��~�c6������Xe��Y�ܹ�!��-^��KP ���c��:�S��Ǟ�
�fl�z��
F�1k��z����B9>oH��Q�b9�K�
�:]̷�d�]V�
�����'�Y�B"��*@��zU������0C�����-N-��hJ��s��/�m��_�Ȃ�A��E��Q~�)>21��{4��Q�
�G}��q!����t�: ��@�n.~Yш=>0�A�̃�[�G��bi��� _}D�/Y���΁�\�u�3�H-�����3)�*�,y��DQ�����.�!��e��e�����ܩ�]��EE�B��#���S6�6���QfK=6�PFF ����+�?�ic�Z"��G����3 v�^�'R|;#Р8��Z�9�%�q�|M�d���J:Ү��?P�����������K��"�4��V������q|���'��_�B�E|-����fox�ݍJF���,"3Bz�_c&X`2�q��Z�_����^����5�H�]5�.�&���`w:�փ�I��7�rT*�5_A�������3ݽa^4k	4���%�<5�s�PB�	-��_@ژly,̓��rB���D�������ⓞJ3�!�nm�q/�J��k_�Ł�S*�"�I�K��|\~(��N5^ks��Rn
�z�g�f�I�j�wݍ�j�SE%d1�G�v�����=f������
��n�;%w�z>�(��qdֶg�- �G�5G���ѾOe�Z���MmW�jC;U9\I��L� �'_�r	Z���x��aŃ�%�p׿R�A�A��ږuP�v��L�Y�Q66��[�(	Y����z*�D��V���)�u�<r���������'�[,I�~�����Uι�=s҂"�(B���e%23(�na'�7�=�LH	�6~��(�.�	_*q��@?��z�q�$\���}d�:�1��M����^4ɂ�������M�Rp�jiVѦ��"Β���F�F%�D¥,�gx��.���Q�<�`�@��D���4U*��Us	o]����a���S9�"��~g�O���U$��ɚ�1ߍ
S��U�%ǒA:;kO���+گ�+�
�L��#�Q���x{������x_z�,|���צ��	� �K�w8N��"s�4i%�bcw�분�8A�M�!9���Vi�m�6�E�7c���}t��]��5mw��?�*�;|��#�N3�oK��^>{�A�ޭ��?��z*�Y�3
Qz�����\��Dt�;�I[1�4H�n`%FO�Ip��N�\�`gu�Zd.�cF�4^���1M���|��=m����e��^��b:�����"���6s��u�B�Ұ�)����7B������F���s�6-j6j?��庮���Cj��*�����<����~j�1�hC���n�+l��r�f6{���Wf�{���N����&�ǩ�Q�䏃���9H��(P+�
D�Z68�H�V�t�ryf�كzT*�rޙf��ԹԻ>Se�>������ⳛwp>��
�69�X���NѮ�^�;c��{�
,,���0�y1���������S��?�]�iŝc�� =�ɭ��?S$٘�
������k�x7u�h����-�OF~�M2]誦�E��ҁ��Xe!s\jB�/߇��\��
�q~�R��k�R�A�����n,o|��Zo���SpN�/&�X��"�t^���@3�ݭ�
������ev����r�Ck��S��!�HLU���>�=RnD؎�7j�|��'j	�O�w\n�}ČD�'U����և #v�0�902nb���$�0���.kz�.7�Y�� �����T[�_ M�o�-�ཱི�֚A��N���*s�2���86����+�S�B��(rj7��?�`�^���Y�H6������B`����7��	�L�&ô*��%Oa?I�Q�^�/���~q�C����E
F���٪��D�t8��3|�p|E���T"�U�]���D���(S�u�������v˦<Q�������,q{y�4� �y�в��4��������K��CY�Ւ*�y�{�ߵˢtF��P�v��E\����v6i��޼7 ����l4�R~���\�mL��U@��b�&����0��fTN�37Yp�l���a���Q�Α�@�Q����[���g��c,�4�Ң�u�	y�MImvq��s���^L�FYM~����d6dfb(Ös�a�6�AK(��涀ȹ�fQ_j��&b�u�_aZ���7[��ity	n>lU�:r�5��)=�(#A�[܁�ղtnP�f��O:=[�Rc��dQL XE4�s_�'4������P`8�L�Y��珜sԧwya�n�Zg��G|�2[�t,��SA8�4^�
2n���k��Y~F)Gv�y~�H��vf�� �� �	D�`�?�^����)�|嵓D0aP:绫�e�-���Qzp�\��m�v2Cf���p.�s�X�ӣQ�!%�����'�0(d��wའ�j���ޯ�O�����5������@��Z+ TE�WA��R���+y��i�[�I�b�q`j�}} u_��+�S~�o0����}$Ik�z�@g��  �"� *Qu����ؕ��7�-E�g5�L��W�j���[e���t��[-0������(��H��s�ō����{3$8X(� �r>��rǰ�tZT\C��BpM���R������e�����(8B�����c���ߑ��͏2ҟt�9��?�yƩ<�Nj骮�X�G�Y>Y|���T�f߰15�c�p�M;6�S�/|�v	�Ӂ3(��W�����U�z���rv�i���?��$�Pfs^���ĐAtd�M��	%���N$l1���f��ܥ
��y;���иÐ���-)�_�fE'_� Gͱx��;4U� �9����M�QB���`�,R����,
AJC�E7#;�s�ҫ�5�����a���T�}�M����(5�ϥ���Kà��=�����[>�g�;@�<f�*��&].�%�1�+"_��2��سA��(�@,htf�Uي�\�݌�E.��b�I�&?�솾�5��8�	_�����Q���s�����*G�~�]��3%���igq��������z�j]w�CxI��?L�I�I�=�Y=n�S+H�MfR\�}m�	�Ş���f�(n�ϻ���3��<:h�pG;�0e�U�9��:�1�J*fݿi;��˞Z�'O�b��D9\oݴS�����@�B���]�{�J%�6Y$��&tk���*X�����5L�-�҉.[d;�S��y� L���O����Gsg�5@�n�.���g>��!ch�`�رR��#D]�j𶦥Q8A/4�3q��ۙ��-���8e������}�G��Zv�49�"䞂����
�S��^yJ�2>�Cl5D��y\o���g�̰R��d�ģ�$��^���].�-���q�!�w@]M�=u�W��s��d�t��H��瞁n��]q	0�h0�3���JW�:k���A�S�� �eٵ�N�ޅ�ڮN�N�J��!�H�%�<���1���=�t����Nѣ����:�6mH�uMc�:d�B��g�pK{Y�᧕jhA@��Ҧ�Ti�Ob~^�!���Z��Tw
*rUw:]�~��*��#���и����TO g{	)9+�1r�� l���ë/���XH�SO?O��MC��&���
?ߪ�*�o�_2^f5�	�a^!��B���#�Bb�.�1e�&`����!���Շ�D��v&J-��q�vck�?L�÷�>���9Y�rU-�b����TΑ�R��ǫY!Ľm�j058-X ��|����>,�_�V��D��-���!��Ow�>m,�E0���%>%�;}��V�*�C~�6d��%�2�4L�3O���Œ� �� <
��܍�l47Z�W�����ƫ��A�Q����#����1�̿V@h�������f)�K(�'��('���jW�����-ݏ<s���7c���|��y���b:��f(X���Dܿ��|smAt����)����S�!*<��g�foLO@'<՚��r���n�k����Ռ)�>�?0�	
�2�Kz��M��F��2Vz��h�8 ��o/:x�i��P���>�ΈJ�%$�ʑ�Ut㕇x\1�=iЃA	�
!��v��T�4<xØ>HU�d�2\��i%q���||�z�R�;.�@��7"Kn�L~jW�8�>�Q�lv���>HW����И,�܄�NQ�N�Y=jo�rtўD֝](�������uN'(�vh��q���2M��=g�]i�.:�Y��?W}���d�Β<�:�(�����^?$9�v�R,Zߒ|�,'w�G6�X8*DPг�\O�rt�I2eZ" �ٺ���ᰦ�9b$��'����\�O�_)��B�f�I�H�F&kIF%P=t1��=�����b�pHa>5�)�?��&�e>'V�;�GOa��zS�G7�rV�C�Z�|�vVpx}�;���v&응�Q����&q�I��C@�_�ѱ3���*F2����2#8�p*}&�&\���zJ�]Ȏ.��Mq~ؑq�3��j&n���d�~�l��HIt �9�7M�mi�m7�Oqa24�"��\$��v�?� �W=6�q*ý�	�E;�q�JQ�
q[��0YW��v�v��/QOvg'�:�iz�u�:eO?�K��<���@��n�֭dN'�? _��Os�E^$���;��,D6�3!���������)x�OC�R5ډn8�::﫟�=p�{�x�� ��t[�jK'��lm����41���Dp�&��(PgF�w���n��k��;�*}�Ͱ|[)�R5ݸ�!��&k���q�]6�k��U"��z�aJW�M��ݠ��s�z&�>Y,8.Q�>h0�p	/�9����-o�V����������ҧDJI���ʈ1,$\��I
�L��%L$�q&���;MǱ�!�Ύ�ȥ/qe�c���N�w@�ㄾ��,!�����A�8[Z�M�|���j�����ǘeN70or7��o����%���>Ce�2���«�ōOʗ�růM`1d�#i_[�����4ۏE��̬:��r��>��:K0E����yGFR:~Y�����#�ܠ�P�}댹����?RuH��oÔ���6� t����#Q��)��z#7;bKJ,u	!�+U�5˺O�U��'�6T8c|Q63wS�{%1��B���^��y��e��,�p[���+SO���9}�^_����A�U�XL�)`��#	k�#�jj�9[�D��<^�	�sӧ���U�������1/�5��H�H�l������Ҧ� �(�,�9k�|���-Z(,��Af�GUm?�~�ο�٦�7�n���^��aJ����ÞFP߳��v�fx��E7��nx��.%%i<���f��������8����^�z6�C�2��{�E/`����N�ɌW�~�/���p�T��j�^S�������ڵ�Ǉ�[N�uV�E�,i]�Y��hL�O��,\ꡪ�CEw�Ps�dN�����_���k3-�Y"4��޼z�w'l�)�]���u�ϫe�o��Y�=U�t/�i���Er��0!�)�N�<�c͹�;��_�!��y��a� ��V��վa���c�l�N}�b�?�sr`�� (R��?��Nx�h��&���z\ N)�zȶm1��[��k�U��8�7o�Π�_M�LN�b��68�wļ��:tWu�a�^�ռw��Z}#x�v��{[�gw�W���b��w*��(r���:���� T��F�>�qœ�FnO7����P0�Ō�_B,%�_[s��KFk���ع
�Ncv�KV�AךZ���5	��^.8=�6��*��:����r�`Jݭ��Oa�O\�~/���R�y9����z]� �X`E*>�"V�GQ�|���Q"ln�S �	E��\�I+_�< Y�kz��M"���؀��`8�*>F��W��_�x˙5Ӎ�6��B��>� �@pmh�x���AR��w�Vb�e'D6�o�ۺ��67���*k�SrM���ls�(Ph=zR�e�;!r�)��_e��X�T6���ˣ���/�8S�B@���:1su�p�#����8��
M.��/�ﯭa�K���ʦQ*�pHֿ�;D�Yaf'��G�"G���]�)H�3׃�Q��cJMS�Ճ���F[&B�\j��X*��Y��F�X>���7Ypda����ʮ������}f7����H#>��͝���(0	��m���Gir�t3x>�!6Bf8L���z�O��<��[���'L�$;����'���V�(��EC=�
��3�z!P����Hl��Da>٧s�e��XP���\b��E��a��rt5O��AI�}@T-ZhoK2|�����?�����po����(��=�ctW&8�.\�N^��qe���X�s�0=��I^��t(H�+��)^�u�&�a��	tl�p� o5��.3�S�koLQ������2��kaaQ�]0q�m_��7��>����"3x.�y��:���f,��IgҎ�.��H�]��c2hL�I&;�D��7��L��pc7��i�����8[�û��v#����C�wK�%�_vZ��q���o2���]���Nڿ\�m�HF|�i��Y!Pj������b"P[��� Y��&z�Y�����*��f�J�<!
�>���M���7\<����qP!��$�r@�h��m���Os0��j��OD+������ 9����u�� �Y�f�vS��;�2"�P�z$�`~� �kw0G3{�s�N��j�����zI�� ,lf���Tӎ��S�'��FX��5����Ӻ��z�LЕ�'���ףR:�x_U^`��R�q�xs�Eq�QJy�p!��h�q&Cx�|ב���$�����Rm�%�1�$ ��Ռ|��y���1�=��_��͒!��/]G��6:D�_��y܂�A�٧����^ޗyR7
H(6 �D�SG��Ǳ����N���ѯ@��"~�'RE�%����,�>@�?�q�\ s�����m��h���n�/��s�so�@p}�J4����D|{���+V���
,$ÿ@�fcِ�x��΍a戭d�a��p�{'�m��
�>t<V8�Ȯ��/r�/��㵴����?�G^���3����?��e��p�_cR�Q�5��:�	Z�[�{I�H��B)���W��Ը"�t����,E��Y�xL��*ɼ}o�
�,��j�z�S/ٔ�#�c�q���;�а�T)+C�F����@�m�;�W����~����|m�d
Q����)�>��,zc�㯐H
�P�Q����8��Z���9b�W��UV�j���D��>�<�Gf�r�w$a޹w�Qt@)��#K\�\��&^�l �Ǖ|��$t[{�4)M0.�5��	�|I��2�516ԛ�r�;�"�Ã��������Z��s� i�5�_�k��g{�|kǫ�J���z�N��æ��pX)�!�K��ꕹ���C���)w�	���� ;RJn�����U���k�J�n�u��#-��W���0�y�|��m36(��EX_0NBJ��Zˈ���Qs� 8�*�Bk:q-k?��k\c,���ayAu�;ʭ�H�yA������*�։�� S�#� �lR��n�w�?���`�7��&
�U�iT3�Ză��e��m�O!��?[�<}���O)кB7�LK�d��Vz?Y��m�����v� ܙ�v���m�f�!7�Q��&�ˋߦdMxS��0��ZuRnϼB�U�(*.�
�����.��3�q�a����
�?��n�=:ς����K��<YB �ƲSXK�7 V�%E��y����Ɨ�Ybz��s�7-������~�O�i�G��/�F�O�
.]$��s�:��Y& �y���#��o*�j��T����㤹m�?F�M=Q� ��Đ�ϘM��+>,!��z4}!�@_ݹ��p����W�-b�V��j{�x&�?�K'i�A�Z\o����]1�YA~��8��Dó�o��؆�*�ptl��.�_6��MZ���8���� ?���7����p%)3M�S7h�� G�8Gw)����!E!D-�H/""����cj<O$p����2T��Koß��;�t��ѼmK�[|�S�ı��	�c\c_���V�oL�ݢ��0����=z9���eښd٨��Es0���;�^�p6sm�M�56����Z���Sʍb�V����G&�E_-��(�6}��a�!�	�0���h�c��'`�p�Z�cc���Jm�J�y�v��t�iU)fhN�X�\4�2o0���V�ͽ����P]�]��NDr��I�X6
��
H���KZ����Wl�x�d@�[Ź��4��Y�h�7�.c��Q�Z�}�Y�`t�>B�8 �b�d��#�Ps-��vs��k�8p��� H;>��p�`}�n�`��r���ɇ��4&�9�50Z�Iݛv�Wъ��Y����