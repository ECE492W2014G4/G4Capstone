��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��/��Q�w���a5P��B�~�/�'̙���S{���^�qѝz��'�hřD~dVr�F�!5�=��[�\�bYzy��d�(5���*���D#����=�6�c�p�GCE�N��+�xh�Eaa�Ƭ�z�5>��>s(�oƤx]C��F�i�TϚo�2���E���W�۠N	Rw��#fa�E����ǁ'�iM�$r����?�W���aݒ�3��L��'�ފ�q��p��FU����vJ�k�~���l���wFpe [�29��Zq���)Rq�� �CPu�)�;��/�V�2��'cu�*�Q��펊(�Ľ�|�3ڟ����<�0�D�>,�n�i�63�'�҂M�N9��������8��x�����k(��v��V�>9ʌ��h���^4��?��7��_�P'Jf5����/N����(C0�N}rpg����@�a8���*c��#�`�/�����<��CÓ�:�It�"���� z`)G�F&�'�A����M)W�]�3 4���-�	<ڥ3�`���^o��y��r�X"���"ķ��U�3��&Z���v$�3��K����V�A2�����1m�
������P���8P�}���� ��p�
d��N��Z����c
��a���W�5!g�D�\��.��f�up�K�)�,C�[<�Y_���k̳?� 6����
��=�3��:]��5� l����l��� <��7�C�U���T�'����R`�W^��$i��j��3�H񽼎�ȅ�l���l���ju'�
2&X���#���#�"VӓQ�u���m~u&���e�G���%����7I!��2
��~��BW������ɤx�1��=�'ž��+�<!��(�ح�Nh���3Q����Y�������
��;�_���|P5��5C�=��j0Ə���h$�8J�Zmsf��ԟ�x��s7{�h��mf�t��Wc�s�K��/�*�� D0�i)9��Ÿ��{��3����n␤/J����ŇV�ZfR�IRZsl����	���X�إ�Y�'v�l)s>��2F�VL�	����&��V�ʚ��6f�%g�P �߶�]��T����sEw~\�)�L�^ ]��O@籛;��҄�:N�ԎX���$�����q�m�~��7�4�Y��kG�qJ�>�8�eT�++�>�|jIK�ҽ�l1&q�n��}pԣ.�����o��K��C�K/��!���L�ޞ1�9�̼�RĲ�G����>@�D��Իp�5�K�Ӟgv�7�T���2o��"�V�,Αd?�?�e��_�6��#�]V@D��Z�\G]���B=+x�֎۝Aa���- 8i��T�N:��f�+͑|I�Ⴁ�r��V�i��P�2�Rj�,}�B�U��xn?Ń�h#�0�s�$n1��)�CZ��\�Z��fDV��7��e?F�͙��(��系_��G~�m�7#���O������ �歉�&�DK�7�LB�%[{&�ۻ�X5'��da���L���͞��R栈	�]�</\��C�V�ќ���z��n��t�\ν���f��rn��b�L��
B|w��9��碲�[��⻷�\_�H�pS����AZ�/`}�$2_im�k[�8bP(2cyg���{ϣ�}�2K(h�؄	Rƻ��;ƿ���;J4�y�S��W����bv��v�`;Z_Yq4'G&QfbY����Q��.8����7YvH�H&�ҭ�=%o��)��=�ɲ�iv.m���l4�߻�� c�0��bQ�!5�0Ͻ9���UY�>=|u`��g��򙭪���	c0~`8���&ָ��`��*�"Ѝ�8z�(oL��⭲a������iF�0��P��<�������w�Y�j�/�"h���jzu�u�|ʟt;!0{B��
�{.�"~���J��3��h��(Y�Ts�'�%�Mw1f�¿o�#��O�ئ&}��4F��ה�N*��w�����t�~��p�%C�����5���i %Eب���qSB֋\Y�"h��g
0݉Y�קA��;�X��X5�	ll2,4�_nT��^�gk�̤�Q����ߣ>I��L۬�v眛[@W�y���:(�g�\�:&g	 4��ƊV�$�������K5u��pU�������G�\�����n�yٰ\q#�� Xٿ���T�ۆ�{�3�u̸d+��>�/=s�F\�
� `ȴ���4E�PD��K�[�Z4�Ih�g�hT��F���U�or6���F}�����S�P�	�ͯ��ϡv[�6��>jO	˧cC`fD�8ao,���8���/f{K1G �T�6�aYE�O�1�2��q��mJ/�!��1��d���ٞ2)/�v��'�a�ϵ"9zA9�5fa��Y���K}k����6�a�)>�)�:�w���8��O;���<�]�����N����	wn�n���5��9:����Z>m=�?��jD�#i[���y(>n����'�{#�>C�T�\ss���E�w����ɇ'*^V:xDq�hk�4�%sA@J?Baz���N�;v,B���ּ�I�����������rP�,E�~��\�n�E��3�I����W�(�cneǖs���=��o ��¼�\�:����g��^P~a�>p�d��j>2��"]�iZ�oKY�=Vӧ_ָ��F���q �x��G�	E�wj)��pԋ�%�u/d� �mAᖒpr�0Xz�ĭ����}L���L]QH�u`���u
�e��{*VUhR���,v�_z	��ť�9e�| �Z}��"�H,�MN���Ly��|V���T�&>�ҏ|�xBqh��Å[�g������3c�޴6�A(���'��a\է�ψ�������`�^���9F�7��-�}Q���
��1�W[/�J�(V����0y�l�
�b�Um�C_��׍W慲OI�u�f�\��ڏ�G��#I����"�DL����!��\�SQ���CdDh������l�yQ�^���W!����]ڃ	Ӓ	���Sm�}�Eɒ��B��"6�*����"�Ȍ����l�e��[�3����@�|��>Z�rD��g>G&��;�9 �-�gɲ&����U�h�{��FT�(����L�j^;�0fX�
h�} p39!	@|֓�ek��6jK`7���lg>�^	(�EiI@
�㡰�s����A2@�b���B�
���y�=�v���1`Ef�c����q��z�`)5�'jUq�;���C����tG�*U�Fg�@W�L��E���C9�֤���kHP�E$ʎˏ��G1�� "q��}�_�/R�~��iR�*r6�pE�V��]��Ԕ���S*�l���`�8(hJɇ���5����5���]P �hۅ�����Q�Ҙ+g����ROg8��N��Tz�g<��7���;E�S,�t>�ϑ\��҃�r�wģj3�j3�].��W }����h��۶���y�0#h�ߞ� &�����i�z�խ�9�^��L�4��\4j��PK�L��mq�c��?�[���ND?1���QS��#G����Pp��+z��领��G�(�a9���؊9 �-2&f���JAYJ\�P̨Օ ��o����2~s�|ݨ  fǃ1ud��!�C�h`N ql�i�Zh�b��F�W�-����tm5�;ڋ�}:[�R���ǎ�=���)��%Q,0�T���<O8"��(Ԥ�*
F�������5�4����etϋC-�vEv�(',��c��p� oݏ&6��� �i���eBzim�>G����>��`�	N�P!��~i�bu|�?*��jG����$�r������V�Q=
��C����K�햴���񨌦i	���_�`m�I7��HWu�8.X��q�N��-���8�)�ֲۻ������-�l�s|���Z<��F���<<�"�{���K{p+������C[��tY��Iq~�Z�=X���`4�~��Nf���p��9b�Y��5�7ى��-�8��^!�ï`?hi;�툞4�>�~l\��v�[PC��Ol{R�E��( �l��	��o�����V�h"����]�����b�"�!�%�A�H���)ÈB�_����BU̧�y�>A6�Ý�H���v1܁���&��{e�����4��sU۬卶5��6MX�Q��>U"��us��*�H�-�|=a>�۰E�9���=�����I���`�(�M��f�B*��b� �������l��9�iz�d���Hq`ʓy�"1�3S8������%�$�����t[������;����O{/�Ro��,F~i}�m�Ȥ�
p[��M��Rb���}}D���O��!����L~�Nv�!~2���wH[N]4�LtYٲ��\6�>T�[�0&�s>��ջ�z�Y�'F�y���D�Rƚ��u"�GǎUA��s�*����R���a�K$��X��V���p8�$�-��At�B����Qo���AZ������yn�)�3zHH��_%7�u�.�!m F���o΍�5+�[y �ǫX{~��)���46��s��u-kGw8ӎZR��@'����U�s�Ҟ���P����?v�
�!�h�!K��H*8%��.����1Goz�bO16�OC�T�q�¨.C<�f`��9pa:��4�� K�3n'��v��Pn�����A��v6�f����X.{覷_5����4%3/j��z`=ޟ�eGL��3]�c,���k�����w����4Β?�$��#��6l̘!2K�%�y5��/���yRgԎ�}tBȇl�^�԰�2t̤ZC���C7o�N&N��z�Q�{��(�;�bP#�����V�E�h��9�iN��ý���w�����<���(F�nZ 2�Y���J�@��GK A=\D����]G��<��v�{��Ο4�A&�^վc�ʺƵV����N28���QaCQ	�_5x�J��Q�r���Ѡx��c��"��t��]d�)+�4t�!�"?y-��Cs�Ҵ����x0��
+RB���\��^�0`vb�Y�q���*��`����M�����`�}]l���j9��@2�rH�T:�Q�WMu��>��cC��d^Ţ2'y����3}�T�N�l��iH��'�M���� aP��L��)y	OT���v`�Q]=�|s�����0�Z�Ho'�ؼ�����ϸº�4K*����{1�o��j�^����(����O@#Z�d ����X�+S�`� �g�yɘ���U���t>�������R�jK{��n�O	��:�Ө"�f?oB��p��άX����Z�b�������JKGz�\�H���X3P���� e,�d���w�Մl�e�J�%��s��2�-0u�(q��CwF�ʏ h�������
`�0�� \�F��c� �j7�y���q�D�����)|7��1����n�]~��5X���d-w��\�	���O"��e���(dcU�ik�V���J$4������,\�@����n��b��cW�����}$H� �:����K�?\`�v����$}e}k�kG~b���ڶ��D5J'�n�������'-�a֒#Q3���Y�2�d�7��w�rc�X)H�T���V{懫���c��Y9%Hlq��`L̙~Y��KQ��yY*Z������5	�?�>�!㪂�A`����|��koKU�^9��2ҋ`qrj�£y�v5eԺq�.X�}��aV��>�`�2���	��8T$�VE#zs���\�B�-�]'�2t���O?�9o`����f����v�ۄo3r��9�7*��r�RM̂�������	��X���@��e��я�Ĳ�M@im�g)Un�c�dd:A��C�|C�T��'�a�+]O�`��٠��A�8�s=n߄-'BK��dq��̈́;=�K8������ެ#�g��	���>L��uQ�芏�'� 0�Jķ��:Ȉ�M���P݆�5�d�{6U�_&òךmM�Ǡ�"Q(��~'���O���X,GSO���noЩX�y��#f ~��:�TL����G��A�|��p�[>�KRt�9�����̘�?��7/��H�q	>[=��;+D��jz����w��6�uq��e���s@����"����o��°RI�@e�V�q��E��n�.�QƕD�s*f�^K�����L2�}��t%n���p���'��L��5�`я��T�;���]�!��4p鐯��[�
E���G�_�XO���x}�.`�i�3���o�c�?Lǎ ��w���J�O��\j�}��b?M���HQIߨ���~I��ȡh�79�[�j-*�C�7�e:p�����N	C��}*n���D�]��;|;br�6O�N��&�-�R&���P`L�K��=�|��{EE^(�" {�*�B���P]�6e����G��'f;M�+��3ثy�ߗ �0�@z��Ykk.��(N(n�S%$� ��u�
���p�����S���P�_�ZVb��� ������P����Tj�ǯ:�:V %t��q�N���0a�LȬ�,\�-���y1%�1D+���W甔}:κ�X�{�ұ�~�t��3��'���P���y�D4,S����!Z��R��k@9F^>�_��]��a�xEs�bEzGEW���a(�P�`K�)���Y����-���k���V�Sl��fam�v�0/���'�
~�����>K�ɥ�w[�+��5��_��Ӝ�(��.Ԟ򰼙�"!5��4iT�[ȳ��"x|�=�D�����,C�������XfY%����-R�63EU��$����(O�tk�����ɱ��{����_����g�4��/ް��Z'�fN���r�����f�,�n)B<�R���`��.����O���(�3�%uXW�O%;m��Hѕwg�	���C>R�~-�2�W��i��*T�u��%F��piO��q�;+p������3�JuQ�ˁ+��2S�%|D،�K�4z�����jB� t�Sg6]ݷ/e�US�@ca^�[ty`���j�����S��?j]��W�?/���9(B�ڏh�r�w�������侄(��\��R%�۱�<��TM���I8Z_m2������Լt]�	����<W���(�-�F���L{�d#x���+\so�yg� �!a6�<�RŢ�Ln5������XX�ө��q�������N���R>��^��K<��	n'�����;��bV�x��ذ�כ���#YA�(=}3��Բ������@-#����	`�ڸ�"V�L;jdUHU��XW�%Ǥ�Qղ�X����]���|�B�#iܷu�`�@H��h�OO��H/4�<����n�9��3����hr��.Y�7>p��$�rx��lűF�u�1����6�=K�hmY�#b��7�8J<�����21�n���G;i�W��>W�����!<��+�N;�wyr�m��D��n %����,��1�M���I�b�y�/� �A@ZGD��8 ��%�;�:K�*�ˡ	r���?;Vm���M�O�`��$�`k��P�ͦ�M&oe���*(�ϗO��g!>��0�X�["�[A{c�~��;F���$g����X�3ޯ�$ciW��,gۍ���`��W����ev��]�`��w	=�;x a�ՄP����d��Rq��zH7����(�ɧ�T�dif��"�L�V>�Ĺ�L�	�"~��oV����a^����B���+�q1�'�?"�;8��F4bo	�Y������E��΂\\^�����o��%�"'%�2N~�Uv��'x߽�n�<u�,?Ͼ-�o?�n��g���
G>%'H*���֊c_CBL�'5�i��*�]0#t�!�ͦ�,�+>ԣnqވX��j��u��a�S��_�d�p !��HYi��0�y��@�G-v�>���gpm�˗ΎmL��Y�h��1*�����
��@xb����52���0t��f�#���u�DEy�m"b�c���������,go�^��+�<8:Ub�!�p��%��Ʌ/A{�S�m�H|��YQ�#L3��#��}���E!25%��Dm����Dx-y��/a�8#9����5�'�w�;)e�z�����^d���F˵/U�_˾M=#�v���� ��X<��v�EA���� GC"�T
C�썇�ͯ���\c&�g���DY�22(2���s�N.�/�+�fH��[ =nB�Y��<�vZLЋ�a<٢9
�|0l��-ȇp��"�;���=����mYU�S<���ϧr�Ӫ��t��LL�
�B)������y?���ēb�g���2'�(�*�e�
Fa���<������$?��=��s_p�)(\5������B_ԓ��녥���3Ѐ�����,�ݴ1X"g�D�#v`�l+���(W�?���mA^�O���5���>��I���9��{����]s���_�=V�<|Ad3@�aG"�kU*�  H�U>i��h��k�L�"��£��H0�m�ww|�؟��R�~`��%���ձ�kcD�:��WN�0�}UY{��{8�:B�-j�}#�a��3����h�WPȂ"�6� 9�� L���q���p)7!��w�r�K}:c��(��tŏI�^�> m[԰�=�iM�q�2`Z���i���<�D����w9�ײFS���n�~�m���;Rp�8�l��8�?��D[:�8��d��5�b�v���fu�)[��S��B�o�k	8w��_wH,�ݯwPMe�ߑ[N�i	��qP�8�*_�@ݎ�%o wmv�������
2� �uX�>�X�[����ǉ���r��������;��rj�W�3�L���i�D��z�QJ�w0�\q���0���ڐ$K�41���4�]���<�X�Ʉ/��Ui�:t;��*ާ"���h�u-�ۛ@`�pD�ɓ��Xp{n�Iv��+��b��z���}�7��HSE�$7��
�oA�e�:6��mh覿���@�8)(��@��5PVX(/��V���wLڥ��K���w|�i���A�~}�*��e��r0ob���1W��C&�|��o����*��у�2���F����K�d �)��������j�� t8dv&�⛷�&��Yhf�w,�Ւy�'��c��:V��Bڷ#^h�h��d���S�t���N�vv[��A���Bq��ʥ�b�I(aX�4a�6?����Lh���@�Ҳ�QtDLO ��~�?X��Xvtn������}��`耕�@hWy����>T䀀~O��23^�o$��$f�y���h�Gm�<�T̂��Tv����
&B�w�1�X.�%؇;�
�ǋ���a�P���rCV$��Kc��/a�+Z����6�M'��̓�j,��j=��{��c|-Q��Ƙ����$׀Hל��̱�u�xm��� �M�pH��{3�u�18~�꽢����d����m��N۳Q����Z����|��FჁ��׹�Y����(N��ϐ�O$�H��S��_���Y��H�OK;5�w���+�dUL|2g��uf��z5Ɏ	a����+�*,������,�x��ؙ]�;��顁u�c�!�K��B ?d�G������9K<"�,����
ח�5�+@5�����q�P˝i) �*��3z�h��Q�d
�X5��9w��^y�v#��zP��;�&U	c�#��q�ꝮD[�pt4�Ä�s���W�c�^��I�7@�K�KDU��qf�y�	�!ǁ���E2f�4b;[��Ϣ���9�}��q�z��&�ū}���`�`eK ��l4TQgE�+Vy~d~����2^�̧%a�a0�M���v�!˫�"�PQ���a���u}|qU�$�)\p�p޷�oPϝď���?���Z$�J�����_��c<.��S�{�i�^�hEvR�n���q/�d�v��8Y:'�����,��,_�T��I���|y���z�(��2���W�|;`��J�Ϧx\2�"e,bl��V ��w�蝬p�o 3^%Y|o����L�/����^Ct���|���d����E�(\�Pz3j8B�,Z]e6�����"wҠG���F��j��ĦIm&Ѕh�`��Q�|j+Z�Կ�r�箏9�|���rk��H�yg�Ħ=�����BR�Æs��	UU���;���M0��Kwu�_�RH�ܜ80���*N(�o��w���&}����LY19����#�����Y�AP�r�5f�r��X���L�#���[dB�X��9��wER�?�_���Vd��ĝy&|0�8�w"�E�\[ŒP]��Q)u6��"��&�l���(����bbN�	��+�(|���*Ů�_��&����i:��2B�T_�G�]޼G����r�q�Ѯ)�X�6����V��*wK���#<H��� �V��۞�;	�����ʧ���T�lGm^���˪j�Jcn��q�6'�\?�}��}��Š�I���#Ì��pu�O�#��)d��_~4Sv�^_����6@t٪a���sc�[�.�
xm�	��2;�fGr�����$yH��)��Y�3�3��"W�ف�4��W�wc��N*�-l��3�?e��b
;;}����C�"EV+�Z��u���������̂��ߕ�����W��R�/z�6�D����9�&�*z�~o�>���q���M>�>~���i��hp���y���9���#uf�R��KJ)lqĩ�P"�P��r��=쎼%��J�r�[`��ʧ�LG�I;�5���8�R�}�,�4�F⪇����
4�ԉ������u>`�j4"�Hy�������Ł�o�
�X��x�[��p�O�)���#J3�^*�K��|L���� Q���ya7���&��z�>�\�C���"�1�(6HT�ٮN�����_1p���9�)4F���T�q>�^J��J+9��x'���+7@J����)j� �W}�Y�޲��x���|w�e�!}�/�����ImIϼ�2dMs��5%[��] ��������������r��i;׈�
T`�R���[��<Q�$M��i��{}��\�.�q�H��>�Q����ߺ6h�te��H�ݗ��m��J_N���k����۞S�HL�7�߽͠��vYX��bRBPwZ-��m�
(;�B)��#6â�}�*E�b
����1���y� �e��<]�ʯ��L��o�A�I�xF���$����0(X�y���؟&ǉ���I������8J\��#gW��4Ĝ�u4c�E`e9ș��`l{�Dqf �+r6^�P�.��ݮ�����(k��*a�05jL����R��_]i<θ��9�`�+�S/��q�$�D�"����n��T��GF���b�j�a!W�fǀ.��3=خj"����T(�Лj��}��9ƕ�z��+��hX�Ӧ���ns���&W�sʔE,�mr��O�R�U�����v�g��"�� ��^Vw�y�ح]�����#��Hr��.�9Uz(�@�,P
�7�P�]/���{�MB�=�ގ�k��yD�5PQq&ȍ݉ˉ�`����>�%�<��0�l�Ƴ����җP��{|�4�I,��o��pL�2�eۊ��H/˒��Ќ����f(ؾT�Su���u@7���O��ߴO�.��6u���@<���a�GQn���h�K�t����.?p�G��ї�t�|�<��GU�B+���O�X5�8�y���6��< $�-�u�)n�~��7:Q� յ����� |{��,��iY��c�ܤj�HG�V����!������m�Fj�e�Q�|�I�x!�Q[$�����P@.�r%����-Ņi���xE��XKv	@���<���J��V���]��N����d�7τ��S�������Olh�_��'�Z�b��U�]s��qoU��sY�O�D�x�Q6Vml�aO�n��z���_����&�?���fĜ�2!aO��طU+Ca �
�%��C�`��@s��CQ��AO��|�8�M�p��M�|ŦL[+� h(XI�d^Ѣq=�Eq�-ռ��I�����W����/�_%^9��2|��I8���M)��w�7�@�M���7�)�HH�=[���s�7� f2!/��;p�pGP���I	k�h�]t����T���5�
^�������D���u�o,�y��L�v��Ov4����9�h"��3�z��7�����F��:P;E����bn��?�DSY�>�pcSYe�ULdy�;�]Q���NЃ�&�l�yٸZw��Z��kC�$���Ũ/`� ?�q��}n�=�#
�rč�v�hrD_��ju���Ǆ��Z)�rAva��sՌ�Mʧ���p��q���p���� �D��X|V�0�E/ҙ���O���2�*Ʈ�?�L�˨)��S�h�V%r�0o����[�̈́1���I����w�A���#���OM�A�� �sRRp��1������3��^6�,�6�D�0������-��*@b��c 4$������E��Ρ��s�*�h=�^�J"��i���7!MY��v��w=��a��m;MA�.��]'NæQ12+͠�����:%����RoܑL/��M��xyD"�����4'4zi	o�C�}u��V"�Ü�:�e��g���8��R���&؁m�ٞ|�)Ua�m8���!��Az[���J),���<�����G�
=�Xt�"���=n�))�ū�h)��+qY�K碑W�O�Z�ޠ���z����$�vD@}5�ޗ��&�l�-d>!�>^�^O�����G�)�E��ځ�k�͜�����7d���7g�#8,3�RV��,s�����?���4� �P���\���q&����̳�h��H�1Լ��2*%�<��4�ְ�-���z���w���쇂�Tg��	�I��ZA���дm/,�
�9��eM���K�E�\\��t��J��������~�C�^���cP��UR����Z�D��@��5��4#=_��S�tme^tѵ���g较{��i�z�_�:�
�����.�p� ��%A��D�X�B���\�{#gh� _W$HP�[ά8X�|~��"�=��]��H�.�s]��P��ʹ&�_����ƥ��;��;>�o-^�+/\;W��_��e��a�E�CʆgD��+�F�.\�� �ࢎ)��D/I+�`�L�B�<s�G����5N'�\�p_��?k�ӒJ0He�k��'���������O��Cz��W7n�,!��Ն�٥�ċ@4�I�n�# A��n�QO���	�I0|�^�h*��r�L����h��M�o�|�M۞��r����,�l��-�"cy��b�2�Պzu�$* ���VE�	�k+��4<r$ &�j�������}5x��Z�8Nς�ؑ$��WR��x�Z:��\���?�(�GE��c�q�h-y��8�D&�C��A�G=&�9��v����;� �~ga�>�7�]��&���+!?��v��9yq�^��@�L��ХX���e�4$�7O1�Zo�4�
y�B��$x o3|4�qE��A�R(T}#�
 Aq⾬�V�t����E=TNn;2���ͩ�"�I���*�/�ז�x�0vat�����Z��E�g�6�ʌc�*�v��U߯∊���k�<=fȭ���rFi�JI]��yu�7�$��uI�HZ?��ײ?�P%7��?��E���b�p&��l�X��_��2�/6�S��^r�n���OY����y@���w��s�B�f*�A��}-�j_�毑B��d��jB�{:>���1�������]�y(w񉦻�(�nv�N~��Id��SȒ�>.c�n������J��Bvm�Aa�O;%�������p��>	��&�Rx���3� 7�q;��!���#��g��J2������w�.�ar��R#�3u}ԫ��iZ��]��Q(Ma�,K�6�0G��fh {�Q��-�i��j젥5����e�R4��ږj�C�27�� R��jp(���)�x��[�oXT��Q��ε�]���!�>C,���V�[��h�n+���Ƹ#x��˸3ր)ڭ��¾NTr�fM�ʷ*�\�f[�9�V���{~^r�:+���~��?���4��-��i��ث������ՠn�tF�{���B��+����A�p�i��j��j��&d<6�������m�[�w.'������g6�D�wm����a�����
�*�Ll�G���Ȣ�`V��~���]!����(h
�z����vXƓ�H1�H.n�پ��q��mJ�m�b�O�a�3��V~�\qke��9lԡ4�:�D�"֖!��������ji�]��ø��/�����P>8���QS��_`� Gq��Aq��@=��s�W�u%,��;>Y�;��\tG���@L� 'R�"���3X؄< '�hwt��a� �?�o2���n5_���T
�$���(�a&q~��bCv�l�{�2������xQ�Pk�S�v��,oz�k����vb��|��m{����;�P0A�4R�Ĝ��k�\���+�:��\��Ԭ�#��Ð�T�����)IA;����eE�["�(h9�v1K�u/����7������Хe.=���p��x�K+ ��9./�
�{��%�#&�$��)7#���hC'��.dAw��Z���P9��9�_����f|}oo)A��w�JE�G��v������ݔ'rq�;��I��;dyK�ݔg�H�o�7���$D��R���ʛ�Z:F�c�"r� -��I9
�:�/[���\��I� 	U5D٘H\�"4`/��fq�M��$�7jn�z<�j�u���$O�])���7�����d�Yز�~���`d���Y׻f"cR�@Vg.W�<;�Yi���Yt|Ƶ���#��F��#M��!�~���|}W�=�=����6K����ѐ�$G�'0n�0�'O}�|%��)�2��ɕ��X���"ݿ�F�V:sNǛ��4��Odk��Z�U����R��N��y�?�h�eħ�����/ot4ƿ��W�6�{��eF��h�����.���m��#�DNЁ�~[��6��:&ly:�h\�h�g�G�����#��f��J,�@h1�8Bz�o��|IO��n���P�
�h��� 
NO��f#�����4���P;\��55i�����;ThS����r���A=���m~�,d=H-�n۞��E�� ph�#sW8����iA����S�����~����:Ce�Z��up�|B��xf�3&/��������,b\����{=pZj�`���4����9�b�b���x~�mW��C���w����Cb��&9%�v>)L�Ҡ�޻��$3�-\hl��������$��5��B�ݴi��!b	�) |Gh�HFtE� �g�O@{9w�W��+�(��0���<ڬ>�,�:�Bwy2M�
~��7�@�y�A�'��]5s�B��ǒ��6����L��	9��⋛9RZ� ��a��m&�3�Vc�
1��2�{g����h"Y���a HMX�H�{��*!7(�ks:�ݶ����]� S�bJ��zF$"�t%��#lx(�(�۴q���J1wʗ�k��p�#?�p�Z��Y���**�{�ܣ�/_yh�5D� 0�b�h~-�=]
��u _L�-�����wT~�;����6+�x�{�B�ɹ`��PK��í�\Cb�&�4�q��}ľ�ޛKe<,-SPٔ�8��I�5?�0� ��j`4,����;(�V@i*�F�X3i��_=��A8���<�x�B�V��7Y;�_��� .ש@]�q0q����0������4\�%�>�c�lq��]@�i���\��������3h��'4[��h���c��Ÿ��;�4}Y�B��u!��Y(2Z	�]�(����+i�q��t���llW__AK[=uX_�2E�@]q��ŽnтIR��G�f�(ӽ���"�C�S�<#�y	�3B�6O\B��D��;�����.7��gcC�cf���nݶ172��ܗqi�Lt�{�o����)�,>�SNp��p����'��ZVA�3M�	gPH�B��5D#�$|�2g�T�±��|E�3��Mߎ'0yȱ
(���O\��?�c��f��Af�m�/�wf7�E�ͺ��F��*��s�r7�ҧ���̙Jq���e��QPH_��&XAA�(�?r-���{�8�Z%U	��7���X>tr��^�~�n3�*>����zzlq��5�5	�֪;�w��c�Zʾ�Bܹ$Ov��,���H{��l�z�:�?Z�	�#%o���^�3����,b�����^�������o�*x��.&꛸�;�Hܬx�EWܦAlO�oJz/&qA��R�ɾ�Ld取�|l��ݢ�?�	�P�#cS�ܨ)�V��1�u�y���C55��]�&��thU�4o�Kmp7J�%�x�����;@Cjv[�i��4GL�ˁ�5�s0���,x��,r����CƓ�2a����Slc�
p��XMyמ.��Q+��y8�2<;mV4��8.�9b�v�H�._J��N�6"	2�@7
^�UH��)/8�����y�E�}՟��3*���N��V�R���޻��T�¿��n�y��vO�jC�zw�m�ʔ�k��
|����!�`�&��يo���֠���%�$���J�%E���y�e;�6x��6V��liơ�7x�i�^
9L)u����u��zu'�݋|�v�Q6$ji؞�!G�^��,���q}�EK6|�A��Q]{�X��cP��>��}�*ᮙ���V��ݤ��v6H��<��,Vu�VÓ0�̗l^7ν���嘁.�(�C{:^`��R�=�1#��G�4�H@�� HT�D�f摿��\�И&�TO����ֽ��9t��{��{6|����.=]��*�;���7MFܴ���}��y�RI�iJ��-9%J�:�Kjf^uG�_l����g���c"���A{����Rv�0M� �����e,�x.��Ty�g��Pa��m���~��{�����0���U�Q�����`m�`��	�$!�A�WJ�B����<F�����[G�/��`��+ӄ�1�<��y�Sq��j����,�*�Mp��U7�eߪ�ih8�:13��9���t��Ry��&��^��p�����c��Q�b�<J��L1|�#�<���4���a%�qz�o��USٮkP�v'3ﮱ@���BH1;�F��� ��+�'VHq�1Z?-zqSᛘ��e)&xEA(����ke�;�,i���ڀ���o��U�<���z�α��?�~ Th�h��XUV��P�/c�bI�{��<!�{�U:��_h�C���ۜo�.Yf���-��+��ʗ
����:'��>�;P Gj+'��>,͒<�z\���:q�-S��?�P{��O��
�s-=m&%#����.o�:l掾���L{�å�	��&%f��cRa���ķg{Fʲ[>|�yaF�"������df��'x�d7�?����JD5�e�O�#�_
�N����o4 I䝞�R�4��I�n[6����� h�EZ8�y�JkU����&9�]�m���	�}zLmGW�T<}(�;�B�
���[�l
���u[�OI@D��%�aݿ�;&����<��6wd T�IP:Rܩ�
����q��
�*7�w3�9����lt���&
tq̛}��C0���C*�7Bq��/G��>��ȕ��*e��
kR�����Q�
w������Qwn��n��I����zX�F򸕐
�V���u�� ��O&�y}��:�F>��rV���MkPi���`2��T��sْg������$�m��_8�0s�J��
�
�g�}�n��JH��J��Z���~��+pͿe��Y� ���>T�*l�ZA�!�ư��� -����:o��z��RL��EJ.��Z�L�f��tiP��j�?M�ڵ�!�<�;T(xh�m��35;	�k$��5@����vv#Ȏz����2A���}���;�a3���LOj"΅9/.9�~�_�wa$��?��X�T�3�������S���1b^eRf�^���b�l�m�ڋ�V��	��-xH-��⦘��#/�����{Ys���L�~��!�[�'pp���`�Юd\��Ae�ђՀK��=����z2�GDy}J;�d�k��*#~�r�x	����G��H��T�� "����YX��OT�;;;��`����[Q����$�p"���A��6s<B��Y��7�| :M��a��ʘ}`͡r��Sܠ�1��P�d[aӦ�6��Ԯ�؋v,��0q�������QO�ٟ��J�w�-6�9S5l|����T�7�7�M��O)��o;T���T�+js ��a @~���a�`/�عtDt~�3�y��%sh�/ː�*c^ X�z�mG8�l�RU+�o�Tqh��\�>|�
9�!��ƒb�҈�*,��)b\�����\C�w����%̦����EؗzUz��|�14<XA�Y�,|�}�.�0^#&�k�R�28�̼#Exf���1h������!�+*��
kf�銉��%nێ�9��H�W-��h=���Zm��9���j�AB#�H�HA/&�hr\}�mv��)�<t=ؙq'�,��?_y�����v	�2$�K0߸Te��ݛ���];���j��w�O((%� 2,V�a]�Vmbr�,�Yv�;�[a��-�1k|�)β����r����:$�3-����us.���zt5u�<�:����):��|�������9��?T��R��L�Gc&�����Gj�K��O�XO�i=ٜ�r�����P����2�vj�1����\�`}.��N#l�����裑�S���VE{ ��~ W��Q�`�'IS�O��P�i��tӆTT�0�S 0�)c`-S@���ϕ�F��/;p-��r��e[E����Cq��l��K��Z�H�V��$�,��M�D �3�["+2��,a�1�K%mq���%����Z�'	V�|�z]X�=�&x��/l�W�W�G���v)����� �K��?Mm��cTd�x��EȌʝ��E��{�{��)�7�Es�>"܆���������?}uG�i�ɑ k�9I�%���,��5���vy�s����+#����=���	�#�%a���+?��9]�J-����[�z~�
�]�v� 4�u���Wɂ6�V7���_RУ|�jsk$�vW����MDu�����m�(
ֱh=ϧ��K���W�]|�h�y�ҋ��jV"A����ƥ�_i����#��$�`�����3��U��Z;9�/X�8�V�.Rw�hĉH�Ec��}�������8F����_�?b�>����Sq���j��7}�e#J�>�,W���F�gc�6��%���r�c�	��ʆvQL�L ���������J���؅'�g�kh���F	�IZ�,Y.~ �@'�#���C��[b�N`6��;��"�y��E��_y��"�4g^G�*yg.<����S�T�D�o��0�c	?�( ׻�4;l�
�Կ�"�殠�2���Nu���M�h��j��^�� �4��nGգԗ)�y@�cU?�B��FU}en�ܖI�X���X�V�<-8��1�d���|:��p=-b��!�F�����;R-仹������XD�J-nSi6�y�	���ozӎ"��ba��4݀fA�;�g�N�&���%ěIQft2��ˉ��H&���2���x��^xwvjcL)3:L������?�WGEo]�?���>&-e�j�SgK�[����<l���Z��~c0�<�����|!2�gq����g�&T?(j�P�*X����}�<�}���@�����č����w.`��ge���˃�$�@�FC�q[����C�ܦ�E=���Ř��p2l3V�1{k�J}{t�O=�m�g�;1���N*f���pl
�OQ��_���t+rQ�J�ض�3��f�dI=60�$k��G����?�q��;X �-�q֗��y��#U��^5E��1��3=�o��
ο<HАl�������ǩٔtX0�G�4bm��''�VD&`F_��7���&���`��o�l���]�vf�����J�w���P� ��]W�Hy)�k�dJD��󒷛��w����Q����PiC�-ϦCQ���4��(�'�0�W��k�T��v�)q�h�X�Gۏ�5?� ��/̽�ڷ�bg��:ђ���T�*��&�-��!�T�WJ)��GL=R�3����h��Rh�پ�5��.n_Y�8�>�t_�0+O�kXa�'�����1�Z�F�l��B2�����E:}W��I<������N��\�V�5�"�\�ؖf7��a�!��������s��u�A-�p�d���!�2t�Eh�s#��>K�Z_$yi�v�K��J.�z�fK�������a�������!�TA��P�B{6@Ҍ)k�;�_L�n,2p\��4�oaM&C�J���t����� ���.��﬽��[W���Mfd'�����G��aW�l��O��P�3�Fz�躿���Ó� �����[��U��e�<@l�~�!�Io���ؔ+��S���R"y �ި��g��k�y�Q� ����#uVƳ�O�H�Q��s^*�ǋ(��;0sGvp��e���vr�)����`o\k��#��ȇlÕ��]��d�����I�&��޵�h�2��
��f�^PטLW�s���w3\ok���Qa�ҹ��p]3�*�MpԌ�t�`���d�|}XIO��b�DAoY�N�3ڦ����d�Kc(dķ@��&nZ���q� R���ks��4,Nl�/!2�5w#���E��AF.�UtG+9>W�K���Mu����L5���M���t��d&�X2"�fqE��8�%	[�����h����!mr������07j��v|�i�30��M=����k�%�B��HNפ�w��,�tM$xQO&zہ��
pʵW��\f���o=y�b��d�| '��d�G+��\:S3��-����J\5V����D�_>9E|@��4U�8��9��%g�����Q�
KbO��bB@{F��OE��2R�8r�t��'��ߐ�ɐ�Ru�Wy�5�R�nNVh�NS!�ԡ�3iᾸ恖��
�q�){��U�R)x�J�������{ѵ~3�y��(D�l�U�27FoC���<��iHʌQ�Ǜ�?��̽C�9e����{��K�D��-on����g�ڕ��
Vn��iQ�&��`��F.�d�N��=CUE��}�j,��g��.PD ����Wp�_��ˀ��V�S���5�Q��I;��M���m~���Ԉ۴f�\3��b2O�l�\��lK��	�缯F��u�Ϯ�(��#jd��Qdy�
�~Q�1��;c�/�U�������s�v+T �x���3�j"����("mjB R�[ө����������?����NrE�%���	} �3� B@�o��4���v���Θh`(�+�Y�[��C�tF|wȊK!��!��_�~�,�ʉ��4d\|�V�jc�Po���/�ARA)��.���R��t8��a�w6P��N8
L��&5�2+RXI	ǉ��rZ���O{?�|�Q���{��_�L^��;�б���[9�>�4�v��'�!t��*aϮWq2�O���H!v3�ئr�����d�f�^��-�B��^�)>�Vy��*Ҫڼ >x���ϟ��>Ϸ|�����W���+���ʠӍnY�N;�\�1D.�=���L�N��wJ=}��j_�XT�ݿT9��^�.R,mL�s*bb�.#R?�WY,l뼰�<����x�2���ƥ�.`M%�GE�e�7;J��
�1��]�ƒ,�b݂���Q���Y%��+;�ԨE���оV��K(	4^��tS@����q���b���.?~�b���_�=\����)���UK�T��Ʀu_pi�;�z1o������vo.�nӬz�<�S��,�()�ݽL�C��5)��g�����h����J�����S�tգ%u]"��.�0�?*�w%���sT��շ5��b�	8 �~��Ԣ���ql� -d��Ģ�.��Ӭ�sQ@89�������A�>������Q1>�h�5�)����'��t[�[�,��d��Ⳳ�8ȣ"���P��=�$��R ΃r��h�H�F�Bm:�mTV�A� H��(��D~J?�K��`��׆<��I��n�3N6e5l�=�{�@ ����O�t��߁v��9�w5��ys��zb p>�(��5�%�{��.�?EU�s��5�_�����/��%�u��0v
��5��?I'�O�(���2�q��$���F't�X����j�Clv�
� ��6OX�!"�n�)���1��L��9)h���R٧�п����w�X(�zw&�F�L)P��͂)]s���Ń�z�q�#]·���-/`D��n/����ę�����V���Zl�cu�O����L����UV�=��6 lo�� [@�#�s�]��K��&�R7�5�����d�I��7Eh^�B���s�6Z���9蠫���O2q
��Eu d�	|s�ZQL�7����V�H> L�\��D@ [(SBC��
���{�ov��0`+��8M"h��^�Y���wۯH�L��!�˹�(�����|��� H���V�/��P�K�e�V���Mk�$�3�,�����G����ɖ�;���yE@��!��D��}�J�8��]�F]փ���R��W�|Pi�7�Nv���������k9}#ή�Ta�R��Js4+�r�����?���Mjs�,hD:�lO>^��P��u��A+:��C���e�A�Z�H±��E8�_�W%�v%�z��R��?1�%iD�c��CXCn&�u�\X��7	��%ȭ=��+b��y���iZ��L��*���
 JJ73vr���d|����s��D1`��{�9a^0Z���f=�;��FR���yN���gv�XqU?͑���4O��i@�4Y���D���d�C�T��$c��Hw�o���$��>Q��_W���h���㡕-�n�_�8�� #WLӡu.��UW��*���G�y^�i+`�2�='�ფ>��Br0��j�A�ip�D7�e�1��V�Y0^�L'x�~�vGa.����L��#g{�)$�B�R'�fD�,t���t@==�1F��	�1�S4�]��P��\RGsǉe"�`�Y��"�S����(6�4d�jm�G��_�w-QC��셻C���W88:�qk:s�o��r����xܵ��^��� a����X~������&�����}ڈ-uﶜq`���!.lܟNfY\ �l�hs�e�`ܚ0`6���Ivo��U�PL��(x��R�LV2��/	� D:p�T���V&T��ѐP�qz*t��2)�x�%��I��)�#�L\�*q�S��J���pP&:Be��[��zQ��p�zy�"ƈ�VR�ѻ�CC7�U�삙ux����9;�#�H��W���\v��9����K�@����� E�Ħx"��^"�b# �Z`據���ġ�v�� ̺;�G�t�Uj���cם.�ah~]�0q�'��]�,����)_MU���~&ݳT�~��]^���n���&��$�F�C�����''���`���S�g��Q6-ؘĝt��?i��߿�1�ј&� �5���-(k�Pѵ�yF�<17�._��P�� �k��+���J�̻�1B��k7	��;[�|�t�L�N�|�BI�D�Exe�2��T�r��.�6�
t�sh��p�����aSٛ�'j��)��~暐(�=�х#	��$����zp�N7[I
g̜wFK���v������Ta`v�(�ށ��LU����$k�:�ӏ����x�DQ�C�!2N��d��D���ωM~��|d)P��)�IO,>�X�p���ȉM '3L=A`��,��.�(=��|4�XOT��8��{J Oڰ�,t6�Exwh&LJ�QY�V"#aQ��Nd �)�2B1)�VQ�Ӄ�C݌�ؠ�u�W��G�xei4�/�%��jzhд����B!��"+�(�K��'�
�.UQ� +�]zF���r��ʹ��� �3���%:����"%O�C ��G��dp`��ZR<��[WWx -�/��F����>�� 	�,������6A��?/�[`Ҩ���w����ɫ��a�巕�� Ԇ'|�]%�=&<Kp"�!g�דZ�G6��7,�+O���Ы���?kF�Z�e�Nt��S�uJ�d���s��|���@vx�QF.t�{&���UK�tN����1�`1��;<ep7VQ�gW>������F�b����W
�}�0��+��,5��2�#�o[A�E���ߚ�$^&�g�v�T׎��F�A6xt��^��%�����6��f���yk���֭s��Zʴ��	p��I;�Jy�¥�JZ>J"�n\b}��(�kӪ�l�$1�i��e4Us�>��i�o%���_�#�,F�m�ɧ��/�5ʤ�sIZһ��^\�!��5�����L���	*i�W	�CUj
�!nZ�MG�t�|����xE*GQL*;*ɜ9W�����Έyf�C�S�ŏ�
q�셳�o"撚bU��"�4�s�}��� �s����_+��2��a��H|��� �
3?�̬ ��oY����h�#F��*B�H��@}s�b�Z��b'9F!�.I��4��\L��4;�0�˛ygo&�f�Yx!����t��^p���ӟ���f�r;�a·���+�5�����/���nY0��'Ŗ�l�N���˷�[�Ӵ6|h]�zG����4���qR� ;���^E.��ɯ���:\9�|�0��+c��\T1Vy9>��{��N��|������8��Z���:��ni4�_vҥ*�S��枑��\Rt�D�c/���O?Y�Ǽ��o-ϗa_q�X��5�NN�"�Vo�$������]�VGVmט�,^H�I��8e�b�V����X����n	�/�� ���B1�Q�Y��_���Y�@_?��\� "�s2Ci�s��b ���=��`�a!�M�*��?\JBmo���Z����w��%�Y%T&<�(���i<�t�P��lz v#i���d1��}e�ѧ��[�.��g�:�L�p��-,JF��{ �0mj|za�e7��eb艅���FI6� sL���q?瞢*���9�Pn���'4���ҁ��
���9詗�9��h�xU
B��J��eCSA	*�{u�M�%�7��Џvu0���#�!SwoU�b�+8#lrE7&@�Y�6Hmb�F�؆�y]�[	�;���v��gyRv�58zòm��$I�#�(�]UW�M{UK�N��+�|P���b�1��π'N����&0}�q@4�G��At%��v����7�VF�냶dP�獎�A��9n)�|�@!/����i/���3�g�CH��H
wٯ�~��@����#A���WZb"iR����`O��
"6�+����n��YP�5�MwQNō��%,���*e��V�K�^��bW���w1��� DoM ��!�h~�l�U����v���L��5�Tim0�sxBw���ÌO����;��C.���Il�S�~�8B�|�Ya,�ݙ�U�3d"�R����Ð�ō�Y��a2�>U1U�,��/`x��e7V�-�2��rk��y��/���1Oa�1����> x�����vy��%6�����ȱ��^�lbx��D	�o��ӆXi��H�F�����<"s��
|2ɺ���@Xw���p��hǓ�	��%����pj��q^�v.�&��<n��ُ�:��jX�Gp�m]�G�`�o!��Hio~>F���[G�����v�A�*
�#IG���J�� kP>���w�lf��/z��D�sx�D��f��n����\�����C�nۀҴ�|!�k�#Hs�_����g��W�_���u��I��(rJ�Jnǭ��;���YږÃ�����r$�:xH>~G���a[*����ʤƏ�_�l){I!tb�+�X{�|<@(3E}���,̭1���i��+���*ɶ�}&We��^6Y/�i�.y���@�oOVY�������x;��
.�j(SSvpXv�z�
c���k�Y�I��M� ���-Z�P@�P�H�^����$�t�Ͳ��z�Q�~������lq0f���{]r�>E2��DlLv���}��sEU~RU�761��1Y/x���n^|w�9
����ͥԳ�+��I&N�f�~�%$����K�_��#Pg�t)�:�����Ֆ;ȃL�i���[�c7&;��G�"��P�r�.$8��f����/ˁ};�����n�s�S��+c�Z�Wz�_�{��oP��6�ˮ�����,
���#���bRѦ'9��_M�p���������(4���o:�~���*zWG)Al��%�J
EIٺ�b���XKM�Xӥ,���%9%���d�"2v���QY��,}E67���Ic�Q�Xp�`V!N.�S��)��>�Z�쌑ǡ���<w��S|�%Ո-��-�my�F��/�j�H{��=oED\ 6m��!j��;�ʂ\�G�Џ9b���4���N;B�M��0�g>k{7&��k.�f!
�.ZG�Ņ=�A�2}A�e/�:Xz:�=H�p���5���w%��ceV��qpYM���d�Aq��bD�&7R�	q�\b^�P}�zW�����w�|p��'��$�TA����#Jw�w���	���Ԭ�,3 ������zټ�)_�M9���rV?��7l:��J9��)ͳ^��6Y)<0�7[���nЖ�"䠤�/Q�-���`82-r��hƋ���Y�Q$V�N�0��~q�D�O���J�QQ7���|��f��R_t�y����9�����Tv�d`�t	�DG,o���s�{=��Ŋ�d���C���3-�~l���n���K�x��pg���Y<T��yRLn�/Q��6�	d���4��Ng
�D�1俯"�$S_l�p�Zj�b2*��-?��A�������F:��AP� 򻉩aC+@��'��[������W��'gꟂ8�ٴ����cG��,C"Kv��}�X��b��6�0�IA��O����w�ׯ���.L�����@�M�B̚�k'�?�]��_L�3���hK�����v���&c�Ym[ �k��a쌝�C���hVO˵�33�PȍO`}9f&h[jI���������qPi^���Yj��5&0{��ZSBA9Q)��}�\�4r���3!�����Gg�����ЋP�}��Q����Kְ�^���N>�y�@Fj��`�W$��(���O�&�T=n�Z�U�ʵ;�^���3]����?)�(oe�&jZ�	o-R�g4��fAh�cj�,h�A8��Q#�m��NGL�ƿ4��r)5�e��"lye*{�I�_ʳxʵ��=h�^�\�(Q?�y'ԧ�M���}�v���Я�]]ϰ9�e*
��Z��ߘ$˵C�T�	[�x�^��.�*Q���;��(����s[1m�|�v���S4;�zD�/���ᒋ�A�j�7�
z61*(������1y��V���at�0���+��@:	�Se8"�Fਡ��E�n�WZ"�[�Z�peȏ�h�/JqN>@�\V�l���G���c'
��1��a�4��=:(2���X��|���M��1G���R!����Gͅz�)��O��OTYqw�V�D%�8��;�,m_���X���u�ß�31-��|_ʺ�J'�[�y���&�Pb���Jݑ�Na��wt�$z�1;��qI,���\w:�t�̊�4�PP�77�qy9�fS5��D�S+ݓ��b�1(����!Ms��<��GK�r�3ܽIZ��0�G��Wݍ�m���o�Ȍ�E���;�d
��;��z�9j,�,n
܃ЅNƸ������H@R�2���%�nO|Һ�ζ���$���5=���.4��~���vQ~ص��M�� ш������o��ߣ���M�mP[Bt�������� QPц�;9f[�x�@w[D]}�x�� g|!/�H��;T�1���@S�k�d�gR��r�ɾd��踧)7�'�����R��`���U��Ok8<����C��g2��_bV�t�$��:�;��͓����M�^����C�ǌ��zģ��
�����DEE8䴯��(��!X�U!+��=(j)ѽ-C*��՞G�-bC���\E���S�i�7�mb9��w���n�kg�b,0˪�����Y�Qۯ��+��B1���o�j��-a�+*G,���G�";��m���� |1�_d���q��aa��z�C5,4�ks�MC�v�=��GVZ�,#j���q7����ƶ!��@��\�r'~:�Ŗ�$(�>կ��$��y���6���?���
���p<���T� ����e6����H��GD,_DCp�<��U�/�:�uŲ���AA@	w��5�,��Le�2ȯQ��>纴�c���)�|UV�$g,�8��3��<��D��$|H��<�,=䦋 �^3[��9m�	k�І��"2���X�1<�9v�H����3@i��нUg�C�(��J�؈�z^��c�C������N&�	�x�7��i捘I���%	�P�y
�����7pid@��$�N��\?ܸ������o�D�� ľ�7s��?n�>b��	�)t�Q8dC[�����U��y�n�
�x��<�_�c~�s�o� �l?$fΕ>��b�vF��(]4|h�#T��h�:�^�fI%��J��u	���

�|	�W!ҏ��0��,�����䆈�@ѣwmÔ� �����QN�0���T3���$z�����L\+ �6$Js3/�_	�>BM3Gh��3j!r���꫐_Y�m��Z�)�L~��R��L�wTc?Q��Q������B�MJ>�þ�G�����. ��C:���ط�ϢĢ(J��6r�9s���"�׮Z�����o�׫��&�"=��iK���)3;��AS�6����̤���̟���Z�hI��@_�]�X9�<Wx�l��bOk/�`�� X��	v�@��5��0l�����W:mL<S����g\�>�I�d▘�T fmd�bQS���K�X��T� ���9��nq�16�X��ƃ�S������ye�x!SH�C�nb�R��dڼ��X̵
H�a>�Q�'X�>����gF���h����d� R���N��Ѧ6ze��aC�/Z��6��^���6iק�V��$���M��X� H�=̛��cm���F!���%�}�Z����ݜ{����'����G?���)�O��:����<�/�W���3���|�^��ǬHF��oS�$�OR��y�3�$[�<?}�F���q�w�����n���a�g�
ɬ�����؞8��풇�F����������L��qy����l�hM���#���%�HҮNP�a� ��A�MˁE=y�v��Ax$?{<����N�Ӫ=�*%��qO�4>rR6��1���+�Tf`[YՊ��Or���������l܄��#�=���@���ޑ\er;,F�eY��+/�̙�n���t�\#�z���`��>?��	���>��"]�6���En��i�L!F7����g��%_��q׋�m�κOB-��vR@��$� s�&L�]�/M2�8
��A�S,����P~]{���<��w@w���ʖ�9?axU��
�]��vfm��_g ���4c��TU�0����PRh��'V�P��z��h8��������q���AzL��piyc��G<B9��j�9��[j#�:�t�tO�
"���S�|e�t�(�q��!*^�])Im��@��pa����iI��gy>��/׃=�蘅2��=��5�7ߊ.�DL�[^6��^�ѿ��t�@n�� ���D���c9;h	j�UE�xgq�4QK��a"��~"�U��@3�sA>�P�]-U<�}z�J�5�J��db�Q&���x�6�hQ-��a��"�tz����;���O�fݱ���-T���|�����;.��Dz-c�j�U_�-���:�EFa��^��f�F�#��t7�����`@ò{�&��+L�&�����d#��1rS���8i�]j�� �
�}L���!�pW�x,f�Ė;Η��H�d��B�'f"�`Ω[�yO9���7&59�pl{��{?�-��<Sg
[��j�3	�l󱴏=j]^��{gʕ��� �(�/��ǡn��ރ�r�T�v�Y^>�L>�HH\^�^�j ��|�5s+-T���L�%3���,�Dy@ �n�u7)����7>�v{#����W��0Ъ����������+��9F��R�V��#��TӖ	��Z)Gfz�{�F-֖����$���Y��,$����ܨ��{��]�W����忟�m`3��	�j�Ob�_���2�'?�� N���a�lF���C%>Uċ���f�^1�s��=�pw~���$�:r��$�b��R���)	0������z'��6(�lgף�hѢƌW���l�F�i��L�R���i���!�����-hxnG'ѯ�YG�D���/���� Y�7C��U�}���B<��b��v���9�y�|��3�z�P0͎�w�qF���n��ǆ�qlr���}�����#-�BC�|�dA����7k���4ᳪ�q,w)�ct���#�*��Il�|*)-��/�֕b�E��=CP��b�jt~-�}��q`���®Y������`Su��xs�T}s@���g����!vv&�m��R�c���AK}����^���E	�NȄF9-��|�A�(�U�^?p���N���/������̱m�>kD�����i�v��.���a$�'��9�k︚�l�l�O�t�-U�g��U:���pZŗ�P#���.ؕ�C���P���)��<� ��X�@�ʪ����oC��؎evpT�Ao�Wy�j�F,t�y�K�7�w�$?�J��:qN�ľ�~h�Ǧ^�
�9�B{�*״ ���f���'*���t౷�m4��L�O���i��Y궤������.���S��1������F�w�lA��-QMrPs��oKι෢���e̧�U%4����������7�j�8�5*��Hn����G����t�Iy�6��ހ*�൛e�|�1=8�)�ؕ���M8�~X� ,m�u��͌�Jjo�<�?#j�xP����?��W�)��-���x��=�a�.����$t�m��Kcp.@)��9i��M̒�C��Tk��Ki�чjw��s��3phl�s")�����u�"i��>�׈��u�l����A��`��������S���a��8�J���e�S&y�X{r
��m�.W}2R��mȇE����Fj��a�=Ӣ2mB]�I"��"!szgc�J:���2�r��D�^�Q!��	�>[ߖ�%���ȿ!�5Za�qBD��@�̥��e�v��Q�x1+�/�c�I}���*#!5��E��w�H����,��3���x�c�L�������p_k�<�������W�7f�u��=��\w>f��Ω����"��\vZ��>�;=,"�2i��u�����:F��x!�CK`V[�4��h�v	VX��*ZZ�uâ������
�B����c��	�W���iAӜ��3�b�S�v9T_U(8�w��DY	0Jڵ��t����H]�^�7���0y� ��0�~��͗��_��鮻����ߧ�1�����* wHp�bu�a�8�6����}�=��T[q��w,����ɻ�������_��0'is��%K�0�ճ����R��z����EM�	W[~+�)�u�.�z��x�%=!WX�k�X�T�})ǐ�{�{0��8�=w�/㫾�ӱ-*O`�:�DMU�%(�<鼁͗��#}R���Ë�W� �G���d#��r�����K�RJ/���RMh��1D���Oـk���N5	�\6�i�Q/V�8b��f墕�^j��%�*�pf(璺*�,(H(����MGO4��Xx���3�BY��0FE,��E�μ������᜖�
ƹd,�,��s�.e��I�����Y���ay�ۅ�u̔%57����.?����Ch�Ժ�vP1s���{{���2���*�v�����*DA3�!e'�JoV�����b�0;N���<�I��������@7/���ڟ- ��ـ&i$���qEcN�k,���Q�{S��+#w�+���9$h~�ǟLg���D!���ω#��@�*oㄖ��c��;��.f9#w��f1M�ު�32�;�M���h-Lz���(����;�w�5G�TF�O�=��"���"��T����>���;��$����/c޲��t�a�����*���<�"��T��F}���@�����H��w�b���2'�ш#9�E,�w�e-�B�o�ˠ�*��m3���0C�o�*�턩d�=
�]}46��:Џxj��^��I���e���M���u�be4�C!�tl֢o�2y{s���nL�(���ך�("�Ғ!�x�T�м��0"l�Ă~ޗ�����GMPH_/Bxc�j��U��6F�b�U�(GV�+RXFs�5-����L����`������'�\�*±ۯ��6��ČX������s,����ױ33B����������'ǂ|Ӱ�KN����vkA<�Lƶ��mU�Z}�þ��U�s���$Z��UD(5���o�{�Bk]�RJ��|��;��pP�(l_�+��l����gPQ����'�cd_o�D#�YV<JJ��$tH�z�'���=�JA��m�`���D�j��ȃ��B851tB¢� ˪�H|ۃ@��=%�cɼ�sGT1���}����O5�-��Q��8���0饫nG�E�D:P�	��{=(�� �I���^n G��'iKqs�~BW:*�N������VP��G��*50����`�Y�X���y�_�A�[5���w���1�0����'#3�\e,/�j�)�7��H1hu-�^��+����b��YFI�}�G�ō��̙Z��6����QLnCW����e���"�kʋQ�""*"%ڸ5Z`�H̾��8m�����IC���9���҂�F�x���0�TX�ղ~��,$;�@���ҌD��H0&nˏZgM�D^� �2pIV�Bx\��3y�����V�ߘJ��7%m�Z���ZY'�4� gD��gr�q��;K���D +��(���u�nYϤ�ƴ���ぇ�E��^��c�w{p�:���g���Slΰ��	�,���a!Iǩ�<7�l��w�|��v	�� ��]-����q��.���|�o�{�*���/ANF@UO����=��R�S(�ۤo��t�IZ&V`���I%>���yL�3������(�v17?�2��?O�)Н�k�_�$���67$p�z����>E4��~g�B�>��8�c�p�a��K}����Q� ����Cp�'��S�MR
.�E���j"����׃��M׮t�9���nt����6$�����9.؀i������#9����l���2�>-���XC��d_���y��8O��=������q�$�Fa��Rz�=o!@Rxm_'L4�+��q� N�T��3��Ǎ�Iz+�����@*a�]lv��LWy}�`�}�����Bt0�F#9���O �Ժ lh.���WY ~�9�����վnp�x����4�ћ���vd�-�ͻt�рq��~��[[!餙��I�ƭ��*��s0���\~��>3�p����3rѡ��j]�ᡯ���%[>�
&iC���U̹(So���������תV�J�I����';��]*��E�*YqY=ڒ��P��t�-Jb.��ˆ�c+�}&qf�A��^Z�]2��c�@���w�r�"�jD	���t��b[���g��.jU ���]����{�����*��v�%������Zg�v����)���=;��&��n�\�;�2��k�7�(�
��YUi4�7��� ��v_w�9�˦���C,�=���썖�иe��Q}�M�}���+n�'�)R�T���p:�j�]���Qf�□�"�*���܍s\�\.,O�lɇ�W�B��s���Ɂ}ͦ-����Z�~��A>��9U�&�Mh�QX+7�������%@�._�n����v�����Cp]0B�+sc�p���?bt�����ڼE���)�As��#��"�{���*2r� �F5ȪB���|q�3y�X�'1��V��(Ω}T�颖�M���cD��� ?x2��Yβ�G��9f�Ky�k�cM#�ǹ~�kr�R,僪���l�ۉ-������q*~j0F+BX׳��G����4�|�BY���	� ɠ飢�iK]�ɿ4��5b�CJպ����>�W3"3��xe�)�#WdP]A��#Y�ZS��3y��[��U?g����H!^I�8�r ��,g����I��Z�8�?�>�!B
��7O�ن��Z8BTv� �J�4���L��L����1���{nI���3}&�L�$T��s�c�E͟x�[{��+f��B����ȟ�`�Ԉe�Qi���c�6��z{<��B��V�|�Z���w��(�կ����`Ã�/�p>���V��^+?�W`#�	�Z{=�u1/F9	�a\BR;'�@�cĚ*�)2�,U�	���ab��/��J�ii9���HU�����3�K�:"�(p�s����
�:zK]�28��v}�ף��(�������u��g���kS;��M:� �R�oF���UR������F�,��Y�w�ה�K8W;������,�t���Ǚ����չ���lhOK Ɏ�i���"��"L�(��[f��#k!7�cp,4����t��5׊=���J6��/W�K7�!�}�QD4�Hy�W�!b��>g���Z�����x�HX��[�)�X����ҫ�Wi��|hՉQ��Z����ދ1�&��33�"R�]*�b&�T�^��z_2E��t��	r��Zf5Qx��
�=/�R���猊yf��Ѵ���y�co�#��5��A��9���e�v������G�`*D�-U7�\���$�g�J���+m3k�B,|ٻ�!E��w h���FP򫡤&�_���9��F��w�; ������eHAM�:Uo1��)���NP�	����'���x��d0�����tfq�H="!2��G�>�c>���ȸ�١�Q��~�Ȁ��x��r�jj�<�.��:q�ћ��Z�t�q��X쀒���[ᑲB&CW�a��1f�)߲����R2Q����o�_��]�{���Sr�u`��=P1ݬ��Z�N�PʐF�H�K����s����R6���u���#�G� ����飢C�4�e9+>��%���R�����,��h��1�|�:�J��X4i�#[2�!�.\�D���d]3�C���o�ѻ9�g�a�,����"F}^�Y�_xb�)�\bu�-HB�c��v3h�7��[�DjH;\�H�*&�����爣V+ҡ�q�h�'(X1��|3��X��e�����%�=�`��R4��_*�-�. �����=2�5�D��֢B�i��a������*�Jxڳ�m���&igLF�p�e� ��u�f*�40����&�����ˬR.u��'fFn�){D�f諛��gsNJ�Nh�궑�Vo�_���6b���ԃV,�[��&���=Qy�2�% �5YΈ}��(�cW]3[/��,3��^��\��W��٣6�5�:O�-BUbz5��6�?`FC/���Lӿ�"�084D�Z��wيᷡ�u���ް��%�c�i�Q_U��'�j贔�����ːp�P�`���,���*�SH�̯ɣ��M���Ue�|D�O/G��]����b�?�������S/����e��+ި̪�WY���9䘸 k��7�W�������
h��8�����"X��3��yN����,I'��l��ů�m{_�{h�G�Ϛi���H�$�k�\"3��Q)S�0B�5^�_1��.�s��!��?~�yH��k����">v��|����8g0c�RV��t�;�VgM�S2xv����i�K�*J�i��/�y.�=ߵ���ܱ����䆴�;�Dv���f����%?��������8/����u/pČn�^p�l���C�i�����w����`�4�Xw�$Z�XĜ׶�J)ta%'j7��4�sv����x��菣v��\���m��C�dP�����2�\S������.*)��d��ݬ��5}F�� �A�Ȑ��F0���>�-���]0����[@Rg�(�R3�!�Nft��\�o�*ġN�%��c�7�b^s��猠��7ub�� ��4�}�ϻܵ�w���n3��a�6�%� �������0͈���Jo1G>{�;���ɽ����PBՑ��l��f�J�ܸ� w�yF��({�n�����1}���V'�'��K�/}1p%9�j,���p`�$�3�Fh1������|tS|	���b�vt�7d�Sh[�����~K"�L%����19�77 a�CQ��e*~��D�hs!4?f?ma�IX_���.FՖy�VB҂d�:$JM6Ǳt�f�_�i��b�V�Y�����=zYPR��S���D��$(
AȍQr�����0��B��0��c���o�����?3���X�8=����rBu�M맛^��`('e�>��A8�4�*��u&��~�K��\�ݾ/L���]�-p r���/�T���	.�D*!8�A�E�,~K3�0sU=jNL�6�7�-��*4�t�
|I�%�]�����wk*q���J��(��,��r�2�N��'R�>Mm�Z~���]�M��ʎ"w3G��E�z��^!�cx�i��o�i�˧}��D���C��aR����jTY|�|�⌰�J3	j������=��O����AT�ӏ+�
�:���n�N�Uxᢸ�=��΍���+wJ����/4��G�B�Kwy� r&;�;�!*�����c�"E۽�0���S-K:��A�/��}��>��A�YN�P[�-E҇��M%�ֳ�w5m��]�Eq�C/"N��y�[``�IE�z����'�-�ʨzT�}�DU^�Fp�Q��*�H���L�*�F�A��-,믋��߱��h_�6��c�.α��9���~����r7P,��nw�͟P��z�xf�� ^ǰ><�T3�B�E(��f]U�Hl�_��x�i-��v�q����;�!A���8����x�=�d2
�k�s\����L�1;�,-*�m�5Te$yۏRG�>gh]�J�C�]V96�å)�p\E�{�n���0��#=_TU�����°��]�%I�x���~A�T���˷9	2(�MjY��*e��Ȗ�^�Oc<-Qd,���{�_�X.O���Y�HӁ�& �P<G@@UbQQy!<�
(s|ҠW����FS�xR���0�����e�+�ݢ�F�8~iu!�N�k�i��h�i�O�p�]}��}�`tn��8������N'0F�^��fn���N�׀�,�� r�|ʎ@��D�)�w��N!���5������a՞�u|}9�:f��c/ܯ�HMGת���#Y u	[E�dz��qB�>4[��(�T��c�=G51��2��	[U��!�@T�OH�[ݜCey�����mRl��?z�MURi�5�(��'8o�"�R�����К��f<w�9<�`�!6�8�G�@u`���b!�($����T���ė��)U����f��w㎩�;�Q*�.��1���[,�D�|�F�e��Z� �f:�8��դH��1u�=�u�����,��@�"���H2�fѵ�`,ou�\5�\+7X ?i>����fr���K�h������2�V�_PSߏ�Ad]*	��o�����?�4��a������h1q��t<��w��i4A���c��<��*ˠu�Uwux_����ɚ[�7�5Y�a6��1_Je�%u~m}�Ы��usg���^"����^"��?��K�U��4�z}�aoVI��H"�Q�]4���(K;f����G^�>Y�������-�;!'*qX6��α�1�>�+?�~gJG���å"��Y�{	�i��L�iXp��$��	^�N:�b#C�=�k�9�v�MU8�(�^w�p_MGM��鮅��h�+�8)!ei�3%%/;�q��Ǟ<\ �<��/��2G5pO���@YCg�¯5�Np�}�6SͯT�Qv�M��FB�#\�U�V��z���VWXRR���3�E���,�F��!�Ì-�=L�)�a��M��y�=B^
�O���ɏ4
��I��n���r$]���N�S[��CM���h�bMF�F �l���p�Ȓ����1j�E���W}��@����ڹm��sR��*�>5�&Q�q���xA�'{��ߙ�%�b�r�'�C"YZO`H���CE�Ư(Z�?f��j�'gF��A��;�1�����#�䶚[F����:Z_�6p�xC�o<��!�kS�b����$ko�`�7bM�mş�;I�M��ۤ�ɤ���\Td_v�˔��6�R���Ƅ\��=�fv�[>��!�w�Ή�G]��'"̇�"�B��f)O�Ԩ�	"�GMe�̻�|C�H8�a@t�g��ov��"���%4�~���������
��&����;���ty��������f�J�l3��>��n#�8wi6�z�.�C�0�Ь�NxT��k`\YN�w-#O������>��P�(��/RA�i�4$Z�U���z`�# ��Y� ^��V+�;���ԥG�H���q��b��Z�6<���̯EJ}_�JBk#������d����z	L��e��S��H"(\[OͬP�=�AH^��q���mM�"��]�: �z�_"®�Y�{�w������Pfs�yk�>1�ep��;�&<�g`�'����C!�Ń�]�Y�V��֯a�?7������fJ�cW�r��*ȇ �MwR���|�$K���]�u���Y�.�jf鼍����B���̤|V�.�˥���Ѵ����Mg]Ns����C�ܥ��t����w�k��:�A�=�5Rլ��f�H�u54B�(B̐���w�.�&n�U�?F�8�*��1�k��!�'��Z��ݦn�����p��Ǻp5ew�քLm����ꃺ��[e�<Ӑ�<6=۞�fU��Y���HZ�
�<�������H℣n�F�3��PRQI�v�*?��qi���3�������-�C�q��|d�D�F2 ��,����>������^��]�:�&||p�%-/;<��M��$�z�%��1|�nV�4�Jqr�X�L_��^po�J�!/@?�I�6d[���҃=�����0.X_��u�FO��W�E�I��Y�T�|��+��1����X�4A�䕼p���@``Ro� a�k��X��3��s��)HyZ �в#�=����UD3����&~�MH�<�^�8���n�
[R�1��@J��rY�'����ਯK�e�5ǩHW�|*�b1Ք?V��6��A�� .��������4WZ�{�_]�F��k�	$Li�C�6�/Hdv�s���x��M��B9��[�74��c���H�U�yM�wǰM��|���w����6/�{� �U�;#[}����)����d-��L:�"������d�x�Y\ngl���8��p-
>�i-S6ܗ�l+���J�].qN^�8!E�y�R>���))'�,Wg��%�nz���l%�������_�1���Z%� �qH���FN봵ȹ/nO�ۭh��v aMv
���
П:Hثs���*��K��YJ$|���ጀ���#�r����%Q��ar��1�8��U��<�j6��(�gV�5W��Փ��]���فnݥ)����4D��E��,�9�G�	�U��Q�e�ʓ�����^��q��� [H�*�90^j������:�@��UF��bǦg:�)gwۛO��;����IF0v�*���8�0�)��A}��:@VäY3��ؕ)�B��qҳ9�n��7����˜�n����U�4t��;��E��'�}�� �ū[�E%_��1y���ɡ\T?<�@���1u*�hd� Kj�N<;R4�Y=�#'��\���Y�z�L�iAG�I,&�Ŀ_��!�Ԣm��:�q���R���m�j0a�^Xᬤ����Y�y���L�WNXpN�b�e%N-�B$�3�?�RI����H�e�c���FZ2bO߇0Sa?x3Pn����ٚ�+���^Ӏ.���7 &a��RO�x� ����T~h|�o�7���!ˣ%t�H��z��6Q)��-2�E�
�=ZwB���~�(\�����r_*�ܑ�>��tu�/���;�:Uw���Z@�"��k���Pï֗��6O�qˊkܩȏ�c�6Q� r�Dw*4J�?Vr�/2�bp�J�q��D^��Veӝ�2��y��4<��$�1�j�vn���y��J���~`0��!>Pz��w��)8Q1�Fு(��s�Z��\��,n�j�� w�H�Z	�ȝW�w�i��1z9��A�WV!SYy�[^y���͠�l��8GK�7n���������#C�僽��>��Dj�WE�4xI��m�r��q�h��1V�Q+U�O�)�|ړZ����Gjmq��E�v]�Q�D����QQ�@h�E<�
#*�;lUʭC�ִ�{ƛ�/�����?�'Ư��>�b.L�d#�%ZY��W�,����9��9��:t��/R]5V��pd6���x�ό{��  ��/_�2=�i�P���y�+�w�mς��}ԯr��1aGJ��B��M�� ����G_��8��^Py0�n�D�V0T���As*N:lI�Vo�j����܏UKA��uK�L�ٍ������(��.��{�O�^�?�K����PO�e��|��V�,ˬ8W��w��珄��N#�q<y�%�f�D�N϶��P���A�=b����$���[v���z���L����Կ�F>��!y��.	����`��f�S�E���XUA�Pe��
dL��W���~2b1��>1E"��<�� �Zm\��]��O�D$�(����a�!�-��+2s2��D��:�;9�v��\&�4�}C���ك�"�k'��V���8�$~����I}���^H;_�Ҩ���r�=�*V�o�����ˈ���o6����*����X���"F 2�>���W9g�E�ͤ��Ah�XJ�SL3�'_���M�}C�,3!gAYԫ[�����x2�f�$1���g����śd.ĵ[*�B�O�A�A��K����U�g3�,~����k���Z1/���P��\~q�kg:�����:��)Z�¢_gE�-�a���Ee���j�����</t#m�����RK�b��1�y,���.�!Z�5K�e��E�q�����AF�y���=p�8�>%�e'����+F� 2��W�+�U���"�$�u֪[���P�t����ʒ���k[˭�	ގ�Uj��fZ�*��������HY�W���;C��gd`�'}�@���������I_�Y�
�{��Z�G�X��=Y��t"�� �M;0��U�ە�PIwf#�U�vW	��|�58ʢ
�;k��0�Z-���IS/CܤO�͐��_:��I��x�2��©R�湩+�;�{"��p�s�i�9�[(WvL6�DY
%E��f�����N�Rʏ+̸C�7E.�'q�hm� O=�	C`�+�	݉�tW������{��}��ˌ�������D���S5KLi����x�m��!���>,`��u<=�,�E��	�a���/q^l!�����8���?���|?�f���Iw~�ЋpR�[KG�[x�sR�ԁ�х��;�m��rEX<}��C71�/7j�0S�ŻN�!x�aj����o���k��6�`g>R�����k�q,��ݳj��1a���J�Ǟ�c*����}���i���pr��\9�k���w{[o���O��Ւظh0sQ���R`<J�A�:?��Ÿ�#fsz��b}|�p� X�9��=�!��1#�[�-�̵Xv}6��|u�MK��ꨴ_��9F���+�B^��H%<n�yB�`#���}��_�_�/ruߐ���#y#�[�oˀO[��pո�/=�Z����0�L$.�9/DR���{�S�2��6q�יgR�2�RrAg��}	�^:�yMkĭ�ME�CZ���yd.�����yMEt�l�͖�uJTo6%��w����H����<?���{�m�9t����m@\�J�d�H�i3��	�WL��2l�ĒUtt���K_!Xp�� �G�@��E^3��tj�W������v�?95�C��hF��+��qB3+8��Q�@�q�O j���Z��gtw	q�lj��(p��0��Ê�Ū8��`�9�����Yf?ʆ�82i��[#$�䗈�6���k�`'�� ���ֶ��)�L�ޠH���1�<Z��N�*,�ҵ��e�Bz�@���T_���)z%�d�A�d���`�B�z�"��)�w�˲l�����;M�y���cV�5^�nCtoN��^���2�kUf4���r��f.��KcY��PN7�d�FA���?�y�󾨌�Zl0y��;zˣ�a�ǉxC0.�IXᖺ�� �0_���a'�[K����>5d��3�ai� jh���0����c�tx����!���3z6'{��e���ű}�ts���RP��(e�d�w���>*7vt"|3�4	�}�+~��E�P�s�&<h����H8���
�fYV	�1;-�Q��Kc.'�r:��S3�)N�h�i���(ڱVer*o�L�#��q�$G#@�3z����7�N��IΛ��Z�8A� ��p��;�S����	���:�^�}'/DN���p��)��:%B�#��,�E��P����b��pR�j� ����䝜uK�5\\CN�BȶA��������\d��]��$��IG���npz�Lq�J��dZ;#h�L{}
m�9[A��j��������n�ͬ�s�peIA�����܇�!W7���A2�����P�^������p��D&i��"�;Q֛0Q?�u�PN���
�~��	��  �bM܎�*r�|,�4p�D0>$���E��P�6%�P�j������KB�遦p��-��W��%B�PY�$S��`z��0�#U Y�u�M�����2�`�g�A��2U�]�6�b�G_p��%��:̏��v��v�>�{��w|���ypy@�R��6�{�����|m��?4�����P��m�S��/��&��u��*�藞�n��9��ށ��������_^�g�F���P���[�A�AT�����o��X�?E�H�%���F�����-�Z��X����w��SQK9�@8�O�5k@~�w�;T�z�����/���(і7�2����~��Yi����(��6PD�k���@����A]����S��f}���IJ�X�1� 2ք�F�����|��燞���E�����B@9@�lNK��� �)�u'k+�A@�,8hA�CL@� v�� �zt�����N+�9����U.4C���ŷ�^��NU?M�}�i��X���*���[&x��ٹ�#ge#.eh�gY��s}�@�E�F�m�7M�����O����)�t���0���8!�8fY!�
QIY%N���ǾcZ���� {�2b
�)On���-�Ӂ�r������=��� ��� ��D�T�S�XS���M�x�#g���_/���g��Ò�������V��z��ż]��2,�h����3Dj��z,9���M��t����ZAL�v/�sXd�ϬBg?\�FsN�u?�5h>}ދ�����@ܫ�>۵�ǌ��G��mke���r���(�#�{�|���卟��Σ(�`y�i6"�WJ��Z���Z+��n/ж$]���ny�X�� �5i��؀���+=9?/�t}a���M�O�
G�q=Q>��n�U}��W^Vm�sj�S��-��16qoc(D�f�}��+� ��=h��{D��X��~�C�D�+�$� 洬��4��_.�_pC��3ؗ��F@UȔ-�c�mf���´ ���p��7� �psnO�O�yo��F���������EO�9�
�<4t�������9�~��Ӹ<�zP����`����k��'{�0kU�1�hP��W��&lT�Lu��.$>(��2^}�����t{(oAl��,KLy�Q5��19��lL�=P���s�Z��-��|�(b9Զ:�>�¡R�ʢ����7���)߰h�Y�� �;?�KG�"�3�GL�#�N-�4�Fk�dW�1-0s�gn��n���}���'Gp�Ӑf�"m�}'����Uɀ����tS��c,=�5�����=�Ʒ ��o���J]M� '^��hW�e�]M�W�4ﺐ�n�ݘ�V]J�@����Ix�c-��b�+DFB�56k Z9zW��;��cm��~>�������vB�,C�M�i٨3��}�i0���^!~��=D�� ���B�����d�氘.�!����P4�oR(�2�T���f�ye����l�o}�X#�(���t_�33�Dhː��ۉ�)4�i��Ȼsu]�.��<�o65�<%�Ss;�\�YƗ�Ȯ @%�28=�\1Z�y���Pv��Âv�Ҁ5�
gH�� ��V���F$��]�.\,�A�,�yK�jĂY���s��.�m�v1���W��[̆�̰+�'���y�r�/O(6�Gؤt��V|������ʠ����ը͗�b����hGi�&mL*rMa����D�� t�ܹ��i�8�R�8%�6I��r������A&D����ײ����Ow��<2Ȃ!s�WFs+lk�Q�.O��0DW���/��D��z<҇�X���:��\�ā��-~~�_��i%"2��23J�sd��x�s��bC�Y6��y!ϼ�\^�o�HZ�3��/Q��rM	�!�Մ{
��ԊQa%����rPQet���h��锃��ty'r��k�E~(��-��n!������X�G�-	,P��ar"[�,Q<��䫥�Y��w��t%�SI~�NT~��V�z�ҝa��b��3��+�|�ƍ	Di����|�ѽs�פ�U��6Q��Bq��`qnT�
�Pĕ"�~�|�!� ��U�x�0�bēl{V����W&�4�֣	­�Ts���dg�h]����gc:�����qۜM�� �כI�dwu�]�?��u����%n�F%=xc�P��;f�m:�oS;�ϏA�n���8��𲀎�Ӻ���P8|���=��É@��V��H�g�Υ5�v\�l����~���x�[�$���1WP@S��#������X�d��j\��
�[a/����U��b2રA[�90	|l|?ݠ�+��=��86���~wA��ӹ�=�|��%o�XE/{��x+(�}P��02r����X�m��
?��ڛ������23��3v�e�둡��@S��RdP��{_a}�z�d+$�)�5��/�r�C��O��Ĳ�]Y�-���x}��F�|�v-:�5�S>���~�#�� Ş�	���Ks�`�7ɗA2(�qQ���}^��,��뎵R�O4y����;|�Ѐ�D4Q�r"�8�L����n�z�L�t�WĊ��{�M����ê����$��= A�ҟ�!)�8�Pk)I�O�Ϋ�[˓1�$�S�o�xY��ܵ�� ��K�*��T�P�*�^v�^�wKB�����$�F}�CW<���RcS{�����H�1�^21&�Ve��Egm-�Z87u�.�r��s��3�(�2�`������K�I�4����jC �
�R�U��b2�%9Ϭ�d�Q��Ԫ+�t���$�X�iI�D�o�K̥q[,l~5�Ք�8`
>����>G%d�#O����ADz�m�D2�x�I�	�s�>apx �n���S��~]����L��V�G�J��qɔ�L�E�}->�ke�g�r�<����?~1��ÿ1����i��M!�\�i�p�bs��5��c>'�2�X�����־��Ъ�����'ݝ��i�n-{��O����#�[/
5u<��Z�a��=���:������C�*.h�)f��2�w`N��,��3,F	�"�L�����`h�T��	M<�&7��tc��	"r؀�������� lK�a�P9��6��R���\c�W<1NmW�u�\�B�ڀOkIg�6�~�+gV��ȉP$e�ԏ=�S@xj�4v��tִ}9N�p?!g����?�t�-�
�id�M1��V9��CWܷ�;�L{�1�9���v�	����'�2>��ݭ��Ly4��'��~ �W3K��5�a�ɱ]�CO�������t�0NO�L!{���ض��I�y����Ơy!�lg�P�EC2�B�p�;�T��߽ ����V
�~)S��L��y��PԎI�O<4�@�r��!s�ŭ#C���<� 0�o�W�8@��QS�l�gۣC���\��i�����!�<|�zVb���i�7VD�w9�`4\�]W�{KF%���Dj�q���]euj[������A�xz�3r}r��fj��!�*B��S[*O�	��&�@���4Z�S����L��=�G�xX������#�u$�q��V�	� ��R�O�����j�;�5�������P�j�m�8S~�ϐ|3�]|�g���$�������*r{�P�յ�)����u��
+4uD��A�$#� �v��}2��ꜙ������$�M�w٨�-zÍl�4��゗:�+>S���i'�݌��и�T�.���.{�bQB@� �B$JH�)�s���a�K�P� |!Y�4�\��J>� \��Ƈǌx4$��W�XĜ��E��Bg�<a���F����yR�p8-{ϣ)"��)�G�bb� K�T�tl�3B9K
�%�uʹ�A���p���&���D�4*FL��x7���.a<1��NZ��a�%{i|A��Qb�XClC?��:|Y�#���W]�}<,�OSU���A�34`m��p	��F��ؕrY������(}�-���u;� q3
�!���j�}�"��:����W��6������(Ш�߄�~�,�oM�Uf�����n2nS�닒иO�a�@��b�]p-��^�YM��
�$%|<���ϑ��yPq������� &M����@��q�	��s������=9g��R�M�5rR_�`��)����=f��#��O��PFH�w��96��ػ��� ������J��y1֤�d��6��<��.<�����<\
��Gܼ��R����=�v�s3 u��Ƌ�14mCb�la<5I��v_��q�z��	��ި=��v+�Fff��f���]���w�y�lY��
`y�碋�o�Fh���t�8��?�l3���+��N���W<L��p�nz�H:zf�e�~��,����^�/��H��A�ӵ�;��=���O�����O
w�d���Cւ�+�}#l�=����߀���cE��A)�L�rJ�͹��gV�S�-B���n�5E��N���*:��_�d�nK�����C{����\`oAE�M�1⢿>���v2<�@99���r�q�(�l?��}N%�v�� Sٗ|>R'G~��f��S�?�nx��e�����DX[�w�~�Jfc@��5���ؐ,�츩,[�/�� �{+��-+H��4�c�k��"Sx�fX�F��v7^ͱƶ�٘��?��tv{ʣ�	X��`D@�����"ug�B^l�L����<�[q}OU]�l�G������r��އ"}�w[ĸ�zj�>@�ئ�-�V�g� �Wc�DӰ�V��i��,�ǆ�X0|�X�'ߖ;�j5�SPү4������;�$U�('J!9X�v��
* ��ѻm���O�H���6ߟ��Z�z�&����
���W�q��ʨ���T�:�Ed�f�_����qW�O޽ъIP�ݝ���T�>#�U�B7�h��3���N��)_��s|��ߦU�+��d���{����?�%�w�^�c�M���v�*�� ����h[Qe}�rc�%��4`z����u�Ί��?�B��EnsO�у~p&�QD�v�E#��VC�a�W���wx�#n����DK����ﮎ<��P�0�oRţ�h\����i�Z�eSb	\$eKt5k`=:��ss�f��c�@es�@I��&孇�p��K�n#,Q�{#�*�9��p��ύ�aJ��v�y�sw$�I?l\Z93B��*C���ar�ƈ1p=�b�b�R�D����E}���K�� ��Rb��10&y^b9z��X�qV.�5��ݲ#���M�4a4�A�v��vtT�;|n��($:)��0��r�`�٭pJ�����N� (T�������x0�K@F�qzM?����ӄd-	$}O�9���|���Y:�𪽒��|��~��汼uiη/��B܈��p����D�T�7|2'���)�V�$�y�� �GhR��<�ذ�c�ɴ<{�!�@֯�\����kJ�"��N0B�}�[�>�腥"���-ɝ��`T�v�@tm�q P�g	\Y��º��@/u�&4LX�$
ݴ�m�$�t9�t�^s%ֈw
�k�@�6 n�`��^kIw��E킲*E�)ӫ_6��f]?bN�@��ƚ���}���G
�6�V2d�t��t	��}\��&��K�.���k��SQ�_�ٙn���a|)��vity�k:'"s?Kz�M���ٌ�(�d�;E���	 ��?-qf7�d40���\�P－���L#���&���9ڃ�r��O��x��#��t�	� �R!�?��Q�s}.�2��������ͼ��b����)�f�R���|�"��y���!$��\���ۦ�B	��l7������BZi"{\�B���7k+�**8M�m��]��5�TPt�PA�I�zT<�Ew?���rHh(Re/_(��:eۯ�<�^���ԟ��]Okg.���eB� �MK{S	��y�q�nє�S؃���B��s��b-Ty`����O��7h���)4H��X��C©�Y� -$�4�Z&��ݜܓ�-cDV����EF��V�I�t�ܪ�mk�$��5�/�+�Mc�]� RJZ�ǲ#��:D����uI�C=���a�aW��?�=@��V^df�+���X�0%'��a<����W]}�1Y|ړ�rL����>@���֙�O�:��u0"*��r�>�nlCsR�e�W&�l����<r����k)ܟ���ԝt�.6fM�?�u���]gA�)��XJ�O��}��XG�x�)F��)�چ�����OHQ%�0�l���%$|_�hRU�	�ƺt�Q�SU�@;,̇� ��l ��
���~�$�7��c��#�ZX ��	����\��c\�d������d�	�q��}9���z����M|��D���I�������Z�"��E}����F���;}Ҏ���?��n@�����	��yfv���ر&�-��x����"-�,�FfOB>mO��R7��߈lA�|��O�C��$89�'C����D�ݣc�q��o�b��.���}�g���E䠇z�c��Yo/DT�Jm"f�%����4��v��/��@�f!����9f����0��#���ߢk�=?��\��Ϫ����t��F&�"[�Vi��X���<$@�
��6h�?�ߨ���/�/��,چ���T�!�7h������$�t���?�Z���n0��1�'��X5�����R`9���U	����,�؄+Cu8��훏��9�_#M�RlPPO��-Z��B����U����Y|�,����<�<�o�|)�ƣ�S�̝��d݈��/�0��f�{M��+!������o���'RS���M;E"�1{^�T+�Qܯ�sCEX"r�>(y�z�ٞ�����W?�1�R���
�