��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�uwC�5�b ��ϴ�	+�
Ct� "�J~���z����<
�����'k�z��ߵ,d�.��Z�Ӝ��2�x$ҟdL��h��ʔf��#
����;�;m�ȋ��[F��E� &'{=u�3jg�b�)��LA�u/5{<	����kk4�w���`+D+_�,Yw���Lg����x�*�����e+H�Qy�8�	���4^3�f�hOi3�Ø!��%���^dWp��[gN��U�v2�S���N�l0���V��IF&��c�eȫ��o��P�wH1���dm*n!��%i���6j�6NU���^<Аa�
l��q����{�_ ���ye��x���.a��_ﳐ�2\.�.%���`�دJΎpz���٩~�B���B�����7�%*�BTT�`8���|�X?����ҔR�2��i��͓!��~�6x���,4"ɘ���rl�߂J�]��׏��sԺc��Ε�_*|jI,X��ć=`������ߨb��F�t�U����sg����۬�Z�Y��hB$R��(�#8�^����
~���1�D4�	���{���(,N&lj>k���` y"dب����C�y��jε<(�&.��]�ѸI�ড6y�NP��vc��P!qsif"�:`s��Ag�V�#��@4��},��u�LOM��
�U�+�������e�{_�f�_�=�+��oþjS�1��Z��"z��{��Н�^�r���^7r��x��Kʿ �����b����iΆ�f?,Np�$z���T�.ԇ8���E�SF�.&{����.	���1��ï�3�q�	3�ܦﲐmA�#֞�����2��`*��5Q}��$/7�ŷ4�k��O��`kT�#n�V��|�,`�uF�;�%twC�{S-�q�� �C�޹j��,��	eTC�o�v���~~e�����w�K�v :���JA;cCx�l�����f�-@غjDhbX�1퇹[	�H_��������fc�g�m0���mM�+��֖{we�~}]cE�)��.����ꮩ�W���u. �d�����p���N`l ՌeP}T�d�m��<fe�&�����}�[Il_[�M]�(i!��c@q����L٨#���#�������yY��+�iG��[N=H�"�F�0�)0#+��X7��E�|U�CF�':{�Mgj�A?뭹�G�s��W�����V���0T���i�	ѐ��F�m LׂY5��O}�!��������&�II��H� �.Sbߺ�*%��q<g�pa�O�9��u�O��=?[T[�*��O��G\����t�S`�t�5���(Ժ���{hy��-#f��Q+��~�Tl�p��0����͵Rd*K���*u»\Y��*��p2��}�W��D��RH
Ln0�ġvv��ܳ+���[�-�$���0�z�� �	�r��[�x�U�?�O�]
`Pn�s,���	?29&0�вi4���+� �k�8RP&��g��~���>��;����ۢߞ���bԤpOg.]�0;� qj.�sn�=�ߴr�����l�'�\��QH��+ý���aOZ�P�P�]���&gU\9��:���т�wu]�,�)>�UX��v�Ĵ���z�bl�L�B�T�XvҀ����`�w��u6��z�!���{����	]��u��cx�s8x<��*:����Q���|�OX`���ͅ�y2�l/���М$A7�~,R��,@�בr1-h�nv�p<�@R�R����c�?��QR��7��
�*j�eV����R�7m��\�S85!Ȟ���Մz�EdғFg��/.Q�?�LP�!�CpA��,}�%��Ä)9�N�̫/B�xe��
7���>]�
�Z�מì��F½�~L�Ph��ՠ�^I9]�i��?��Q�~��(R�����|`]�w� ���-��6Vi�c���Q2bVfg�4�
|�Ko{�B����#��/S����xG�Y����9.���̈QQ��-��L�y6��1H��\��&�C�2ڜ���<`R�w`�7ۄ7Õ.F������ͼ�����ȹ��RS*󟥧~U�Qm�I~�1�G (����0H,�KO�,�x�S	w���.ܘ�����BG�"���ߧmW_{X,�Q��W�Ҩwi�g�P�א��S�	�$Z�z�o���K�r���8�9	�]$�
���z��lLuB!��� �ww�3Έ�_|'n4"���?�T��76Ts�^�X����B���!�.	��h�{mz�i�[�j�MZ�B�ך��ۧ�\r��uN��K����e��_���j��>���,N�W�ip���cb�>5,�b;�$��%�C�+�
�;��8�S�\b���9���S���F�t8c���P|�\�������[������J.��t��k�i�qsb��f�J*�3��h�a]z{�m�<������=�J�U\�s��(���%}��g���b��[P<a��׏� ����:��:�/(0p�M���I���9���{�-�(_���'���'��/b� �fϨ���^����i��9�J ���/Y�[}��1����Fƻ���P�����wy�e$���ɾ��F�/��ĸ�~��9�H J�d��������%G�Wтx5���][17E<0�@`v��TH�����=����Ji�)�cwp<̣��w��կ_�:�\�E~o��{�{#�ݭ�R7〬ծ�,xE�:��")�v�����=�	�W��P��,��GQ�������l,�*6"�����c9�D�VQ]�7�.��3Q�Q�q��kN��D�},d�b��vpgb�T"-N�B��!D]vki���}� �^5�$��.����L�"��KP�	���nr�b�W.cF��v�|С ��9���{��&!|\��4�k ��s:6Ec�X����o�Ҿ�G�O��aI5*v��A�4�"'�:��=��m��|M#�B,C���6x�p�yp�E�smؖ>����:>���DH_h)��՜����V[˽��pm�oL �Q��d��(�^�)LO0{����/��� l�
�wO;8�olB]|C�ݫh��Z�������|��pE����%�r)ը�^��d89�c����T?JwXz~a෧,u�&���3PPX���֋�
�ڻ����Sp7������n9�<z!j��i
�cJb]qPQ�CIy{�Wv�Bj`�������4�4�^ '�o�ܒ#Z��� �9E��rO��#'{���D�֠���o"��R�~�l�[7�.��qy\�{zD�oDq�+������g�لS�
/ڏ��"4�u�v_�>Ub� ��*U�$W�R}{k�g1�ō�:�`=e>�i��e?3֧a�R��7�h�h�{��F&#c/�����Z�����O�2ϧ3A��o�
����Vl�<��+��Ɉ�f��2:)��u�N��H�!D=�;�n�('NC:
���ۏe7'�� O�(J�v��7O�,���#���A�y��q��pńBO�]���R�h��FtK�^o�cV����&$rX%�1/�H���+x|�wVK�K'zT���6��+ՀS�����X�48�"r��Jlr����U�|�w><`2��?�����4��H�9�X��}��2ZgŎ	�nL$,�+��Dۮ��y�ݞ���D�̽7��K���t���g�/#ԊS�{���su�bE�MDܥ��Ǒ�([��u����@�FI��>F�nf5=p)<�I&�P�]�D�t�?��݁��vi�׿C�ʖ�5���t����j�1�t�;qfLȒ�����S7��:=g;ʏjܔ���@@G��)r �'�E�i���J�1����fg|D����hF- ����7�U��m�w�gH�*�6VX�521����?�9{�S$�gZ���\!pJ���kG�0�.�?��5�b_R�h�{���X�8@�O�=��3�Nt���Yke�bdހ�O�4Z�US5��v)ȹ�C�Iȏ
 �S���W�^4G��
>�L=:��P���&�Ҍ�6A������G���v�5��Ẋ5����ϒ|ݪ��]���]=�z��E;��;��?�BX9��U@�tɬo����FJ/]{�f�	54x.�	�u�����)~��[vds���f������*w�(��;sމ��;)A@�����n�K7�����׫����E����>�;BT�����	�)�?h�����`;!�������P�����Ç}~-E��
�I����8����*{K�R�)ɒ�݈9aR+Wfv8*��GyU�l1m�W��HKH���s��*�Ƨ��ꪌ70�>��ʁ'�r��O_��>"Ր�:��G1;i�f��Ӵ5=�L����I^��}�
��@ZB�V<�����/\�E�k�et:���&8v˖U�=��E�oƑ�ݧ��3����%�/�{'ᓷ���=�Q$� K%�`�B��{�=�	���7}�ʘ��6�������rn�{�=���p����-������3m��X�&����ʲI>�}����Mș؊�����Gߚ�oL��lhv�]N[O��Ӫ�S�m1`VT��]��Tu]Чj#���R�
eP�@�:�.�UM�/�a]�p�a��*D�kib�{���Oً��>����4�3��D��W����=D&d�S�6�M����}��?�u�ߠa6 6F��q��	U����P:=z��?�ݶGw[��EM�B\	 %t2/�����E������)P�����y���B�[PI��[���L\�Ob�U�t�i���م�7�l9��@Q�D����e��0yҔ"�P�ُ�)����MB"�Kr��0[���L�㠫�}�  ��J��^bS�*q]����IVP�R�Y"�k7W&9����6ݟ!�����%oJM�e{{_X�� �Z���q���=�H&W���|��HK{ԇ�~����}�8�d�c�K�ʿn���БY>�v���w�J~˄y/����/���%�����3ߑ&�e����>o�w�e?�fe%{�B|B�-�d���d�/M�ԾS(���#��UF"|����VԵڜa�FB 䇁�i�D/x�O�=�����W<9&��Xw8���*���2if�������Щ�<�+",�������[CX�����G�Rj�o�g���Gx���9%]t#���É�x��ي{�ց�%����~*EW4��"O�R��j���@��'^�o�}���]%�͕ib<Ft�u��f�s=���</gܥ
�����#}��<��y�[�M%Z�R�"�4����v����~#��u��rH��L 79�eZ��÷X>H�Mrb��t���$>}��K��7�-{�`�O���*8R��,��WG����-��J��g�>3"�<�	 л%�dS����D�Hc?���%�F�u*�9Gﾑs6M1;��W%
��ʳPְ��1���
${ҕ���p!�'�p��E~��o?55dm�6�x��a�1�)*�LV~��$�WaP_f�K+��|���.^$z4�4�}�>�gK�f(�<�hb��Z��G,�a˭�9@ ��j�o0?�zD������G��1���*.F�4Z����;z�5�ރTK5�?ke�&���w��BU��c5��k�uV����kLyV<OS��÷�uD�x�E�=u&�3�]d�1 �����-ނ�#ַ�:E?o�d�fg�(���s�ފ2k�����k��H0��C����'#+%�Y�O�I�ݴu��cj��)K�3m�Q�`-SËX)�2|��,�&EZ��''����):���p�ftY��O���w0M�(�:	ov�J��U�&�R�d	�:݆��%�/��))�X$��9WM�Qt��-O謂4;8�#�q��*�� ���ʤȣ�x��'l�a��4����OM<� 3��e@�R�(��@��Zr��O t��b��0���Hu,�һ�`��6�<>;�m�>�����}���qa�-�Nze�LU�2ؖk�I��I�����`�L6�Am���%
4����'=��Sd�;�j�~�r��?�B=�M&E
�A�ꅹ�=&�S0��9���W�F�1��
�)O/��o� Q��}�u�D��E�Km�E�*lM�2},sO�t(�j�:-k&
�2��v�oX���v�c�"�Bw:��w�b�(�"Ӱ��:�/��.gF�σT���6��	�\Nĳ���M�6��?�[I�%P��_�j3h釃*��v�H�{���S�~rO����i=��7v�M}��4�2pOiuR��k=H��������-ɼ�;[QHg'.=�i�Ê��Gk��g��'('>�_�9Jc�= �6U���	S|�DGW�q�:����>r=(�`�٢�r�i���j��r�|��\�y�M����b/R�~����:���Y&�#��\��\Wҍ�7ER@ȘwH���G���hX�]����f��$�aȦ�A��k�P���3謾ب+�]�-6*S�B���
��ryݭ�����vz
���h%�;��4F	E���Hl
kF�I��+s֪X�'"ڐ2قD�8���@�<�f��E��k)#Us��D�,�����KL&���^Π���k����������DV��r�>,f���p�<#�A������T���eǝ�m�LJ�g|�_c�\c/��徉�k��ӽ>x&]Ѷ��&��էYd$�9x���1ҷz����.A�_��&~b��c����΋��G����4�Q�;�$пz��HE�˷m�z\�t�g����?�7(C6�kK��_>ʹ�k���!�}�4GԄ��(6o9��DIU��k�4�E�8��rl���t��D��-,Р���ـK_PQ"�*��ƓTZ0-�i� ��qL��`��|��Z[��3�����
�
���}R��Tƶ�Fy\�Y����?�2���m*ɡ�[1�|���v�>�C�w\@�ln�q����潜���եGI������QM�H��2O�ysjJ�3��P/�PH�-U����d��w�^���E	��hκ�u��q��~F#5&��{.�����[\/�� ֽ�����Cs��[i�[�2Xj���7Mn��|�}�$X�+��LLz�&���	ov(G�(�ƕ�k��"XՆɠZ�o#Q7s�=��KZ_uBm�7�����SEϳECͿ<G�O�il�/dC`?��kYo8Id��*�2�%\-���δ���=s�<�^#i��jfC6�.���z3�7��8�|�{�a|&T/�P�z���(��?K��z��(���W|�������1���S��'	cy>�B�i�/a��Z��y�-}���e�C��f��B���{���<U[�*�y�����<� !�C�2�^l��-�4���I}gۢ'�(b`��d�)�d��ƲT�]p5�u��M��2�����/��}�=t=���g1�-�Z�@����*/���彆��_��z�5��$0H\J��*��"�ݽ���g�!BF�~/�GC���`�Kw��W����H��4g�<���v��]�d�ճ����E�1r��,�!n�L����PS+�0�w8���BJ��� ��Ӑ�0T�)b���5�6�;*�q�l~�
J��K������"Y��w�#�iш�z<��I�d�\Ҳ�0������(�K���
�������)&d$�_E�?-+�v�Rӏ"����uc��_�ǋ�'i.�2�ݺ\M�06e�&�h�������_9�]H�S@`6��cN�$qX��h�,��;��
�����=D���^��|n�8Ku̐�;�6Qt;�Y���
�D�4��c��h�q�g��"�o��Q��w�Ur�7�
�q��{��7�@aq�	4LQ���B	�$���Wi�B&�v�c^N�Z�w�lDf�[�ɛ]�ޤ�3��ƻ7U@J�[�/��Aut�9�'�����4
��W�bg�/ xѻ/Q��465��թ�坪�і�P�gf@�s!��0}4K���Y
B����#T��l�E��_�e���*����pR����H�D6�P�f��9�=��1��~Ka�߳C�����qZl�U�5�� �fa�*#G��b9�ɫB��P��/�q�wƥ@����/_��-uöCe:��`�r� ���Ԛh��療x�HE2_p��4!I��3��V�4�ïg�c�F0CVY������ȕw#��\%k�6�DW�����g��>�~���b�.I]���ϊ)�G�n��&C�?��䉻��H���aV�v����lg�c9M�� g���SՓ~�L߀�,؇WH18��Ƶ'�.e�?t�ְϰ'�'G�52�5�=N���������{��Q�t%�����>z#��@쬴Z _ɗw�������j\�'Wt�6A���-��{�29�uh4�I�,s��&��@��P�>9A(�M0��V�Ғ�sf6l,Kx:$�xV�.ό���@+��n՛��B?���{��a/���e*����w�j���ߜ�<�l���f�e�.�ջAuWb��T�$M$���G��Իg��~#tmf�!&6	�VQU5���^�z�s�M(���O��JH�x�^��u�̇�bǜ���R���9-�|�@v�u�ß��yI��S�£����^�b���t�Ir����Ü}L;A���@��{�d!?c�T��\â:5��3�?E�=X7�J�"��6�J��m��&����Qd,b�6�t�2,�3�`�Ɩ�������IVz|oջ��tZ#$��G���Ж�T�U}��~7�?��q�L�8������d���w�vN�~��<�r)�\�~�`~'��ZnP��i��硔�AV����R�ыL�)x�!��	U�N*b;T��u����<1�B=��*՜4dX�=t5�D�D�j�������m6:�'QI�j��2���;�+։I���3j�x���Պ�L�G|���Wq�%�-�keCP4��[��o�xQG��0��8c
k�yb9J�G�q�H*���QςB��j܆�Ewh����K�\_�I����A׀��O���$����b����?;NN��*�[�G�K�����+8I9Dդ��p�&�(���gWr׶���/������K�p��!��y>�x�Bq{8R�	l.��&����������]����K��R�h	��U=T\����8i�i�!,ۜ�Z�#MzP�xf$�!N�^ə+�e{$W}ov�x���7_������7�4]"R b�Oo0���8R�M�v?��m/	�{�����]u\٫Bv[��C���&Z�ӄ��!������Bc���X��c
�����r�с@M�%`����+��L��"$l@���"���ٵ���fGur�aRX�#��k�K��חn�y�d�6OK���3�%'�bk�~im2��u�ғc���$���� ��Kz�*~�e�*K���8��oImOh��m�a��̞�R��]ZL����y�\spՓ;)ǹ�p�
Nb��|သ���m⧑�&��I���k�9d�X�@ͮ��$�說Q�&XF����=�E!����=r�Ήy�_A���I�xh?���:Ԧǈ3�A,Y&z�/��񳞇�:��mjJ'�"I*q�}�V:��mOn��8�z��h��@m��~7������;�"�N#�h�炖��.��,��Ꮠ3	���8��^�O�X3�{=.77U�������U�G�J�]�D}Jac�M��֢kV]O
m���l��+������~:G���HS����sj�vT"䈓	��{����GȖl���&���d3����<I��{,'��W��"*�IA�D�����U�!ڗ ��B��A�r6�M��/��,�$��x�!�n���O9�y�!�`��� �-e9�׫�l���)cT���� �gPB6��x����ã��8w���14�?Y��?�������UTG�8��
�����V�<�/��KS����wt?�n�wi6��t������i���D{H.�yh� +1%ȹ��wC�/r�@�f�j
�t�wcXXJ}>RX�)�OGX9u,/���n��8����s�`�O���B�%a����xʈ��E8�`�-�p?8�?"x���LόV�Ĝ �bP��&�:��|H�ǜ���Iߓ!��xE�@��q�^yA�=�wE�~����0U�h�.A��Tp�H����K��a��
����z�����*�v�|]�����樠���ߏEL��dV%�.e����=��b�����l��|"kE��S�N8v���H�<�Eͱָt��B",ka�6���
�� ��A:�j6�C�n�)�I˳�K�I�@�~��V>5Z�_��ߒE`�D#M�#��4�v#z$|s�F&b�cv3���2�9�\X�l!`�����ۚ�n����Oee����x�Z}��Yni�y�l!~���÷�gW��UM�?9 5��O���}������\?�\�?ih�}�đ���'�G�"��Pp�g��BR#���>_����y��������U�ų�BE�h��i��nc�*9P�tўE�OnE�E_}i��V+�][XK��2�X't�bI:���'��
X�/��2�Vm0c���.W�U���h��5�L�R����F�bc�@~*Ϊ0��n��u�5�"T�M�� ��N��T���ٞu
�h�֍�܉�U8�޴qTF� ���7AY*��W����	h\KV�|��&ס���%gt�+��o�au5���V���;,N�&r�6Wp9)@I�Mr�&6'E�	!��U���Es2���"����TScf2k�<:5S#s#9M$da�w?~Nn��u}z��{���|��oq4@�c��Q8H����B�pa�5�5/�	�U>�&��B{�Z�P�~vG#�37K	�J\`i����=�#ard��5vb
���o[D�	E��)3`~/��_]Z�0"E�>dDj,�fB�.��5�[Ġ�OS@z�Ѱ%rs\����<�V##����<�c,����S�����T�D?��c���l< �R��~�q,��n�����H��-� �,��%�&"]���v�����7)���|!�ݷ�+�s"I�roзJ2�7&���G}8���W>��e+0.`R��M*�٦�@�=B��*Y4(�U��RUҒA٠���g�a�u
��7\� �"J~���o�otQT|�A�y˯�m"_����e��ˌ��;Mܪx��ץ~.L�g:s�V��9j��/����1����� e��/_\+�����Nj�*-�<��ΒI�8�a��g��|�5���٢^�ܡ��E��DR`*(�t'd�Q�8�$��q�-��}���C�����?-�g=�-��Y���o�����9�N#=/�l˧�����^�0EEh������#>Ob�@ԯ1�J?��ۂ[iھP��zW0�)���Y~�xjxx���g�ľd�n���t�4;u�'���p��2։ֳ}�K��� ��!r��ZB��|e�'01s ��߶I]݇JK':��3_�*i�,�^[�g���\�G9[�gL=��Q�ќ6o|�aP����t��&��հ]��j*��ݽP����L�z���#�4#�b����J:��`_��ήY vE7�8i}��y_W�4�]�6�)�2��t�RF
-�� ��Ӧ��6�X2����>�=u�G ,�;;P���"�F��>����TFo��9����u���I��J�rl��k7]�)����IfD�WD��E.����8��3q>jBi*:� F�h�{�k�4K��R��mC=Ʊq�::�-��m9�ӣ�2��o�Kқ(u%��̞�0v�hh�]r|����a�u� ���� �'��sg�G-�k�y�թ�)��ݭ�Dw�8jJa��됨^e��X�ĝ���At�Ϩ`���.%�A�J�-1��x�z��B�����oO�q1YYs"�%d���&ܒ��H�٢'�������S˧��x<��h�뫑��ђҴ����>~m��O=aS��f�M	��~�W&֨��?��������	9�U�[ ��]d\�9}=��V
]%H�6m����-U��}gCx�����Z"c�����~U��QQjn��������d��W0�}l��~�iɵ�����G�y
�4�񀚩�9�+%��;9Dk.h�D� B=q��1��R"���x�u���\�ȸƖ��%��S6�j���g����v�X6���5�B����s"�ǹ�ɑ�7��3؉~r���s��۰!�׵�CUB���>�K
V��cva���?����5�3���ۄ�/�ir�=�/�x�M*rR'�\�q���}�pӂK��x=��u���C�md�H�דuu3Z��(E*EL5u߫b�ql��4y�pS���UZJ�=�UCDJ��c��uU���'�/������;�m��5�v����Q�	-���'A�,A�۶��Z����dټ��� ��⽐/�����e�yDb�kg,�9�*�b�w��qԋ�C�ꦭxg}+7�Z�Z�dg�A���/��gJ
0���H`N�+��+!KO���ӟB;�n0b�O��6��g45��7�~�/ۦF���6�&��,�ˠ��65k�4Y�_ˢ�ꐨq��l�owP�$p�zk�P��E3Q��g7z�ya��dk#~~���"L ׾v���������<��Rt��|�"��qU)U휄 k��W��e�C.߼�Zs��|g@&��QI��U{	������y��"����Q�x.I�spl��h�~��(?l�:�Q��n�V�y��쩣ɼ]E�^>�P*K�I��hI�N��$t-��I���6w�]��Oy�$��ˍ��E�!8&q��4���F8�j#�has�y��V�ۓ�X��`ܳ�&��.�����D)!���]AX]�Q�{�����)7�8)�*��2��s��A��{����Mǆ����@�:w��e�f[�Y��@� L��@<k�H��}��L�x�E����C�����f�E��c@QM���- �v�Z��'��,;��9?ˏ��!T�=y<��@?�^�/�,?Vgc��B��xx;�=����=~���	�搯� -�h߁ѩ)��RK~�-�?�y�9[XJ��gb^w �hvd���~��Ԧp+� �nL���%Z]�a}��|'2��R�zc��6�3X�@��_���}+x�"�f'z��F��p�A:�#Q2��.�:�v{�h{�qfet#)�st$-�������4��k^K��^�t�d-�'�{���p�q׀h�;�+b��>�$�sݐ���Q���V7�`����m���5R
�@>AR\��g�SXi����� ����r�0�"QKl����OO�|�{D�h�6oD/�{n�~&��]�?+E�5���T���6�Cbg��r]V���o� \�ݑ�{�k-�����ݻQ�S)�]M@���8뢄�W]�P�J�oa O��袍/VV)T_����%}CE�q�j6��!���V��d{�*����Δ�.�\s���Qf�m^W�+n��Ų����Qo��fS*���/y��[�M��.�^<k�:�c�|x�%g������+��\w��I��)�!�*�XGm��p�7z
�0N����*�<�����ke��<$]=���S`�C��y9��·�)��g�%��ܐ��=�n��`xpV�� �?)�&���ᠭ���}�#�~.�'��	5׿��u{��(�CLJy6y��m�ȜT�'�7jx}��Hk���pk��j��C�O�v��{��A3/��Aaj7���R|#'�Sg[d�/�-�/}l����~IS|�%��,N�q�,��,��l�?}l.����g��%Zrm��o�获�0������
�bw��VL�H��EK۷򩘮�P'�����Z��?M������2�U8I���]�k2�$Z�w	/_���aIN���R�n-3�����-u��=�`�J�:���m>��#ZQA�.��_�W-����;G�4X+B���ND��Q Q\[	�$L�:d��ֺ9̼����\���-n9ب�U�k�r�r�*�A`���YX��S�#5�~���[����/�AY'�m\wh�bϜ��,�
 �C���
T��]A������h���F��t������X�Eݰ�l���Vm'-�)ٕ�m�unE1���V���ޅ�]RQ�O�\u8����U?��o
9?�ėQ�:�YY����_aD'y��%�ˑRjU�������Y��\�g <y��̮<�X����#L�B#���.�쥿P��c	z�K���ӵ'$������Z�?aZ3���y�h?�ڛ�N?(��]V�r���M:��6�����q�F���|��=��k
>-�nGt���u�>#�3=.Fs�U��1٘�ޥ	1Y�52/C^���Y��q�s�:�� h�/H5a�/�6N}YSu=O�O�$z�岅[fq��5�4����k��3�8���+x����A^_K	���	���&���+�x���:�:��k�CA^�b��x�"��@P_����L
��΃�o��ȅ��wC�������v*ƗV؟����as��jQ�X��	��8j�i�g�[S���V�uP��2 |_~8UcK2�TN��R�d�FQ�!{6��u��;{e2�K/�*;�.Ayb��W�*��Z��
R�ն|�BQq������v]�v�؟e��Om9�����I.��V��mǿ��3�o��ͷJ��R�ngy�tg�j#{��{l�������u(2A(L�x���r��#��I0�;��8�}c�!&�����P9N'�z�J�r�.`����'l!Oo�1���j
�����PTp:}9wnW�������"R���gb|�BeW��}����a5����P���1���	�"� jhdce�G��ZeB��� 	x�OI�kH�v���o ��R[l�2�X;�Q�?��)}���Ԁ�.m�jŠ��7e+�3R�T��V�F�V]O{�u�E�+��0����)P�A��OQ��	�6vƅ��_��|�ϝe#5!Ix�� ������/����xM�_��:�HM)Wy��z��{���w�Q�����E���X���8O�N�ȹ$I�"�3 _%��o-�H�R?����"�@_�5��	"0kB>ԯֺ�zYc���崙"$�M/�RIM
'`�zֱ���� �=}g�u1��`�GEBq>Qѽ杕�t]4 |��xXT��v)�o��`�4���'j��`)O>��ܤO�~~��/���N��Qv��4�����s���2���7��c��b��
��F]�\�I"�h�������d��PAR��U�
�� �����~�g*TJ D\2:@��xg���0r� �!&�yi�����7ϰo��H��#,d������2�K��U�1J�s�Z�i"�h,�,�j�P�K��/L?�+�QS"hB��H�4�\��x��/�@ί�m�V����~��jq�lrj�>P���>�4i��b�]�*��h<�L�u���H�a2�����~���,�s�� o� R����oz����7�Z�Q�I�#����F���n���b��ě�jR�����-N,�8�ݴ��3ߕ
;�6����egL/��%�y����?�����W���ȽX٫E��U=��=�)�)�b�.gDV�LfR���<�$�a�����U�͸��r�R�־������<ҁ��N3oA��?���7�gG6��r�_?:e�/��8r&pbqV��t�7�[PaS�n/Y�~��Ly�����ו�7�cx!s�����b�>�î�2���q�����y �-���J��^���4�U�A�O��HOQa,\? �>�n���,�QJ.T�J���$���帍�����tiΊT-Q����i
<~�*gP��XՋ 2���Z���`;�%�9;��7������.`�/�D���݋Gv��i+i����셸��Eј��*�|�mu =���}��z��F�
aiG��]2Ov��5�\C��K�z�IP��Dnot+�LKP�I	ǃ�\�´��t��؂1Gm���׈���;vi�Vؓ��1��هCBa?B����k�O�nᏓ�3�6X�8���_�l���8��"i�?����q@�XE�c������|�pS
ڴE��&��cv�6P�l�l��a�}-I�I>WI�c���3�X�$5�5 f�RA,��q�U2�;,|�����Wwmx	�i���jc��u�|�N<J�l������}i�]�2�3��ء�Xǎx:&u0��0�FUt���MC4�	��:� �rp��F���1~2�{��|��A��K���tL���̘�����#9PѰT���ў�}R��&&��C-oq�ˌ/�"U�ϟcʲ�������"��>�MR�c+c#e���^�Ѷ���	�+��o�.hmjt5�#�ީ��ό��N�j	s&|���$Z�����74S�o'�)&H�?��'����t�p�(�@���_[#��:[�����Ј�D�m�aE���s�L�W��U�̀��/�͔Q�3����{wˆhok9}�3�]s���r�qI���%{�o��f�^6+�l1������S��4�i�O�z[�����hAm��.Lt,�M��bPi�_惇��U���ev��#6�L��j�Qe�h	w���[6��	�H R��!U2�Y�Qk�ύ�L�#(
��L�ڳ���za�,:,����M�ĻY�KRơ�O��3ʇ5'ҙ���ꝭ��q\���P����{mਲ���St���d��,�a�x@3�*g�n�O$4ݺ�̙6��$\
Ut	����X���,��wQ�Ha��QX�O*;�*����f�h��O�L�S��@����=�2�����M����?�hV_D��ہ�8�g6���_���}�S�<����AFX�17���@�6�e[�����[��Þ�P��n_m�h7��3��!���r��ϗ6g�h%����em	I#
5�.�^�g�, "�~N�4�7q]":�W��]X�?q��?� �_�>k��8y��XQ`Ҫg�ѻp�rnр`
h�[R�@�-[��3Ǘ1�F��\��fK����q0E$Y���9�(Q��A�V��*1�E���>o.�ʃ
U�,A(�r���9 ىY|����J��� w�`ζ�͞�Q�� 3����忌13���:���H��S��?_���j�`m1,�|<9|��Լ�D����z�W�������^t�$���H�^�qE�"յ�X��y�0�}		���i��R�w�򇁓�ܟ`��H����@�o�|�'��̈́��Ee��͍��W�v��d7��� B?��/ע����:�7c��] ���f�	2H*+�m�̾�:��5�`�*��Eij�㐩��A�t�D�o�st��-��D9�uI,�a���4���*��'Ӧk��'���U��HD�x-1��'�J����Z8kځj�s���H�
����f߽�.u�@��[]����6�c�c��Ƕ�=��.�Z�E�K�P��)rin�l�����&0���$D�r���D'�$H���O����d�s�.r �å�B��ө,m��*a��K��57!�_�U`?`R����d�J��&����
�7��?��.�+�|��
r��r��ld^��6+ף# ����u{A4�U��fٟ��)&��p�5j��@s�g��� E��m#̂đ��tv�
�P|�ؔ�T-;�+ м���مqD{{%b�3��0Nː��^~U�c۬�! � �yG���!KaK�iN��o@�g�&*�S;m��ҋv���@W�&�ncQ��Q�2\����p�<�M��[��.$��H ]�]�@���n<����e/X�h.���������J�8
R>���t�&�@����b�$���n�����J�����ۛ����b����="Lx�Ah5��?�iίR/+6 /Ȧ�k���F��L����ݵ�R0s}����W'�e�֮;��-t�6�`J�_���('��k�S��P���)\�5�l?I���(�5x�����< cނ�S�{c1x/�o{>�qO/b���(._�5/��j�Y;S��|S�<���|���ѷ�:rlk/c=�vp�v�c��`{V\����=��\K2b=)
w�G��u����8V%Z|��2�����N7G��VtjP��&�fG<Q��4=c�ķs\�h�_0��梍���k����2�JԘ3i��x�(�F^�u晰,Ԇ��/�I�|��N���4�Q��������Hx�����ސ_���@��r�9��&O-����#��?~���q�A
�\@O�I����������3Jg,��L�o�������)r�>���F�X�ydצ>�c�Gm�	-(�RZsN�z�=�ã�׮H�� �:�#O��2�Q��.��+�VI�� �'�uR��S�V��!���D�����>�,�=���ӂ�����O>�LbIR�2�M�6�c�"�PG���'��=]�+p"fz�P�]�-􎖝�W�5��!-��w�z����!�?�Rh	D�D�:��>e�{���3��g[ʄk�(hG�%��#�G�W�8wѿl�c�Va���mu2�EzV�����^�
A�*?�$B�u}�+{��s��^}-8�%��_����O��ʬ��Z�d��v��{�%���s��i��z�{v�+d�@��S8��#��\�^bf.c>�$��J_����BC�Q�Ǒ����K47�`I���(qZ�����ܢ�-�|�DZ"� �,Qe
$�^L���sL>R5��gdR֧9v�ZΥ��R- ����(07~N�#X�|�~<�	JlA�$o�$�ذnֲ��gZQ�Y&T<�z}B��zK7��X[9�j��y���������	1��ky��\�*ka�k���iy{�-�����ǎ�w��C��Ϲ� O�-v���^lY�c'��a\˪
BI���K��`T���l�v�2��Ǡ�e���"A��v߃p�#�O��
D�藮��)>��2|�8<�0X�q�	W7`k�

�%����_�&<_�t<��h�;^t��UC��\��G�Є
)�Lc֧!�4~�yv����p�IK!O�CK�U����}[��H���;"��G��YK3��h;�j�e���@T���ؑ���|jSb+]&��?�~(���D���H�w�jR�������WL��Ԧ ��;��&b�)g�bBH{��b�˃	ll��zo4Hb�7X%�H�$v,M:�h�H<k�h��s��k73��}�����X:\��B���4�-�Vh���x,�Ȅb���ďY�8,�Q�T�H� x�Q�q�?d*G�S�`�������0`�ާ�%��J�����]#���@��1��o�P�VWn]�u6�Z���X�ݒF��#)���з&��Q5����<4�}'��5�_=9�O�_���ǈ�ݺ�χ���u������-!\��Z&57��.�
�9-D��s��7,�Wo����}�!��YAA�>Z�x����o;�I������}��xnm+\k_�� �:���[S�z��r�`ѐt�á��b�J^tN�u4�a�-F�,3�e�Əx+{�RI��Z�q~�!)����y�_�
������8��v}��/�Ϗh�S���NwA%���#7�3qo�YCr����o6����'�L56�_��_��o@�,.�b��xn�SaP�y#
�[�i9��F( n1O��"�%��A{F&t��+���!S���x�<o��Wޡ�N�S���,}�_L�?:L���ڕfŶ�M=H�Ƥ�"м�x���a
�0%�$0[���_���4����T�p�U���)'M���}�`n8��)]���|)}�d��WR���c`�ê������ػB�Ywܱ�6P���@5x�3I�/{o�i@�G{��mNh��.�v���n%k��ĵI(� [h�f'3:6_K �D��,�qQ��B��C�#=VN�d,ʜ��}ʒxЗ��eF�N�[����^��;>g���%�e�����`�ϝW��� C��2�v�=R..c��3�Ǿ8���y�=|?-K�Q���ȹ6X� ���{�N��3=Ƞ��L�\�������N�[`Y�[�t�`�2;�@RQ��W���@����Љ���GS�M�,A�_�b�4c�+��?���k�ftܕ��N6�Mc .�3'��?���V��܁X����ʣȔH'+�)�B���͍r&��#��P���^��R�p��M�	��I��U����X���Ύ>0�R��d/t���d�"+-�[�E9 �<�CݽT1-��ChQ��)ƕ�5Q's�\)�����mt����)'%�v��4@j}?H�qt��ބ<l3|��N��ޙ��){?�v:�[	�>�f�^p�~��2Q��1��Z����/w�}Ί�e%T�A���{"C���8rQ����u���WM���s@`/����'$�oS)t���&��;3(�M���ك�qs��5h^%h��P@G����9*�x�j�� ��ÄIP���I�T�E;Xd��i��������K��'���ߗ��`>�S�!�(�N�d3��}/Ȳ^rd%Y�ݥ���Nc�2ՅK�*�����IF,η�SgB��~2נ ��N0�o��ڬyn��5b��,e�~�d����7�Y!<*��KDK	ņ)�q�V ���#�A*�����lpVi�����~�%�\�h��e&7��t>&P7�_��b�)?����~/�kg��I;��!/#$OكRj�V��x�N�́"(P��Df�b��5N*��%�ɳ���'���3)��Xf��^�����Z��m�J�Sn�㬾j�(����7/��kD#Pz�,o4Y8��N�R�Vfn���y�4ር'��˫P��eo��z��!] �أp���&д�zǿ�B� �i���|�Q(�Ë�����!\(0Ef�����y�2�wц��k����}����C~�����2�%�i�酥e��2�1�PD�U�(j1M�r�Q�{���߲Z��_Vo�E��z�Z&l�BϮn�a���؍9mLO�(�u��h��7_P�0���̬9�����G����s��I�[;U�Dm�"X�`	����)DjH[o���0mƁ�
�!T��1����k�.A,����=�Z�F��cu��]���j��wwq���ӄ�qB}K�c��ӧ�e
�7���BŊ /�읕���i��v��ڡ<���^h�2Q�4&����t/5�A}���`d���)TA�ņ#��@��2��&I��Z����F˞eDnb:ggv�Dߵ��p+KW���\�N9����{�uX
Nl���	[�7Oת>j�B!��K�bpgdq��Ь?�[���U��$�quf��(�7�(�?�1Ƣ���:�\A�!:m�aze��d�K��"Y���������Q�'_%���癪�A�ʑ�ª���Ā"L��PU�y�t��O��!��'⎮��~��0��*���8uF�Ե3!� `�00!M�9��|�bI�єX���X�Ֆ)o��{q�3�LT�ht�>�?�4lk�osc`�9�&ٶ@�p������)�et���Tgc��
%�[�ڇ�3�]PE� l�F���� �)E��+�g
DJ�뒖�΁�a���@�+��Qō__�n�$���1
0�.Ֆ׷�1�dϵ���l��{B��oH�0ߕN�cW��B>|W�S�NT*�q��X=`��d6;�,��͙�\�������GOQ*�v���e���t7������,L�eh7�w�'-.?��I�y7�R�l6�4WU"�/F5�T��JĞ(��a��O�6�O��MS�N�$��NFg7���G��=�XN�ϤⳢ���6a.�R-�����[ȯX<�/��
������A��4�/�~$T�⅖Q-�LAɌt8G���@�xH�I_���L��RLt��6?"j�X�7CG�T��3���@����Q��7z��;9�ʆ�������K�b��zrը����z�� �<�["���قLO��v]T-l�������@�*f�U*i �:)��Mp,�徬����
��=�;ǁH�ll"�S���a9Ί4�|I���+ͧ'�4/,��p$j�=��bHoy��~!�/1k^��A����M�k��[>��h�����,:~�@�tZ�G7)ެ�a3����Y:7��Ž��3uW�if=xI�Gcڌ>�듉G�m��?���tGa��>��at�`�//:
XBr[I�p{^Dr,_fo{k�%ב�vd��� H���5=��E�X{���Q�y��h������\I<	f�@y	L��Q��3ݢL���'���f��%���Q�ܶߎ8t�ɜb��_�	_�JV<CQ�"�^�xa�z��ՠ8޾�2�ˤV���9��X����^��'��ق�W��ly�	���b=�L���a� ��y)�$���|=�c��,�y��oT�O���/0�z��.:}�Gw�DNjO���Vۅ����G�)L�X���.� ��-Oe�S��j��m�'��w:��6��~Ѧ*���g(J��/cK�N�X3�B�!���A2��p���_Q���z�#�#_.Ι�K춑���?�u�kNa���^.eD�)�8q2T:�W�I�``��rg_���b:�[)�|�:6������&v���Z����/��2*^���b?F��/�2V��6���{�|�M��u���P���x����9!�s��}ݹ:�|�Rۼl��P��	��o�ef�i�� �o]��Z�Fɇg����#���yT�Y�$X�S~����Ғ$z y���-�Ȳ���%a��8�\�H��'[t�M�Q�3�s�����ђ��U�� '~��Dd e��`�^_B�o2JOA��V3����SH@v����w��D�wp��v[�)r�J� /��T^Ѝ����t;��{-���&�j~�N��������ؑu���a��5 8:݃~���η�ST��[p�
;� k�aTďw�-C��{K8K'ȋ�VǱט�'+,��Y؀Cȯ�@*+�S�W�r^��<a�KEt'c�e�?B�������1�4P_	��ow����n�l}'�
[*��s� ��t��DL@�-�g,�'g��D����/�"�1� �y�A0o~��;�|sCD�`
����G��vP�e\��e��A}-Tv!x��%5X5+FcG#����P��l����4�LAv��Ȃ��]�QB��Ba+7���(�a�Y�S��߹'�}|S�$��jc�gJ����.1dr��~;?(�2+ Lw�'���p�S�a*�`���³�I"�Ot� D���/�R�A7�����?�:������^~���/�~'j�jkÊ�1Jt���"��dAl�:�2�-|�=����0H�{��(��n�<El�b>Z��LXc욉#"1me�S�U��G��ܛ����K0h��n�#��V�u&�Ca���W�'i�����L٥��EFV�Nl��%0��aە����{�����V}q_��=X6�F�Ѝ�B��n�z�&�ʔ |���D��+������;�E��9K�	e�_6>�M�@C��px��~7G6�;T��N�J��G[��T�U��O����H�(�.�bNP��?
���E����b�SG�1�.J����B_I�)=�6��0�x�j�=Z�I�^3�6����F�o���AyS]	�]��~Gj@:�z�f"�2p-�*j4��)�
�^��˯�?�&�$���_���7�$��(��&��O;H/U�a�L:��᱇��2������hV/�ei쭅�yrоZ�LRHz��	� �WK���t�����Y����b�����BU[�?�@��e�ݯg�^����3@-Q=����i��Q#(��J�T���2�.�WV��ȅ��n�4�x�����	5�܇�x.&��N5Ydf��8S���^iج��1י<��$���t�W���7������L�µ�P�u�8Q�@p�_b �9
�)�z
g���^�/������ʜ�����zZK�z����`n����� �sb❜RB���5�(��Z��Ιk-�,�o3��<�������!l�y�3kH3�m�Z���ҹ¯u&���m ��VC=p=Z6�ʘ%��BͶf��.�����8g���Dg,^H so�YH��A�2h3������������S��i;}-&��%����9�u��L�f�G0�y4?Oz9���ܯ�"�UXt�5��_*T�Ql�L�Ҹ�$��`)�`:��ag&OA1��	A�~L�ە6�Կ����9^U���;�"#}�� V"N7\$�[�s����!�U�@��sIOH�s�����o��`��A���_�ڋꑁ	��/UX{���^�!o��9�ߗ26>3T#�`ڨ7s����51|+̓`��/3�;��U�ei��8�:Z�%d\�)�3 �N����+��'��x�_h�*�}�.k�F0��\IbuS�w�_�SY*.���"Cy�|uѹ!.N��WW�ĢY現3�1޿m�&F���:u����<c�}l��yLx�p���M�	�WK�蛱��2���{B�>���`w\�-�@�Y��n��E}��am�hO#�-p����E-
���e�V�ǑW��e��w�fR��[R�?aǏ��	�zř�jtC�C0p7~�=��F|�'�=`�.���e��j�)�+-g|��0j[��ϙ7z&䉀g^�k���Qrٴ��+�(��7����{ٲ�_RB�Co ���P!1���&g�X��Vؙa��1��'�LIǉjs������@8w�^�b0��*�O���/��� ��7\�,�nW���uB�2;��N���@��S����[Ǌ��Z���#V����?��D?�l���۬Fakf��:�jQP��)*-��P�*��q�at������s׏�d�$!E���;��圾(�N�H���O�Q6�P[pE���h%��x��d�Y�F��m�y/voq���O~�)xD��Ng2R�����4@L��b�%���۫�"Z)���� �	�`�e� ����M�TĨowFwD�M\zQ�����N%?K���Ob� �;�<�����E�ǡ����_p��Ս�^m�7Y�BL�;���[̆m�Ô�x<���!��6�m=(�}�@A	�b��yk�*
 c�u�@�fR��{�r"+k��^�~6ĄC��_!\�집Q�r�X�z<� �H�B�u#L{�����޿'qšf����Ms�H�q��jM�V;dO���\���.�Y�K��ze��2^4c�]j�����
J��H�VL4=`��V��_q8� �CF�w9���`<睃40�_h�2��>���M�eG�u7�μ����!��5��G/.��䆿H3r\�`��
��M�&$�6�z�Y�8��k)�%~ � .b�%6�н��е�v���~ �'Y���1�(�j�5��r��f��lA��D�і'��2�]m����Lt�%���#Zv�9�p��\����s�X;�B3�
})�fC8�*�����;􈃓�e)�?.'����m������d� ��x�O�O��P���b�ޑ��\���F1�I��&\�{c�:��U��%�Qe���Xw�_7��*�̏@dsλ�'��r^�t:1��R� ?𽭕M���T�[��_�ŧ��>L'����}��Vm�c��6�{*3_ş/BP���}�M�S{��d���O�����!��a�~m2�5I�"�0�/6��[3�lj|��裀xb~w��7��bP��ut�g���>�,��r���&)�f���h�ؾ��*�MY{F?k��jB-�pk��n8% �q��)t�ؤ�O�o����6ii�%����ZuNt�3���'��J|.ʀ̆*�7���]����{A���s�v��p�`�IR̝�m�83�(?Gܤ>>9052����tDS���6��� ܞ~�p�d�'HN��&�>�B��R��]p�".j	�Fv�VK�6�8�:��]�A�}%��C!�m��I9v&�38.lJ*�L�=b@��|$/`2�|1p�����KRyI���ӱf��`�Z_3�kp�K�pF�t=nFbE�w�>o��s�fl9��ɹ��bz�z?�)\i���;�2�W����`���}3�Ir͠p
�c&��65wC�?�c������/B���0� �I�M6��ŤL��I�ڽ ����h���V_*�I
MQ��^�,.���R���	�/���lb����B���bW�Q}�������W�ѿs��_��I�y��$�iB=����q.�x�_&'�(��\�m$��&�2?/�t�-"�,ҫL��9Z
'���LR��(}`�\���
��;T���kU~Ϲ��c)��� ���8���i���N �{��絘1����05Ba�6�.��.�|�g�N��u�L1"�1H �\h)#-��Ԓ�$�h��T��R���B*��4|;;�c��w�G$����R�U�th,׮'��A��}Z]����ɓt���f�v5��-����%=p��p�CT}LJ|�Dv������7H*L5	����'�J^��J"���K��>���&S��z��m��D�N���M}�5 ��ٛ1�����5呪*����$"1����r
� ��M�[T�T�/�2X��2�l����	SO� 	X��2�0��GػWZ�J�w�� JO&�/�Sg�'o���� ���>��1�T��O�֫4s@�����_�-;�l���k8,ČA�I����3o͞�i#����������J8�A�L:�YG]�q���Q�L�륺]�?1^z9�չ�f��ad�?[F�o�j�ʌǲ��?�����s�?7S[�L,�!i����;��k�<&��8��t���R
N�L�K)D�"Ci��������Q���/ f���d�n��c~g��5{ܢ���n�O����P��[����<P���K/iʵy��3��U>�AT��������$$n?ƒ�o�>�P#%kBgX��N �xVf;�R(ZU����#� y/0 <N���tp�-���ݨ�3��R�\n�x�~3���t_ɀ�x��KV�FE�N���ی��f��[a�.lkk���aR���6��ٞ���%���Qb�������>?/�`
4�����&��o�N���5���`�@��R�3,�_��C?T
\T�����w-y%~��� 9	l[�F�b^��9���
df�[+�椑UKF��JS<�o`���ev7�q�@,�����A��Cg��f6�q���~��3o���qE�{G@���F��=h#=XA�5:x�o���*��A����L7ؒ��
��cj�*�8��%vL�� �eg�0 �_��",��0���5�8�XN�v�t(S#5���}ײy[��CJ^/Y�^��Ykf��(؝�JEՏ�T��+S���������I��&e����y�̙�b)#"���[ܰ���Dh¾��<�}�iX��i�w���kO�O�B���ͩ�$�
��B�n��#�<�^���z���Ӗ�&I'��ƛ�9�7� ��=v�9�M�TZŏ��!'���q6Y�k�W��[�rQG8�L��&>%7���Ӱ�Ku��Iͧ�i��*�S��Z����o�_�V�֪jn���O����n�L�]���w�U�)�j���C������`�ɑʞ���	v�iF��a�O��j[Bd���U,���Q��j�$˵����^����E��W$x��;����2l���ˎ�p}���V��	<�����m�t�q>�AD��Kw��Y���=���@���Om���:�(Q-;�g*��ThayP�Z׹��E���6-Vy��ac����>���F[)]#���]�)��,Y��Ga��[YdҸ�  .,�z��t?Ľ�������N�w�]7"�K�/Q�����S�+OX�{�J!�&������kyP��ӣ=�AP����hl����KO�������ZyK�R�t�KJ��X[�� B׾At�Jd��80Q׻^��:&0�:h���_~�0U2��!����$+9Gl։��]�b������*�y��ܒ[��F��dF��9l�K��h�U�~���������\mzKc|�D�q�dE���:_"ԋCZ�Q���{��㌕,�ev��͌�9Њ K2��v9��ZEȭRM��&ۚPT�Va˱G�=$��?�{�g�d�j���l�S���w�f�I('��~!��e�	A�d5/�ڃ��EO ƙ�����!�jݲ)�^Kη 2��I��H�|
�^�c������elѼ�V�� 3X����B��-�8�h`4�!m�;�T��N#F)��^��3�Uk���_q|��a���YLD�m��Ǟ���`!�i1}��w��Yڎ�$��'��Ծ_�S�_ɴG�Pe�y�x�,j�.�!V�:m�A��*6�_�1��ۃ����R�H�ɵ��3���բpv�fD��"=y��̓�cM?+����ڶ$v��Lx�/�3�o�rhC)��4�\�����K�s9z��#���˩�]fq�'��XJ<�ߖ�
j�f�L`��
�蟘�J@]�M+�P�ey�f�(�i�>�0�6{�":�?�؊�ON�9��p�D'Viܠ�M>)T`|Sv{��#�F�3��$3%fvw�t���%�~��9+Ԋ*�v��q:G2�W()�xxL�z�/,lZ�F����o����ͻ�]'��|$k��:y���|>C�n�� �Υ��� �/�gm�B:ܴs����m�G&��3��#%�^o�G�}����� e�)���|*����TR·���r�"j���a���ދ����r�����ЗU���$#S{cP&��M�nLa<`c��3�rW߫�i�;m��j�8��=��fZ�	~�3��=�S-f0�,A�������|p��x6�:l?���W)�6�ͷ���
jp�-C�k�r�ȋ��n�W�(��Ly�J�;�4Fe�?L@ɦT����_��Z2al�Ш�5�y�W�i�I<�EIa�S��p%�e�L��������e9	.����yA�9ۥς�;��� ',���r}3U�V]�\VK��'#�_�h��� f�:�dc��̖R�%��2n�o52�V#Ҝ�@����v��bF�q�����R�b!jZ=�a��^��7Ō������G�1��^9�&��-3�ź�gb:w 7;fh}G1�=����~=m������*h�ڛ�Z�9^�Bb0�,��WP��3Ӎ�.�|������]Q�������#\�g��a��7��ɬ�
�iJ���,~;!���P������i�:�K���y�[��K(����5'H�hZӻ1#����O�d��c�*U���`�
{��⇁�i&M��+�j;�Ѧ�<�	{��_NY�p}_�Fi�<z�������׎�L�'TMI��g�mkê+�N�tX��߭�qLRh�|��[�AT�]l�@�u�-[��|��@8]��X�ۮwI��l="�e0�:74�}��D�m5���H>�?�ɀ��u�%�1��	Hw���r��萆�#���xs��DBA�կ���xA>hz����q#/��j���|4�a�g�i���p�F|>Mg�����傢����;(�['�O׵\jb)��$�25@F�4�i`5�n��۔%t�Ń��Y�K>m��\�����̧�9�$�%�#�G��Ļ�[�5�����3���I�&��O��_1���Q�{N�n0Z��f�HwA1�I*X�]���O���'�V'��ɥRt���ݾB5�˕1��?��r.��t^�G�|���/O�5�P��iP�N"&3���v[Ħ�)��.�����Gj�?����<���S���D%E�7�w�C0�Bys��W���h4��C�&�G,pJM���*g}���9\�<$���[l�{�9*O����N��r�#*�͒i8Z�R�:by 8��VF?i��#MW���Pk�\�Ѕ��:r�d�vrraDd�	q����%8fV�	�!���W�DK�ڕUY�����z�ʡ�[}*2�p��=<k�x�7Lt�`" L��j�s��J� ?_ =�1��Bݖ�ˀT��\$�Eq
ڝ����r��EQP9	pD�'�P�ߋ��������վ@�?�e��hD��C=N�ť/�s�)0RC����*o�nbDa���a��+�S/p���'¦��ަRw��A�^d�3���E��������ݨZ��t�v�`5�����ڗG���L�/����Ry��a Bfj"a�5FHn�yh�ΐ�Op�v�	�@��Op��&)))t1B�VJ�*L>ea�������D�Z�΀�H¯�%��Y�b?6��Y�yk�q.�
�TAg�Y��YA[]V��xG�p#3�nO�I�HiUe�؝`֓�	���E��M #�2��	\!]|~�I&h�~rs�M?���}�����l(U��{�T�%e΂��ݶ|��k��n�	��O����N�V����� C<ʤT�����23�=���D��/����e�Bϩ�b��b6�������<o�� ��=�4���F;9UX���>���js)��*�-�V6_����V��N`�l�d`�+�[,�vv-� q��~�N��]S3�hB�~ݤc�� �Q�ޔ�?��\�T���O���Һ�I��L6�t֝Q�r��TՐP��O���D~��.��k#y�qV�s�����x�qj� �O�{�rKqũ�r#q2�����zR5+�M-�<�؞��b����Rƌ00�ǀ���R��%	q�UN��0�����Tj�S��K��=Ћ����-�5	Ͻ<�Zz挠ޡF��#W% ���0���K9���\_l�=��Rj���ZeC�Z���M��>Os��cT\�vG@dg��f/"Um��K�2ӄ�a���x�{Eu$�Y�aќZ��b&(��
ϹEB�X(S�=��s{ח�݁4z�+YQ������\�*�^��K�H����0�|�	�s��Y����Ԣ>�9x�`��^��
�Ʃ6��V�^$���,	xS�Q���.�\�("�Ư�)���/�+�M2}�B�r�&;xE���G��s���i��4���&�y�j�VC���H� r�$TY6�+h�o\�s~���*��c����������~���5L����Nz+( {�1�2Ҭ��-q+	��vo�����d��\o!Z����p����@�y:�谸gf��A�84�*a��M�
��J�M_��~�u�9��3 ��C�)1hh�����&k�_�t��d+�N@r���ZN��H�'��y��ԉۓ.�c-wqkt�`Z�jN�ւ��������1��'҇M�y#MПXꭝ�<K<8����w_Y�8����+�i�_XI"��t+D;jتM�Z �h"d���-PA��M�i=���E�&R="M���9�����:y����،H�[@&0��K:�shȧ�� )H�#�O Clk�kԴ*)ԥ�45	h�)���r;;���rt���pEx����c���v�m[ ���W \���	'D��-�6������yӒ�Hr�t8~�jY��$��Ӝ��k����&[����3δ-���?�����]���w箆k�`��~� �)�Rb�ɪ�?�[��h�|U�4����b6��6$/��驣с*`W�ѵ�]�$#ˊKb(����c��GB�����uç$R��*�[��g���0�4;���3�56h׼��T`o��$5��ȍ��%�^Y* .C�~1�|c_QQ��2P��g�x���m2Bel�g��\���k��B���1@I{������)��b�>0į��gi��aJ���]5���_,��(��RkhM�*��U,%�щ���z��_�}���0�+&'l���k�����]���u�91��h�&�{�ob_�_��O�� ��N��_���dXs(�`(CV�wЗ���=�k�3K���i���v
R���z�E�&Z+B�w0C�� T4���y��a��B�; ���.b��0I�	o7��@������LXw��K،]���:}�dA{R�
�iB�9�E�l�T�=��4��C=��h��묓���x�V]�E��Zڲ��B�C||VI��x�k$��=��&&/ozn��xz��ֹ�Α�)�)������3�k|U6M+�c��*F�Z��� N�p��x|۫=h�F�ѳ�u%��㥜��s�7��7��?�H�.&��N�^���4�W(ym��4P~N(��e\Lh(�`�N�nRKE�LQH���6!l��������b��b���L���@�Ja���2N��"vSGA�*X��Z��x�*&yd_w/�G�L- K��Z��noS��O�%s��>���j�J���N�뽑��.��y-"e�9e�z�le��h���	O@J�3�G�M�{�8E��&27����[�k��@�bQ���E�N���A>���)O0=��H���y`��KR��K�xO�B���S<X%Q�G�����G���v�*A|�f�r�������LW�F�Y��TkF�/R0�
�
.ױ��Y8۪3�<�y��1~E��q����.�&p�N�0+�c0�ґ�z� ���}� ��G)yl$�.�dY�F��[�n)D(�Xe���f��`��Pq!ς�D��a��~�C/f�j
-
)�z��
:j#�6Ϫ�k�Q������s�^�
=�i�)����+���&��l_���0�����E}n0�lTn��p@��Y�9��x5�1l�~LgQ�Pu��ZZ =�-n�{��w��a�zf��w�ȹR�gB��}=yM��y���$ւ�Y�H�4���n|�[�?\��@�Uuz���N�oKF��<��83�O��`�qgm�Ֆ���{`+�r���6�kO�����liM��g���ZM�tQ�gG��[	C3c��i�=D,�������pu��"b�:�KL�_s����� ��D��,��%o��R������-/i/����n$n;�)��R��#U��PD�~����7w���{�`��B�<٢����1�̐բ0`�������q]6��YoP�g􊫲��ڭS�'v�h�s�,>��EФ
�b����!�������� ��-RqҔ�KE����<zdqS�ᨬ�&�����s1�/��!�z�J�G��}e�?�#E�p=��K��D��b�s�����a[�y>�&NF%Cjl��Z��"h�4�k;w���%3/um�Sg�Yqo��
_��U�Fc�Sql&W~���b����Euo	�����?)�pK胒g�9]>��Ů)[�P<O���O��ܢEl۾��ʾwN�ԛ[���2-i̱�	��DJ����GAKk�6R��F�c��4?^?�!��p�86:~�O|��08���<5�,X����jL	NW/v~��W-��`w����������{��\�,����h�-�C�%�}ר�R"6����9���Rq��N�#������^4���jk�����˛\pN	�ĩ!�8���n�aY�f�=��o�՘<� �U"�+����.�b�ˇڒ��Kཏ$®x�ίq��w�#�����L&��*�J�=Tp~\;� ��)X'8�}�is^=N�z}4]`�1�����^�R=jf(�E�D�r9�Z��lr�4�n� Y���s~:�/���n�p2cA������� ���"�X�YY�A� h܀ɾ��P�WE�EI�`�/}��ǯ�� ��ֺ������v�['�/*ݐ2M�B��a�o�_�<�S���O�)H�Yd���*��ogJa.� ��n�bPh��19$��VF<�ŷ��v��j`����/���h��r�yx�ƒ��~��'?��[�2�At��^ �Tk.ߩ�&>R= ��~���Qwb��sA�~
��X�[�"y~t'�G�&�A������8�Ճ�&K�q�5�T	�A���H�0>����sFnr�d�*�m�5��
�YJZy
3��g�y��i�?
���~�]�q�%_���By��Th|8��3Ënѳ	�%������{;wܵg��Fi�o+xX���"���Ux�	�*� �
�5*���47<Qy�Y�;��\�ggS��!L�6[Y�,l�ɜB/�Ĭ�p�p��;M�KO�⮈�+���+�˞)1ܦ�M�׵��{aQT.�E_�������f�җ��j�����s�оk��g���|�`����]��d�Λ��������&�G|�V�_��SQ>�@�mg���v��L~Oҗ��tR�!]S��w֢��Y�́�x	�ޭ;�3U�����)ÆK��I6�`�~J]?`9	+n[X�lP(k��6R]�ј���j�*��ׯ�W�//�MZӗ���F��"c�2d���(�9D�fV��a��?�C��e��������I������r4'
��d@�SWȳ4�|��/��[.Ȧw��j��{\���G$�^�>��nnκS�Psm��d`��+����|����92)��vN!�CI}o���'J}���xPΫL	����LӆA����(�q'�9�N6���䵞�\nuJ?%��L�X���d���34׉�8 ��?����#f���J�MLu��G6�愀�h����vd�'�J�1���m��v�����X�T0�CV�PU3�̡�5|�R���=���?A������)�/�y]Y5�l,�D������ ����<��NU�~3s��{'gɥ��:%ʹ}��#�e�7��i���%'�����P(n����
��`^�)~˹��<,�ɢQh��	�n��Ҿ�c"Ss-��ԥk�Ȟ�l�(Ў�2x^ƕ��o��]�i7�����U�?0r����YYdN�j��t����,�� QiW����ٌ�6�-0��c��(��:��Xn�CT�@�˟���9-�En=��!��O�jB�m
��ԕK]G�������!|�%��x���N��*�����]َ��9�d��MSGU����h��J86a̒vg�L#M��n`����sŨw��1��}�����A85�淉�a��.!�ì
!Q���ރ���I=U>S�1�.�"}(b��9w;C���5W{+�k1�<�9�8�I1�!n�3L�LҰ*�-����rS���U-)�39�ۃ���	�Qt�$���s�ɏG� ,3�����d�ϗ��Ý�[fT�QU��%��is�K`�l{�5k���Zj�<g�oR�Βi�����b�#����� `�B�u�٧#A%/k�j�I�m�~�.�:�9�ө�=&0�ZAv�2�qi:52�Zs�����J&�zEu�Tl;���^���f��p%Bd�1��ɦ5>4lH��I�]pt�@���'�V� �?y�����1�4�'�6Dq���F���Cðnd{��w�Cw*3�=	۹�#��ۭM��cDm�٠_���g�K���U���8��0��B��#���r��q��������3�a7V�,�l�������_���h-�ǧ�\'l�	����XQ�*ݺ�qAytvo�X��������%t�;08h���W&S,���R��=��3&W������ n�ԃГ�ǱZR�Z���%Ao���q��MKb�������үD�0l�*y{�#�&�e�����@�D�p1�y���_�YPZ,�0��)&\�a�q©�1~H��B"�a�	὞���=	�nYK�������NǤ ORBI���5"��4&�O�ҁ+ٕ����+������4�1�0�T�0�� +���z�P!U�$���TJgv�>�����#�4��T	�����Ή!Q5gDU`i��Q��=[`t�t�s��
M��F��lSY�@Q�ϊ�t+Nj-J ٛ�/�%��xpg
���2�Lѿ��5��aͶ#��k����α*����D6}��J.PϽ^D1ݿKf��1�Y�a��v�-�.��/л�+�?RT���OC}�|8jܝ�� e��f�^���C���Abe�)d�o_���&�o��I�1w"&#_�饆�m��=EEХ�&��ъbϑ߼�ƙ&��3fjN>(iL~k@��U�n��B+p|�+;�!؎o�՚5콟5�����M��L F,jo�mexeI��#&�?����lʩ�m9bsR���#��͸���ߌ��9x�^h��&�V3�U'>ds�-����OL��s�e�9U-}!ߐ��ʏ���#�;ޫ$�3@<XG0߀L����w�F�:v���k�k�E�j��Tڿ��AU�~F�XɢѢ��n�����a��ve�4dF��������Iq�@�9v���;��3��S,}����4���p��V4����v��rw|��	F�~�P1�Լ
��cbK�n�+6R��\._����s�J�ڇ��-�'�[��j��Jb�e�рaa?<{��������O�M��H۱QIGm��6`V��m��=]�m�)N\���bN�b���o���IO�dֵX�ߥ�O\�4-kg�@I�~�e�H6���3{Hd����~|�k����#�S��N�(YS� �c�?����s��t@�WFԒI�Ü���h�h���kTK~���Q�е��v���5��
u�Ex�1��)��G�e��)[Hh��E�a���Y^y�,�>O�*j��Aw��^u�H;�S`�g�ޛnAP���bE�Τ��*��b�H�hV�*Z=h@�c`���\� &����'C�v�����{�=�|gϨo�?�[H���!�rϧ��g	?;���|{j$���*�4�/A�z����Yv�n@_f�f���o�L��@��NF�i�b��c�U	�o�z��؜?y�
�X�7L��?d؃�/�t؏
�E=Ґ�ʠ�P�w}V"@��3�/{Y��о�Ñv��i����-A��|;��p�^	ZCg�i�j�+�A�EBď �h��\7�	X�F���t�F/<�d���or�<r�w�Z?�����r,����+Y9kW�H�ܯ�O-�6���W)��i��=u> 1���#x�Ϗ�N���~\N�+tr���8Y�
cX�|�3���k'5Ж�Yק��BwN��!�ѥ�v�S�F���X��F�SzoP��m�|ᑮڎ�M`��M��Y���.R|�C�*�[�^D����O�~�u,p.���׹BK�/m�'w�x(��o�c�}g���������xfc�uOǩ9��pa�Q�H�t/"5�lF�����ﱳ��E�4��T�=��0��5�4��
\��̇�P&��� ���q`�=�P��9�����B�����wl��I�'�%S�&�U�q�P�w���$cG�A�S�n��1��n��bl9���x��L�U%\hfV������¦of؆ V.�	낒Ya�?��#�g�lh����f������Nr7W�!��8����o4	q�N=Yu�f���s��?�9�#�=rӡ%�mZ*ab��0p��2��,xw�0^���@3q7|=��fQp�l+��U����ƭ�+���3yٕ��sz�Q�~M��43�'(1��ߝ=����pJ;L�j3��N�9~4������z�yD
Ź�w;*-�]��O��u5'(��M���؁]B�N�ijS���۲Â>	hrV���h���^��t��:R,�m�o~Q�PfjN�~r��|�u߬