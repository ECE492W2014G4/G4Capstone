��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|݅o�@
�nI�֛TU�PP.�����+���u�Jf]�ϫ(#��$�r�jO!�Q%y����m����T}�R4�?/䃭0����AU�(�ƾe��������f�7�m��v����of� 6�{�
|)t�]з;�Y7�^��-��f���s|J��/k'�U"�n���Ҳ�`����R!.pT�}c�p��_K�Y��TSY��O��T�TV�8��3����#��f���@��>_��o�}�Pm�gqU:|��n�ʵp�g�ɴ^�BM�ɒ�g�/�\�X����IY|�� ���L��
���E��v�# YJ\�H���]�LH�A�d��Ѣ���*���|������&���%���Q���Fca����hY#�M�f���k�L$���dP���D��6|&"%�F4ަ#�j�#�	2��"9ۍ6Y�L�;"G����	f��4Y�.��=�ܛ�쿬0�L[[WI�ŦQ�i��sD(N��5�Ml�
 }����r�Nf5��@RE ��t=F���������FKj`9�x<����������V��{�����I�� q���FǙ�[p��nA��(bw�B�������=D"�4W��>����kK�Ƶ�|7.�����k�����o����yV�4���o��E΢��rP�n�i����b����U S�K�ɾG��⩵�qɻ�#n%2�z�s��5y�J����* ��<TjD螱�G0o`σ��(��CFȬN�قV5D��><	%8[����������Ϧ�Q9>a(��5�xjDN�B;n�a,�k I���~�r .�U�[�:��wv��*���Nb��-V�vw�'�ь�$�
�ۏ�Ǻ�5պ7�3/P���҅Y�_`��Ƅ��s9�#7��sB��;`՜� ������˃k;���i2�H&nZ����+*L(J�HM�A���ڵƮ�]�s�^�6��Nv��#���$L�~�Ri�S��E�'@lKKBb��H{���z����� �H�$B*�m[0E@s��@�qby}|4K���}Ǚ%:f��H�8�@�:�|��рb��� �?Ϣ��b~��x�#�+T)�9l��67>�[�X�&ojGJ�m�]����)�
�pn7t���Wl+ηj���PbϮ�Q
jg��]�W�d�!�^�)�P�\�ZM#+�7^� QJF����2���^]��Dg�� [���i��4HZ�ZB�8zfm\�]��!���ݜ�o�3p������e���_���r�P��mt?�̪�_��r��y��D/[���!i3Rbդ��;M;�b	�"�<�Sщ�:t���i��a�V����'<���)&�q<��e@%7dPW7Yi������&�!��;l��Kr���O.�}ob$R+��*+�3���+���R�@x���'�%��ŉ��#AM욻�����Ľ�z?��1ӳ��
�v
QC�i���*�O���۽��r��KN���(�ZY����u#?�X���s�?(��~�n���6/�.9�x��턈�BI>�%�Tz)'���ٕɘ��u2 �Ra�U�L�������Fs����
�X���,��1��h�Z�c�q/E{ם��a�����.���A7f����Q��-w�49���M�6V���pZs(��|���R��>���In�<���'�!q[�Xf�J����ĺ<�sL!b��xx	~"���U3�L����X�~M�����I�b50N4Zcm���|\�s�����Vgg�6�k.t��SU[�i�3~�����cR�yq
�CJ���v����D)�����#'�&ť����N9i����,�t��!N���$�
H�2F�:}��8�.��G���KU�i۪v�kw�l�����4�$]��إ�yɪ���=�WZ�RH��Ǐ?��m��of�䄬|�Y^� *O|Ǔv'�& ?�e��16}���	z��6�T�X	0�����0X)H�I���m
�dUd��U�{V��K$��p��z !@�$}2#?s-m[����}�?�>�dY=Ԥ0!���t���(�),�ɦ���@J�9:�;�~.��T��f@F�k��Æ�Y`_��Py;�`��ҏ^�B*U�E�ʇ&�Po�Z���g�U,�-}Bߕv�1�l�0{�Ҧ�̩`�ؙb�z␟�4��nt�wXA�^��4��,nd%KbȨ_��/��awd�(�Kp�����(��X�}�s��Ť�m�X�B��,�4�uw��m���rٶZι �A�KC�C�>U�`�J8]D9Dl'.I(�o��j1Ӭ��o����qc�R�=�(�㐜�F��6y�K��e%M�����ͭ� =i�+��Ԛ�U��A�ͅ(pS!38e��>��&��A��*�ۄ$�gg]���*�K6��˝��β�=�H4��+j�ܘR"pb�
��`������2|��n����V̩�N�h�+�TX��#mJH���|V����7ZB��{�u��"k�k
�mNu|��Ft��뽻��w|+�i2d��J�˓=�^>�"���na N,WJG�K�B"�*o(��x~=��3��ȥx�4�V}HVR���	2�)�!dx,����D��^�3"3� �+O^Att(D��v?�]f�N�b��ˊ�ʘ�3(��~ذ#1U�>�W�i���xg�z\�7^�̝S�|!Jd��kQ�V�ǡ@}�0��z�a�����[�'}�gK1���[*�l�l�=J�ڴ�v�t��%Eoa�Ǡ9�g���럻�T"t�Q�*�\}�D���u�R��n�s;�o�j���[��<�ƻsW}|��ӽ+�KOd�2A'������ `��_�#&�_����K�`��۶.7t�^Rؕ|�%�ό����A�h��wJ�m�K��G=]�n�6�#�<E�@wvQ$�[J�����{���'8�jj�b����Rp�tXX�NT�8bb2l�pR�� ��-���'����dPX������%��ɐ<\_p{L ���f�X�(���Ǿk���ӻ{�L�����"��XK�Z9q�:5�)�I~v�q"x:G��<��c���WҾ��V��C��~�;��`j%=�����Tv�����S3��E�R�~[�7�sF�h���d�$�����9��R����DM�l�gH�t�(�Kr���2��,� �f�Ke*F0H].�Ǭ�[�G\&|\cqK`v*��B��?*sI��0���L�T��g��^��a�<�uQ(!��gۨ`���up�Ÿw�m4�/	��i3-�׽l���f��q�v�.�!Nx��@Nդ���M"x2���P�z��K�:��*�?�$d�H�ֳv����b���~&اN�~��:�ѥ$�@�n�z�g�`����3r���=��(�זf������>ϊ�����x�u���!�9'�i_z
�}=���_P����t.z�I����@ 
�ַ�H�N��������
�D�<ѨeH��M�ea�u��^���n�.Y��C�k��U-,x�G31#j��5D$���bɿ8�i������1ΰ���p@$`��G꣛���o�C�r�¦�j����cdİ�7�Q��߄j2	�x��V6S̭�����5U��@��Qt�8�(;�1R�x�)R^�(n2�{�	�41��@�����!�+E�*Ez�]����=�l���J�R �gۄ�n���w{ŠC�P6��2Ƅ��c�FV���V�12B��k������N�f;�,ղx����,��U�M+�>���1�t~@T����i�U�ʢ=���6Q���͓�'���x
�:E
k��o�����=�m��)�8s�����Y�2&�[��c�.��-��Ю�uKuͰ���Pl�?W��uҫZ��87C�3�#�Ϟ�tJ1o��]�R>D��֮|*��)�φ4������?cbR�$<�<�W��=%�ًRѶ;1I��́Eϑ�O�M�ؒ����ь^;Z��\�T��!R�Q�^N���٤E!�}7_�jΦ�n��s�8hp� �GS��Ȥ�yk�Kp�7^Npح9����j(�N*��#_t�V:��C$k�i�on�N�-di�7�ݥ�·,)
X����s&m�1�i�`�)_��3��x��t�򈥁�P�H�`�99�Sp�y:��6
r_u�l蠥�����q�Ȏ���}]�"��|�U�Rq�Ӽ*�Ƙ5d1fW��� ܦ�DN��{h����V�.��k�����(5��9WJ2B���v��n�e�Z����+¡��aj��2�{K�ǣ�O�:j����'��֩ks���[g|�a��G&���xiQC:���!B�S��-o������v��/ ��V?℩SRH�D\r!����!hMX�>˫���6mA�Z0�?R���HB)��rS,�=�s�.��u��/"��#�1)�ʀ�"��֏��7�mQ��e��q�o�vjva�p��<B���2�
��	T:vxI~� �/�/��*��FJ�T��ɨ@dKQ<o��$fgG����V�W>�<d���`�!����3�
��Q����7R��=�Y��W�b��TN%�f��gkȝ��x�ֈdJh�ǒ��b@+�蝋\����BR��+*N� C�U(��0��)s����Z�S���x��gG�%����'HPI�� �Amq�����9z[����eg JZ��t^Ng{g�C2ěM~N<ө�����`֟, (q�����%�~�']���l\�4	h0�w;�56z� �f@���S*겕���s�8��`g�ō�T��)�����na^R�[2~�P�81�Fɛ�<��A��E�^�E��\�;ϒ���t���_�U^��M�2����]&�ʰL�N���J��m���5�BQ�Ӭd[:R��m���k��Lu����V@��b߽� nX�ss�s�y�5w��A�#rF?'��phF �:�8�|$4_L�Ly_��*�Ǔ`zw��O��X�KD�<�1�-�vq}��zRi�&\������%�0�����/i	S0�Kq�6�\s��a�ė��QHEG� �E�)�XA6��l(�>�ņ�c��*��>-:��J���0��@2T70�ivۖd�ݺ�70���n��r���=`�Z�,�t��,&�K���l<1�����Q����ܛ��5�VB ��/5�=|���K��]��u�I�d���jP&�_���K-�k�$+)�%����k�??���w>}%A�zY+jW{=`�,���J�d�w�7��IW�$#���e���G4n��l�O�SE�ѓ�͛{v.D|k�Zw���!S[�/rdPJ����勬��t�=M[ .&�
�U��F�,6���ِ�]n��w��V��,��4E6* �9Wn��Fx��ƕ�'m	D[l��e|��	O�Y@�i*f���4����wŉ�R������Vq�|�r�̋g5ȉ�q���;bs�X�kg�'vԵ�5b��?`�KJ�}Ps0���-��~jĚMo1m�FY�Zg܋r�1�2�wxĝv����`lƙ��6�%��-sң��E'-�(��Z_��Fe������ŞHFy�V��#|IP��&��˨;���5�@D��E��$��_��&cj�ίԪ�{��d7���3b2F��yI��s��M`OK��Wա	u9F��`qS��_&o��,0��2�n�x)�z8`�������j\ۯ�A7p�Zy�⦉q�"6��_�*�)��H�6⥙x�&�兑�ܘ� �zQ�^y1�?���7��/�E�����dܟ�N�b�~+�nz���e�)l(�;F}�y�m��O��|��t��R?�2��9�����fT7C"{靪>��G<ɋ�&���uz��5*�����*��P�����v�ǥ��VT�����e���A�p֬������h��97�����B4}h����p�C���0bɪ��"��&Yg��5������ C����έH�sk�$J�U+/.d�DN5��V(�a�DOn��vZ�����lם?�f(@ɐ�� �y�g�&�7���*f&fH�_>��\�J��%��?]6�*�gR��?�ć����xFi���!�[?��]b|[e�Y���kfyGjj�+ç�vj�Z=ǽ����ri!
ڍ�x�9��ܚ��Ry�r�����_^,A[tr���JӅ�2ֆ,�k�	��Z��5���&8�������6�T���'������as�ܐ"*�.��aV��!��՚����I�*�y��N��]��pG���w��v2�?7�(�m�_L�2�<؇��*�m^�}4�1�^j��ݰ��GLމP��?byFͱ�)'X�?��tShy�m$s��D�:��x�t{�e$���Ǔٺ9t�8��.���4�v��]F��IhܕM]���c��(+��� ���E]+���Æ��.hGӞ�Aߧ4Nߓ�`?D����At��B���@����G�
�~D����IH�BV��A7q�w�з+���ml�_�;vq�m������w�q�:6�M�*달�9��ӆ�6 �j���8���1�Hox��v����MNP��ݯ����%��y%���NKԊ$~eț:^A:D2��gR��%�RW $�����sX��>���ሌ9�L��:������4�g�?��	V
�7����|��7i 4� ��%xG���'����H���/�Ӏ3�:"�"7�� 8`���6Z=դHtJ|1�|�i��B\p�L;����CP�R��g�E�p�2�c����-�Vie+v�X|�Q�	C�)	�9T�V�c�M�|�f��^|��&Bnf}z�l8��RR������3Hg)����/�й�Ӣ������ɤ��*�k�)tŭX�����-���	T^�3�AJ�ĝ���s��v��	��R-rW�f��j���m�I����SX֗^.Z=Z��"���a#�Ah�s�Q'q*�^N�-_���fy��YB.�O�w0��U�m�HC�GH%z�]�A�	]�5�{��	���pӤ�Rڭb蚉�TY�V�����|�l�����E��nb� �o|V.$#�˻`Кfl�F�4���K"ZS�&qΫΌѰ����/����Q�)�5�]���_���ĳ��S�IB��Go~BY�2��Y	��~9tL� �$���z�,_��m.��/��g�u tipFfߧ<U���1�9��U�%�s[x��(��m��ce����f@��d�XZ����U�n�lRZ)�����!.�xp�TL�Q91-V9:�b� ��,�bybC��=ی¥��N9M�Dj�����^+G�w��֓]�*V���b1�sݧKYZ@����d�졔,�+1��^��T�|��ٟ�6�[��!,/�ým����%�c��vm>��0􅴞���C3��;?��?�|��L[��vH���y9�P�n�i'�+��t?�Vf�j�V��b��c�,J�������0�S��ׯJW�	I1���.z�3CD�BG��>SZHN^H�p�_7��6��+�N��'����w���0wKy>�8��jp|��p��M�ŰH��9UU�%<�&���]�ih*)*���R:<�c��G+E-��xC����~<�q=�T��כ�n�{>�8 eb�����^;̺J�Q�0�Ց�v�E�~�1&�+\ʆ��+&{y@r��˗�m5�&w�����a
׶Clj1N�U'!HExY�����f5����k.{7;�G���՜�����a�éǙs
����C�z�s��c��u��c�|!ԉ�"[&ɸ� ѯӲC �K�#�8�{�%gq|mzYh�s�O/� L�a1ӡU���@�g/���We��(CǱ��p�TY��2$yT @QT!f��i�P�`����:�_C 6�J�J�B��i�{%Ŗ�<�k�|���pR�WOa�cw�cڿ�Y����o"!���>��b:��<$�Ж�?���mw%��
��߫yϝ芐m�u��zn	��rXc9���%QI���toR�4���SF���X�dw�y�yO�}+%�{�eʞ��e���(�H���ћ�,�m䟴�YD��������+0��m���dL��6]$��I?yzW��-�U>Y��F���s).y���ؗ�@{��1umո֧8��vN�p�	�\L�XG��5ө߆X�g���*WZ|�؎?�:�ۀ�-С�eĠ[����n���QW���?��ӣ9j�}�;�
Ń�K�.I��'�;������zG��U"���� ��N��pп��B؊c�<�ї"-A����&i\�y!
��)Ɏٟ����@��h��gR��"3���_vK+ojZ��*�r
�����3}��؉��w9�HL���dA��5 H��Lk2x9��X��(�ɹo�����y�B����¬?����,�=fɫr���0TG�g�b����UC#M�Ɗ�9�=��i+��w��b��ݟG��*4��#��5(YdHe���"ҏp隻4���xIhv'5TD~��v��H��kSV6[NS{�.g��B�6�D�k:%~�2Y}?
��d�I��JBzkGӇ��)���f�@2��pG-�nњ���nz:�b��M���h���	������"�6��a�K[m\&h�E�T�%�$�T0.j+��%�OeM؟{'���t�\5%�+f��)��Dd��n�Г���e����K^R��j4�is��0d��;���u�?2*痧Ȓi䴫�'�%���o��\zl�?!�_��N2��^��AH����'P�T�eK3�O�>��D�ʛ�h���IJ�@E���_b�i�A"R���7����P�)� 6���8�IE�^�q���d��u}�H�AE*���y�
�4�	6��$���ۓ�/�����~��=�$���M-i�0ڮ��E�Sl!,?La�O��]����5��u_�Z�x��6�������$j�.E,�#��|z��p���UMa3�Y�$��t=#�y��n|"v�� D���<5�M�7�&�*fJZ����q�u���:4KF��}�.����PY�k<P�����(�ȨJP���GyoA?��l�V�\u�O%��޹�M��퍻;��N���6!�%�ju��[#Ujd�O��g&-L4t��P����!�[!���A���['U�j3]�F�N�s�\9:���+-�淋���`0�L����j������q(�A��T�R��?	�.���}��6X��㲝
��~�Q�V
#uJᤘ��y��λ�ip���$�"I�Nn���g��tq��P��By�?��1.�K��8`�ҙ�-_��{�O��;�i�Hof���2aL�m�E@t�,�@�;Q�u3�%��47s��ԃ �����<��x`��{��70��^ܢ�����O�0��e��5�p�[�5�J�V2u�ie+Z�&�9��6��W��8ג���>�d&h����d����������f���	�L�bv�?tS��ݮ �)��F3fa����6e�l]�2~��~Xv�жٕ�$^��Ť����|�z!��_�`�/dZ�sP��wi�
�����P�P_�����"�GKe�k�^��\�G"E�&�ʙ���M+BU�kg*aS�ׯ��t)�(O���T�8v\;��1U�o��������D\���˩|{�f83�_�(�r��C���0(�ұ"&8yy&ɽd�MVm^�ٻ�#O��@�;/��廉�B�B\S���)x�0Wv���{_��Fe�yZ$9噙�`�;5;��Ẹ!kM��p>��dPlsߒ`�\�F8��^���'2v���[�%�#������j;t���,i����'�A
��U��+a�i^/bisp��~Ԋ)�\�'�S�L��t��oا��?�}Z�\?:��@�u�&Ȯ=����G���&�c(�b���Cy%t.�z�E��OiM/3rb�4�_��Џ,�DɯB����|���9�M���I27xp��h�q�y@h#��^c���'!)�X(ވ������2��S#��Yb�W5TcU�B���Rw�݅=���n�v���P_"�*H�����ҝ��ؠ�G<ƙ��Z+�"�r��tp��疌�?3���������"���B�0���K���a_Y�C�l�c�ou����ẽ��y��45�C��B�-ڨN���[������� ������(2)�'p��|��Rx1K+�O��K�H��'슏��Ie�ZM��B J}�1��ϔn��6r��|�WE澍��]�]����D��/��BL�V�"�d�w�$n_��3���õt�E$��`�r�Yh�<)��L�	�xѶ�7���-��H�P�Lz���	��jqd=��im2�{Ϧ�5&v���G\��՘��^TZ͒63
���>\_�����]{�Y�?��At;��ͫ����֖#:p�w�IL˓B'��β@Ѽ?�����U����r>ͨrX,�ԣ떜�̈���Nˡ��ԡ[�4u�Q3��2k��~��'&��~p�����o�̹{�G���V�m��P����L*�K���!��5�s%j]��Wx੕ZT���J�E��'��_B-�T�>E���W��\e��_���~�q��z=@:p�dx�A`TVFG7H��>���W��U���w*P��8��D���6�^�����y��?o�O�Ϳ��`s(�	�0���]�#\�b1�B�*7lż�,I��"#���Af��q���i�"����������+�o���"d�)�,Vզ�����F�Ц��� sˬ5:��u��)���������α����Gn����Eg�2l�G$�k�o~�A����x��#�� ���Q~��
�̅�^�?A�eg-� ��#�']��q�F�'�C���4\��RE�����W@���s�~1��:����3k%��W^����L���]��b;���T}-F	���\�6�W����l�0����%����/�\_��`�"w�VE�Ԍou�+z~�(�N�ۨ�N";8�%����ٶ�J�z�W�}F�]i4����#�UK8�ʠ����r�I�˝E2r�Qvb�	��d�x.��O��g�YA�NK���P�Z��<io����5qP�wf�!(�f*��@K�m�Xn���[��3CѼi�vSJ�ѻm��*7/����bm���v}��s���m+�x����͕b�\�N�߃LnOȱy�����9�R$��t�'�q����jsXc+�/G1��w��vP�!����Ĭ���y��'�Ľ#F��|ejk���aǷTݦ���gCE;�R,�#F�RPpA�X�v�����Jz�2��Fe&x�˭�[�}L�)&C�k䕵�pVJ��ar�[�3���J{������c0T� 3��$�G�l�|6^L
Als�=no�>�9v� ���Vqi���.�s����F9e\�q~��+{�f��9�����򫷾�w�>�������՛a��V�e���v%%� �������1�m.J=8D����H�������2�c�פ��˶���/��i/����P���_�^Ë��N���E����L���V��˛i��%J`+7'�i<l��J�!e{~6�5��y�0y䭋��/J���N�:$����N��I�`�|��eӣ.���yM�y.�>�`^�3=qX�D`��4Q�?1���(+>��k�����u�ly.R�Zܱ�ۡ(g�7]����$��v�J�`�;}��f@��'�T�#?[f��淑C$�FB��;؃��O�i�"A�Kk�Y����q���xy�ߍ�f{s�`�	l�A&5�27��礭>���-����H��5���1W!�����/{#n�j�
��S�}k{*W)n�U�Tmu���C�
_2^�W�7��$ɮHl�A	�+��KN���H�o��J?���ǆ��Co�~YE�B��Ȑf�����ő^u�mN?s�7��ʌ��P�����N�O(��O� ŕ2������S0W\�M��&=T�!A�|O�I��}/ęٻ�C��F���c/]n�ɼ��¢�w��>�.5 �����h��LY�R��X�y��"3�P��#H�z��?/�P�5+��P���H�p�M���h?B���ɽ��pV�t��Yڞ����HJ��K�Fh� <�ɛ��q��Q����k���;GW��.��F�G<��ڠԉ1[u�<�������Z���on�h�x~�!���^wE��|K�T]ns�<:-ʈvF�٨�PET�̯�!�:�9�M^���ٺˉ�
��R��q��~I�����P|���V�|��նM���$*(a5I&�:����l3���`^�
K��65����Ҝ �MN���	A
,��2D�����0�*��nH3���'�m����k}9��a�cs��2OF��L|6r-!Y���+��C�_��^�Њ�kK��l�&-S}�>���X_���J��*w�S�3ث�Y� r�j��faMmV���PTB2?:9`M��'6<:�@�}�V������=�&���(���y�hh�I!�1�S�R�R,����/輌�_S�
0�hAq��*�&�\d*����0b�W4�������~#b.�%�E��b;�7*�����������c�nR߼V.�V.�64�v�3���<��DO�aГ�n�y�fS�?(@K�C�~A��Ne:(8�G��BC�{M:V��@���������Ӭ��,�~+�ݣ�<.����bC�@�Y����4��h,
��u���=gY�����<�K�O�����=�?�C�3�#�%R(:�+�����
������ٲ��J����ef]d�v�g�9��'�u*o�NƑ.�����Ay�c�0g}�����E�b��q�إ����D:����B+����Vw&Tx{�i�Z���D���s=���"���{Ϲ�ӑq\w�& ��ŷ�e��#��@=JF���3�z�3ۨ#K5fGk�Ӗ*2��?I�a_�mi���m?�(H.�/��䜄r�$`���eK�5�:e���7�'@vfL�>d~i�߅�R}����k��12���Ƹ��2e�/��2�@��-���d��j�m֒]NZ��-����-Q�u��w��*"ԜN��DE"n/J�����7������Gt�2ef	OB��x�U�^L�2�)�
Q����c��5���F4���|�JF����L����N&�Ճ�*6[kXY-�ޙU���^��k���v������V�z<��ۅ��\w�
�A+�V�^ π�joqSw��G`�6Xz�X�����T%���+.CQ�4��T�Һ����A��ⵏ	)/
��<�uOr9�	x�Cz�^�0��,�ߝciB���+��(��W��-�9-�O��3B@Q��o+JL��0��z��_t�n���M�m�?��G������9�V16��ѬX�U�f�R!sC�0���2yV�[#
÷��L��]l�E���AS>�Ff�a�r^�v����
 '���=B�.q��4���-y�?�؉���j��Gۂ���,(��B��w���H[�y���D�|m�E��^�Q#��V=�aZ��*�)���V+�G�U�]82.aGM�5A�f�6"�_P���J�b��V�(��l<�6I�)u"$���[ё��Q�#�q�c��c��U�k}*���.ȉ�O�cq��BZ��C�nh��o����B>���7��IXvY�#_Z/��k�.~� ?��5���C��A)�*�!˾~
���&XL/Ā�_5̍�>�dࡠ[5A��t����z�s��$�.��|jD��\��
]^�����y-A�%��0nMma3��gs�yBx� ��8��CW��l�bɡ:2��L�Hޞ�ج`���UǬ�P?�Ŝ��~6��a����V�wV�#
uW�͹!�����8�!Gln��U����G�xgY�>M45u2�����<�ހ�W���~���p�?�MU�؅���_��	��[U�Wf����ITf/�Ԛ�<|�:��Ϝ�-_����_v� q�R�Z��ݨ���Af�J0g����Xr��6\�7�ے��t�Γ�be��B�7�0�@�B�i�]=ް��5_�3���l��u���RO��}S���Ӛ{���F�I�d*�q�wXΊX�����*U�k��x@- 5ry�ǀWM tee/�x�Zǒ2#S����ZoE�5��yX�PFx]N8�O�u���B����{G��W�ί�E���6�T�������+7U��Y������:;@��altM̶g�ZiCA���.�M)�5�Zj��ӊ�l��ּe -�I&�"�i���Ǽ��*�5~]eU^���}��6q%˒9	H�r�A�@7"���e�eY/�<xa�W3���j_M��_:��O��#���2_�R��iD��a�U���r�^����U��=�4������vz�g�F"mh*�)}V��-�T��.��f{"�	747N5�mh����CLBv��o9Sl�$�S(:n���`�'KT��\�	A��_����?��@6�C�%H�3F~�_��~Zn* ��z���O"�%-: ���LQk�	p�O�ݒY�`,�g'!�?5��G�ȼ��ǭ��� .����0��ӊk�i^�  ;���:"�R� n�!R�X^��`�JnA��/��������������"����i(%����3�<��L���@����E �1m��o.?����G��p:s�I;����Y{0��ͭ�}����q�3�/oI�-P���ޤ��l8l������c��dF�`҆/�u�����)G/:ۏ��kF���ˎب���)����4߰�O�5�pP6X���թ��|?��2_�O��b�`.�1��̊�Lx��l.5֑1 ���[u������𸾙�:4�ov���>d��/��pٔ�"�*&�����9+�N���Ƃ��+4v��k!F�;,��ڎ����7���n?�����]*�wM�eML�4w����5��ihK: |ڇ.v'J���݄1��#�~����7sܾ�ѭ�H�o�I|�"�,��"����\�l��kXb��?W������T۪d�Gh�L�UM�,��v1>9�:3���"�Ma���+R�h�74P7�'Y��ð�fk7<�c���i�4��Z��o�t}�a������������Cu!D����á#�:j
)Οr���G�$p���8��UQ[���^)��2�bx���`�0���
 �VԋY?F@�B6����u���U�%e0�=k���B�+=�:��Q{�}x|�|0�E�v��
iT1���FO�,��A���y������b�^2�_��z������/�˱%���lb~��� ooY��.�m�A�zv�c�R68��W� �����:�7�L�-Ǿ�$R�(�fJ����h���l���s�;�F@nƜ�dXX,3�?�0��k*lqU�S����[/�!�lʵ�sA���JX�|�K�ׇ�ۇ��h���PB�7`��Zo�Uc��5��b UG�9�વ���
�\څ]k��� �J��V�s��>b"$����tP��ta��7nS��yX�@�K��~4��%ܲGh���< e^O>iW��H=���k{p��SD�L����u/�1���P����Y�>�|��?���w����HXi��X�sA.*�@`+*�:[[�KҒ�X�3�pT�!�y���ъ��$����G��l��ĬP��R�&Cr��xH��ݐ�Z�PDUɎ;J����^͘��X�C��^�6_H��IM�QS��Ln����h����i����2��蘌om�C�{� �"^��*������7��{����Oع�uyu*ns���*p�a�n?z��d�k�4;�=^�(rf��w�paA����`��ɸ=J�����}�I�JJB��R������H�,�!�0*�hL�b���ׁ���"E����ulV�3���Z�V��\u
J��χ��ȳκD9�.Z�X�	[����N�s'�ДJ�Np���LK���F�\�8L�Q���$�RD3Hgrs�� �/{�R���/��L��F��{�rx��#�������Ut$n�h�Y�z��m)�oq{��	��)��jƏ�Z�cq1�/Ƨ���Ƀ1G�X��`�d������X��J�
��,��)�"ɩ�?c�����o�K��q�nux�2���s+|�z��/N|��b��� ��l�<�������
2���k��/\��ť	����.��ڎ�V�{(������m��=K~�Ĺ7�� K���_�2P�
	����ߺ+�R\���u����P�.�<�e�n�-i>UA�yk( r����RÐag�5�0�S��q:��i���Kv!�)��&���ͱ)��}BFV	c���O�վ�a7h1Gc�Z�~;��wAK~hւ�ȭ1��+#s�!~�u�0Tp�oz����.�mCd�����q�p�µ�D�UI�fO.�P�z%癸�ӄ�M��f� ��u�y���Chp!=l~����>�D��F%ě��W)*�,喂0}z �kRO�o�rp��wqsC\���2cj���	G��J��¥o�Cz�������~��ǲ��lQ��a5�#��
u�*�g���������A��h���"w2BM�c��5fJ��UC�3@�+&��pdBonM�"�����P�')��/qd����7���-�l����L�6D5;�f9�8�+2�b��C�?(����~cV�j#����9o�F69�]������/�d,p�9!�+�pU�F��=�S�B�c�q�P�zm��"��[3_�c�v�t�Y��_�N�>sR�n��c�Pue��׉4$�c��$u��7�#Q���k�*xP@v{��e��Q�U��q� �j'(���r�y�
�����⼌@��U_�^)l'�Z�c{t�Z�ùɏ���~a���oM�sfe4���e�N�����I*�+�U�Wd��R`b�L�՛5;��*����o�t���+��{4��s�l���p���u���Ҍԫa_+K68�@���b�MLcs���.dG��#�%r�hpD���
*2Lť�t���+f�ɚE�O+N��	��%Ɂ�[R�n�Ŕ
���'C8и�"	�V�bɧ,#V�w�!�1Yz�����f㫖��*{�0���0_�r�{wP%�tҐ���BRg�����dg�B�)aYy������ɉp�#Se�N	ց2��	7�RŮG�5*�L��w{�& k�j`�e��B�ބ5��^�)�F�9�$�ohQ�zC�3�L�6S�%�`�~��c*C2������̉�~7ޕ���&>�;ɛ*:+gh�E�NZ)��=�r��"�:-�"����^<^'s�`�\��k	.y����t�P�L��!���U��A��=�@��ڒ��tx���^M]"�	7̹��>��ӏ�i�n�t4I5��^���s	��O��>:���\Ux����2ߗ�Ҹ�/Z���O��	�p��w{�L��"v�	�9p��^���"��R �l%�CE�G�7�I�W=[�Y'G�dD;�@`����V���sa�R,XjQ=���������ǻ��cr�ʮ�� y�IO�f���]����`cp��]��Ц{L����%5��4�V��m���@&_���
�ρ� =��RF��ou���꧓�6��<:N�ލC&�L,�}�SϱCZ�c����>:vÝ)Y�{S�*0ID@9T�����=�����S0��b���f�aY�+S�����b�{�.ݐd)��u3��#�M��(T�_15�� �����3"�F8l��ګ��z�Q�Ȏ>�kdQ �M���E�	��Sq�>�X|Eyߵ���?o�!��)`�*!D�6�V��j�%����;D�7e��O��ɼ%04!�n��FSP��Np9�^�.v��w�P����P�.��FG�i[�z<�d7����+�݅f͚��= ��Vs�{��vr�5���Bߣ���/�E��z%�%�v���N%H��d�,w2��%��F����;�� ?�Z"1w`��ܤ����퇲��M `+ep��e'!O���vOΦ��>�'m_��ڝ��� \�0�e4��:d� k�dUʩ���w �����4.u��CjG9ܖ�Q���j|�/�5�3�dx�@뚩+$����u�-�n�=o-�ԳD�_�t���T z �W,$���:ҵ�S,��w�7�A�/)M��i���.�?��H����t�����Y�Q��3Lz�G	��E����Nh�blb5&P
÷�E@�_y������<�@��7�qb��������>Zp�3\������{���
����3�!��L����|�:�5�^��'�@��Q���$4G�2 �m��/8<��(���/�O�N��vt*2LE�'ߺ�?(���q��j�����܏^C-�Ũ�X��a�8~�������=�������hƘr�?{���S|",�(x9I���P
%�0%��ypv��T�MԀ�.��&�Aj�,���>��ka�� /-�,�7x|���
�R��w��ϭ�S��fˮ��9n�~Zݯ�,X��0�tV�u�5�����20�3jy0Hr��غ���|B?/_���^��░0�*�)�Cr�a��WD%${˂O��j,U�d㊯��W�5H]I\�����Qn��� �̒G����O<d��'�Rk[���/7�"s�n�zZ��J �����Z�9�h�4@��B.UL��m3��S�p�z�h��4��e�	��x���t�8���J���/� �/�l�h�<����r�]�eĎ�Nu�;�ͣ�Ԣ$K��9�9���D:�܇���2�ŕ4� #=l�YV�ڞ%TǊ���3*ڎѽ�����!Xh�`�M�d��h8� l���J�=��X�eV���[{���_��$I�_�����"/Jd��5�xțm�"�����i�����5�#�͆���>�������'�?�My^Y��.�Q�d��N���w�6S~A�t���	K]Ƭ�lO�2b�r�v�v	h
-��#�BF��U�Ji8M�A��3�ɟ�Xh
]�G�|���P��ρ-�����ߒ��23�]����^��k��M�q�\"`_���e��n!=v`1eC��$&��Y�h_foq��Lz������V�9L|�/3J<��nU$dU�V+][u�Q�/�8�V���}z�7��?��Sk�����[Ĥ����R<i.��ZN�Z��=?3{^$���J����ajQ��þx'�p��r ���7&�i�+j)�h[]^3`
�O:�q����4r�pˁ8��nB�D���u6h�GD�l��1���q���Is>V��� )p���a���l;��R��gkǸϬ�pI*�ȫ8�{<�bA�s�FG�y������,٫�s�B�[]�r&��ٷ����6W)<��N�s�3�uR7g��/��)�yl��"��۶��K�U�^7���R��M�|f���ư��]����sQ�x���M�ۧe����� ��5�f��~ʻ���	�<{�	�?[��O�QoVl��9��n�P|�3Z�QW���O�FcMMߥa��4
 �j,�2���D����#Ҩ�uqTV��<4��ju����y�Qs��Ԙy���蹺7짱ӻ�>4�d��)����bu�_s{A��(}u8u�Ҟ��'��X���h��f�^���K5|��c+p��f��u�?��^P�����U$9��aP� �d^.�#�6�{*�=���m��Ww[�7J��O�@��+'Y��j���	�h�?:�.�1M�]���p�%�����О}v�4�-��
��Pb��Ͱ�ҟd $ܝ���.�Uw�=!)l�#U6����1׎E�a ��W-����q��mï�wJ8/�z�N:Z�?`���J%��b����0P��F�cO ���,�)R���b��zL�Υ���	�s{]�w4T��k�Q
?āJ��q�M�-��}�zO�(/�qE��o�[�q��*Z&������u��{�C&N@�A赠PTGA�ѻ�Rw�\	�#��T����Y��;�~��zJ������
6�F�����L�o��1��#���Hx+Cp�xw�9|�'����ܳ��K��<�_ `2߽�?�.�K�lJ帝k��w���k�aV��F8�F�S�Z�t]	ˢ�`Ԧ5*��k����mP�o,���A�Ѧb���~.��E����(ez�D��K�GB��	h=]���o��(��A?š�����Xs:8��R��� ��s@彠�%J^Z�����۶�ђP�\T`��{�H�M���3	�4�� �TK�賯����q�Ӆ�l�U_��]�t�{L5i��m8��fN���l� �y�bF��6� �����<VR��@��M�uZ�_-���)����F��]l&����-�=W���% J�r4��L�X�W�{"���wJ�.-��܊�����Z�SѬ�$��64V�G�r���aPҪ�͛����q(�N���4�n����Ec��XK�
�)�k�J���_fȾN?���Eo1���/�-��)����tY�&=�`/��0%�Y|�ORa�Բ]�
���n��ފF���Z�(�A�JE��ei��)��L������
�C,�wi^�<ahdű\�j�A�_�{g�0��S�vtC'���
21�َ���H��/p[����[��[6ܮ,vtm���D���GJ�Cq����G�
H0\Aj��(����A]|�gL{SA���B2�R 