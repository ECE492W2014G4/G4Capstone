��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P��v�"<ߞ��&'��k%P碶�R�ӣ�sĞ������FY&-揍�2�IԼ�<	�󉲪�Gx�I:�7�Ó� �狈%hX5<�'�1�.BCs6]ޯ�ن7�<mʽ�������#+���?��G, �������\���n
%��x����<7��h�Qtt�E�T�g���B�/�n��&��ڞ��DSM����X�_:8���������y�T?�3�v������QY��a��S�H�^�r*�'�)��w|���낑��*��Q �Z��ZM�Pc���F{�ei
��L2��k��޽307=����3/�E����jaO{K@6!Pp>��EnK��ȯ�@��N��-���A�ɸ��h����H����@kL� ?M�h�h��_%>���o2�o��Rݢ��|٢�'m���g,�m���ְ���uYA㍙�v@r���V�<����K���������`�� �|��Ϡ��"'#�>��o~��_�����P�ߟ�����v�>��z�+��3�i����
C�4�TR�hG�ć��HQ�,��qKH�ʐ�C��$��|�6�*@�<��杊�]�x��愙��+.@�>?m���.�Ik&[�7���z?��
��O��9���A`T{��o�"yh�8/��LEa�a����3DdN@zLJu�ۚ���^ޱ6�w�D|]%�����44���&W�Ȧ ��b(�T?��~�!܅�?8�����%���׺a���$ŉ����;�Y���h��Fk��c�W!�	�7�!��ġb���ߊ�ŌRe�?k�W!����mw�a�zBf܉[��Л}oE�8��~��O��t4�W��{1�BT�=�ge'Gϻ�:�g{��������F����uR���u뙬1q�y��u2����Ydhd��x�T��J���>�/�}��z���FN�:?�Wm���G�Yu�@��|^�������[c?E.4t�?��6���7�Ծ�6��=�ȅnc���V�E��Lʮ�͟^�p�25�0m�)w�V���4#x:�����r"����Ӆد�yd��>��5$�%�k�� �!и,u^��#|��������MI�6�	�q�ө��7FU��<�Б��6��!͛��#de��L?�T��g@�D�J+��U~��
:�J]���/�ķ����2ч!����7��{m��k�i��G�C�܆��X�d`}FNt?	];�f"���^"�L;ƕ{���5(��Ss �q��f�@?$O������s'� v"-mGwɅ��eQ�5�4�}�m\����PrE[��S*�����0{t���5��ˋ���}-kv7���+)�-�ǥ��H5Rیd�o��'y<���Z�	xxz��
T�I3�� �v���/���*� �T����B�qy�F�_2@F.imF59[BD��}m���5�ֆ�lM�s5nv�T�������+����'L~�5��e���+oE�������@�t�M����21Zw��ta*�3l�`��b�Y�!��`1f%)B�����p�����N��X������g��P�I����_�4n�Ӎ���v>^�R���l��f�\ʔ1����?8���h�ɥ}R���l'&�鼥fgrGEHhӧ��"C�G�	֕`$�$�g�/a�m[�o'Q�6��6qBL��zXPj1�S=4Q��0�
���ZH��r���]e�b�
���v%(���-�;A��9t\�e2��!�<�ͳ��6]�nSh��l����������.(��:CQ!~��q<X��f�^�$[�,���(�{u�ܚ9eQ����3�GE���P0�D]�����3�C��M�9d��0��'��M͛�e�@���%�!i�{j���l���8-��h�z�^��iǼ���%�@����{3�믱�D�r,��mY���lA1���|e�_E.-��L��v���!#�9Ze �/�D�)��
�m�e�����<`6f�J���H1��0��笖�oy5��C!�b��U}6�W�4(�1H���u�ܪ�,	���]T,��ڣ�\�x-dG��'Ѣ�4���	X=�O�%�
�	t-x�)i�|4�h�4�4��y�6����6BtQ �?8�������Y�9�g�L���1�!���XgV�"��=Z�����h݌V �����z��]e�tE��$����}{G3>��bh�p�G`�b$��]�ƎE�����P^p�^���w� �3�7�+��}b	Cq�"���+��q*�4��9ٱ����~g���[���PZT��h�� }�c�ҒÍ��0������X�NN2m�R�� c��~YC{v�?���]� <2�0���"_�������M�Q׻:}(47��*Y`?���2�1�ŷ)v�}
|�t���.g^��k?�>�$?��1�	$����U���(�Fx�0�utU�*v z8�����e.�uS{�"�jI��v�@�Y�+e���ڝ���DW�|F	>��1`laȺ�:�m9"3=�D�е�U'�)Y3�;#z�bǤƶ��������Fp*vR��Q�-�}F���}�S�z�e	��Z��V\�SK[۸~5�y�MHH���!���!2��l���T�n�cF*���E�O�����\|b��>'�hkl�t #�89LA�ǜ��6��`�b��)�9��"K� ��0�U����1J�d!4Ħ�Q��yCy���6��[~L�Ղbvl�dɂ<.���K����Q`������mDW�I^_����z�����E֒Y1� ���Zӽ�u5PΝ:$�1x�e�����J����P��+�֍�[�D'�H�꜕Ә����;��	8��e�j����4�����]��Ȳ�rHU$f�P���O�"�V奟LH���Ӎ�jp3��8���{&+M1P0�-�}rU�N87Ԟ�nDtr����/�l5x�j@���-���L�m}�F;E����
}�rcWA�Y�q.i���Gt�И*��*X�qs�b�r��t`��p�ټ�\� x����.=��H�4�C����=�o2ڛ\UH���irJ�)������#�tH @�t'���.c�A����<&_�Z~j�h�k����:Oh8���Bs}�Z��u����;IV�6"�I��2�B*x�:�eѨ�k+��\�2���9zE�\��bJ�L�Y��}��3���T��*�w=ɸ�N��K��� 'th�[?](%��5�AL�u�8��Z��oR�Z�G�#���^�ư�RO�^�=5���ģ��J�C:�ͩbܥe8���K�����7��A��4�PP��҆g�	�LJؒ��rr4�͟��~�ΦȶM�{װ�V�"x��'���n�G�&�9Y���O�!x�������P7�W�cg�n�3TL�(��bT	�8�d���9ͯ�v{�d2��Ӻo7�ᐟ�=2��i�޴6<�k��_U������g�"�r�_���f�-~�{��At�ɀM��C�+`o?�ͷ�.u�̟$�����KN���
P��`?KV��B,��j��b:!?N�Nԩyz��p���-#=m��U[HN^dI��[��қ�����^�۴wq���a����W��9k�N�r"��!��/mI9~�(����#:m��[WF^�s-�� 14p�;�#�����.��:�8�����δ5����m���X�0�ǂv&z-S��v�]m���$�)��ɭ�Ě�"��a�ca]u�V�v��sl፳�T$vo3'H��=��LX}��(�&�p�{w�L�r�u� �:���z���TY[�.���ث���o:bZ�.�Dc��3�������Vh���m6�*)t���� ��h��GZ}��QU�1J�$o�^Wu]S�	9{��e��M݊��rh*[r���^��1;�M�T,����`I~�~��=�Y��쮲Qp��e�b�ڧ����@3���M>4����l҅�[B����ȅ�&�V�|�u�c����yy��`3.�pj�oѷ����[�F����W&7$Q��ͿC��Ҥ�<�l��Lb�W f2l��y�Q��X���AO'S~�߿x~��S�?�⛳�D�wjZ6�F�FyN�$�7Yv�Vgl�[�~�6��(Њ\�5`^���3���Ϲ'�醕����z���!� �2˕ӝ�H���qq�U,n)��.{��W� "�����ۥlC<���b�CS�����RO��E���os"�@�c\�dF�I���{���P�/l>�ڃ{��N[$�!B��]�>�ITj��[p��(�G�����u��!�G����$[�Qxc�V9���J��/B������9~?T4ŻZх;���-n��x����O�T����ɂ�N�)���@�����"�<k�?5ˋ����Ϸz�{x���?��_�LҀf���i|U���+v|��o�����K��A������.=&Z(&x̌#���?�X#?����<�$�<#��z;�$t�s����S����F��A�����PMYy�Bl⟪M&'{�t�8~mI���ؐ纷��6��Wzz��9�c:���T��[|q՗��x�!69d�>>���Pʤ-˵�rf��Ć�?�5�q ���(�� ^�bNM42T�6]G�i�Y�� %��AS��0�O�>�L��n{Xl�~�i�����&"��c�s�1��P���Q9>�!�!�E#����Qt��u�u�4�X
�Dn`�Mu�p�"��.ƛ>���a�<�8��l��'(���i� -���I1���٤��Ub�Ϯ�Q��#�_}�"4�Ƶvl<�h52v�jGc_߀+�̾aM5��M�E�l|A/���a�G-<���a��U���e.-�G���T� J��	�j$J�@$��T��pg5NҐ#�m�% ��6^$?�������'q�2+�@)؃��M2#��Blڍ���{
G$q$�%��� L�(D,e"C	bDlt��̇T����G����J� q&+I����6�.�=/� =^��'O����Z`�"�Vl&�6���En��I�g�zO٣WNiO@���V��;}x����|��_�p�`B+��&=��i�=ssT�1'�|��W�2Pu�!��Uv�%
e��~�Sn.��Z%�އ��>ď�KL��H��߬C8_y蜕gzn]��Q����� �y�X7��ɥ�+0
%NB�������&�1�%p©.`�{��rbd��N/D���<�a|�1	rD�+�t&��&���.���{~q�7��y5�E�ɒ���j띿����r�d�m:�ФKK��rYV�侌���x�D�W R	m>�IP�D�$A;i7�0�2�~#�-jۖ7;Dp�4{������@��<|���wj)f��␢W�IU�Rq��^���CÎo��-��=@I�"yO���'*�!�YZe��3�e�Ϧn�:/'9%��Jb��
ό:���� w�����g-]�"�1m�b������T'�j1"&WI����������5�Sc%�_W��c���m����/t�VɊ�	'��h�Ѿn��yG�z��H�r3�D�d�xYii�&jn���H��3p+T��5�$�%);�z�
:�f�$�@�v���:�A�ʆ _��W���w�&F,=8c<��:.޺m��!�:��.��O���$���M�NA�'��;�챾������c��u��(��_$������Y W�"�:Pۊ6H6%\��P�?ݜv�G���Kىx���W�?d���E�3����^>^��J8<^�����E=K`�O]�֔��N��[�R_����G����#���I$�~H$L����6�˛K�����"�?[�LY����x��uoK��
�7#�;ǿ,Ѵ�o$��@�tI�7�оX��;���t#�Se�u�k���jTⴝ5�t�]�w���R����4�#o�?\��&�29[m�}�,���u�x� =8�qeiPJ���S�L:�<gϔ�]�V�R7�'�A��d�ѯō���o0w��NP�k�'���e%\�i;P+�.�א�p����)@ �r1������� P��=RRY/���~S�ł��Iw����R��S��`;�����|-
��o�/�o���-��^n�B�7�@ W����Th7�c��w�nM���]��)��'�AM۫_�$:���et�u��� E����g&��D��r����p�2���@[�0��� E�g��ю"U^�֖l%�M�6Qu�C�`)m�&���?a�"����4{=���T��̙2e��H0+XS>��������r��u�:n9B�1��4%�f�T�d����\���WU��N�xuVF$�$�ʀ;ݜ	*g�F�~{t��TZ���;.R+oGN��V�r4RnR�!-����P*S6@��*����'TOXu�����'����_%��@���rW���n&�A���?�&0Q��C��'w>θ�ڍj�h�ͼ`y��LkU�����|�q���'�\�k�`  `���V R��癍ӱ+���_L/��E?�{. ��u��6ߨ�g��\�4�d��̺Y����.���m���т�i������9),O�]e[��ge�`��]<*�*�T��>Sǐ�p�uU�N�ӐK7_�>�}��'�1֛�.H7�Ym۫�=#.��~�Wf�v��~�Y���b��XK��Z¬��/J�B�*l條l�
��3�](+C