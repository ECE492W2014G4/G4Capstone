��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�"��F9s�`&���a�oq���F�g�O�]�<ݲ����eCL��D���{�5��8̝DFI��Zp\m|Q��
�}�6C���UnF:<�jΈ�2�����<����sf�k��,jڙ�����2��X��Ss�HL��	�������+g?���N�Ż�����|�v7�{M��VNB
��Rs�゙�Ld\��X�'��R :�J���^�����kMkx�Q���3!P}�e���Z�Y?.�U{�RP	�)��lI{tI(S
7ZF7��R:]��Ѥ�>aE�_fiL���t��,��Y}{+�ae��)q�Y�+�|9�i��ӔP��"!z�+ !j�V}aV ��.���e��O��G��[pQf
���x�Cx񍅜䈧�!!Ɨ�VL�wf���Ñ��n�ocژP�5�_:��3W����_g/�j�.��=#ݮ:�X/�b]fnY����l�㗈c��b�����!��Xk�/	��SHgnG�;}����Z�jH*�����@�i���2���dR�+�D:?^VD���~\܈�xy�C��y����dz�g�!+kh�I43�4�S�T���%R9˵Cv'J��鴽�G���=�Ǖ^��ҭ�ג?��f�' �8��_["�}9wV��5{g"oK�k��g5��k��+%�)X�^z�����T��5{�G1����Hp�Ws���b	�y��}'%��^��{�nv� �K;yR)
�Y����=vn����\τ�MЈ�cg �ȥ��΂[����UPq�!�S烑��]~o �R�c}�����Y$tn�6�S�'�;��66���ω�Ys���2u9�cW��r���N���)|GW�$<�b  q�R���mqCȢns������c���N+	��4�x�6]8�����}�Jp�l"�}3Rn�]����0����Ԅ~����2���i��9�dt���?=`O��M�+��t���c�'ޞw�bdjX���rRX6�A8�_�$������Ϙ#c�CC�C�ƷŹ*"�a��x��j_<��&Ԇ�x��_��00^��� Nkx�0IA(+G����v!�Y;Pʰe���JO���u!�4����3R}L�_9/d���ʇ��Ǽ*����������Q;�S��Z�lK!=�����8����������E_7��>�.������t���	#��vk���[���%:�;{�b��k!��ꌊ�w`u7�Z��*�S�skn!ɺ�㇊D�UF[*\��)q��t��Z
�.U�"���\r�=�7����w�"j�b68t��EQEtn�/�>�����b">�S��DÁ�=vi`
_1��ܞ0F^�p������U����NO$Z��lY��;�#�f��jh��ֺe@("���!f�tD��/�i����`���W�[�Qo��T�=>�܂�CW�s�\���
:�����w�������7�o�N�kb�S+�&|��-�	&8�&,��p`m�s1U��K���9�Veg�:1��s=���6����=��N�U߁'��v�N~@\�#H7p���Fa�?A=m���.��4~��s�U\��Js�9ѤJ�
���z:Z�q�F��TT Y�E����X�t���bez&��B���4xCH*��!������ľ�^C�SfGn�U�^H���uH����x�3�ҙg�UQe��1W����}r��.UA�N�o-�n:�ݟW���K�O�]��m.i/ij�`^���G�(TA��e��e���H�'n�z�`gV�Eie�I|ђݿ�7K�f>b�d��K�vv�b�c�!��*r�T!�^4�}�#�I��&��ʾ�)�r�?2T!��/���	�-�M�y�P=ˑfw��tY�� �,7���!Ѓ({jf�����!ݹ�i"'�g�]�������m�46�����y'X�WߘF�t��C)��G[�U��ǡ�4K���sd��oځ��X�,�dUe}���Y���o��0�8�1[ s���+=Ԥ����/��Q�u{�����\-�g����۬d�oƳ�kP1��m2�2�c�YºO`Nac��Ⱥ�� �3W��GL���%|H�P��ҋ������4�//�_����hC�r ��\�S�=Y>֤/Cg��24/uꔷQr�N�b͎�F�!f���H���-���&�#��B �e�� ZKXb.�q ԋv"0�8�E?�F����C e2\�P&�ֵ�93��A��P���A�$U�3`��GG@�'���@`13� ��E�Ի�?{r������J� �G�f��K!ƙ��u�)#���Cڮ7����GcW\aĵ9�Sň�{}Vb=کG1�(W*��#�k��Wu_��W���ȧv!z�A�ޣ�`�{g񪤐_^i镧�Z��+c�$���� �L�c�k�V�7�-$�r�;]�-��(�#j�K�i<i�������`�[�"��X/lY`|���?�vI'�m��h�/�a����d:X�k
���2"��^�S��~BWuwlq.�X�j8ͦAd��.Nl�ɜ�5�$� �:ɁA0�����5��$�.T+ʡQ��ۣNʴ�-�ꫧ���aR��{�{��� &a�4�S:�So�O�$��Y��=V�S����r�T9$�`��2E��D۰�,�[L����<�_�k�4�G�C{��\R� �D}~���G�����2ߎR��O�U���)��ۓ�"<�������Z�~|ч_o1X��nՐ$�q"X�o��͔Z�V��fBA��MG�v�4�r8�)c���E�q���o���\�_rK�g�W*d���`�/�_Q�Q�A��k�1jْ
�)�ci�n���EQ����W����y)Ub��JT}>�ð�70��<e�a�rͅ��LfȎ�t?J����2UB�ƺu��2�(Ґ��b��e�g-��j`�"V /��G��f ����ꍡ=?G�aRPU"��Y�c��:�0���r�~t��G������vBE@+r���B6H�P�i�
*ĺi3�eŔD�-o�&5Q��C��%PkmG��%���&��ҟ�����?zK��f�;��kY����1���\z��ۣ4�C����%&ARnT�7��+N�=���?� +��B3�P�"������;?=�����QG���P���n�˖O�+�S�yl^�4<�Kp��'p ���&с��֏"��1�v��o�ێUu�uN����v;��*	R�8��}Ou=@_��GG������U7VN��%������Qj2�'>����YmVϗ����R(�<� ا��2H���$�kq��>�ǆ~�0棚v�\�,O	wM4�5f�?�(;Q
"�I��:��r ]�z<_����Z@�ߖ�N"�ϖ	���x�.�Za�n�ޘ�N_�_D�����ؓ�O,0H����`��'abc@�4	I����3W#�rЖ�+b� q��E��"|�M|:V��M���~XRU�ϝ�F��}#��&�V�&��ve3:6Ti���4���0�VI�D[U@tO�G���`��+�=u�GK��Ν�����O'�.�(z0���ԛ��(��C(UO~��1�w���f��f�Ǥ3����U�����6����40����������!��V8����޷��_��ܪf]��03�愋�M)9V�xڅ5EfbYr#Vb�8��\��|������Y�� �9���-h��p!,p�q��Cv��vݟ~��%gEl���S3���~ΐFJ�7yoT��W���]�ˏy  �F;r���:����U��Z�񈈉R���LV���[���4TEu�����^B��2ම�\\�!
�t�%��q��f��g���V�{����i;�F�k�� �f��uD2 �!�CLd��LՄ���1�����q��w�#�}3I�){篨/�aq�j0r�qy��[�T�Z���i�4���P���lL�ּ�\���!�1Qޮ$}��^�H�5�Ϸ�\Z�,�%^��Z�O0bW�f(����7�\
�d@�z���ʇ�8�k��5�����	�N��P���ʪ��@{v_�:F�a�-�i�?���Kp�|��TBɃU�Y���-�_Q)dew"����Y�'ׂ��[~���J�er�y(2��(\�i(�F��5���ڷ}�X�ɍ��DGŚ7�� ���=	��4���@���L◵��go=>_^Z��iv=��ey�k��M��x�j]��P���˃�'�����&>�C��"L���v��.��`��3�A�f�i�$��%Y��eɶ�>e�c��b�r�j���!����������EVYZEW�$4��O>��e�m41����-j?�ŭ2�.K��-��"w]$�}�iI����T�+A-���h��wV�>*?���GO���	��s�����Sa���px7Snj��/����d�i����[�e�C�;T8����t�O6U:< �
�/A�/�$�k�|���B��y��T�W�+�����PLe�=s6�{4�;{������|�N��Cpv"1řHP�E��Io3�s����1���o}��6���nb���|�=iW�1�hٗ ���:FJ�G
�%WV�|���R?CY��:
��	����F�pH�^R�Q%w����$mO�փ�:x@�'�.ŉ���N�������rR� :����"T~����Pw���ʶF7�KJͻI�*[_���հϘi��߆8CI�5"N���c�F�{O�Q��"����uc-ʫm�4�mfc�*;�2|E��M��[��;Ѓ(�o��ں�r��� ��5���*]�������"Xfxe��w$r��/<���*�s/���.	�k���I�M;���~��G@o�'J:uԔ���\n9��D&��6ͻ~Xa����l��ŷ.��eM��9]���ˬtu�wb�Qh�|�3=��0�4�UX�O�k�?Wf Zd�ზ�-q!Ac>�0f�|$�����1����QV��7wc���գ��.7CZrH�Ȃ}�[]���$r�:T����K��}� ����CL07�Uf�o�A+���4�X${U*��y��d�yi+��b��yQj:�K�?r/�?�Y"���Զ�1�2��4n��6ױj��9{拣۫����ح8�}"V�Ec�YH{{Ͱ��pl�Zy��N9,wX⓷�!Q��h�ͬ�W*�ma���撼g�x%����s�ʺ	�������tݵ<�X�����Q^�U��Oܻ��й��a����|@C��bR��p~rdJ��V�{R	��(z\ZB�,*K����og���n��k
�r����a|��j8-���I�Y]�4Xi&��Cj�
/�w:�MGŪ_k��(S��(�t8�1j%�<��fa.����~bu���$k���#p&;���1t�kZS�]H$���#ӖX�G��h\�b�՚�e��H�m�^�?Z�au�sQ�38!__t�(3�ӿ�cN�s����yһ�&$�r��!�r���tF��M����m���ox���9�媛��ƴ���t�U7Ƨ龀�d`�Cy}՗��v�	�߈�Q���k��;��~���P�}_�wuQ��N�[�b��!�t��3:��ixq�A��K3�c�rN��@�����.5]d����U�G���d{}`�ʾd���"���?%��ǕL��^������t��J!af#�����GR����rJ��Z�l��[�KS�U��4��m�Y��[�c�|��E.�L-��H�����f"m����؝����d\�E��<#%�ƣ��In�8���I����Z��.>?���brӹ�}Qɱ����5��6������yXu@�ؐݥ����ϫ*A{_ȣ!�"�!؆ ��dg�e�ӌ��e�����R��\B�%�q����{�0��� �\/E���z�X�L����c}n���l��՜��kv����;w�[R�bW�}�Fك�+�!�@P�x�+�$ފs�MϾ�$�^O�85��K��?G�Dj10h&m������h�8bi6@�2�EԞ<�@�
��j���e;6���+h�榃���vy����Ȝ����-ʥ2�Y0'�Y�}�>ٙ4���u'�
�� }#��N��ϣ�d;�v(ѵ19>�X�No�-.���Ų�V8T[�Z��IуV�98����j��k`3��u�Ay�(��ٴ�����d-)=��w���*S���-���;-o� !J���l����.yVF��=�t:M3��ƌ�R�3~8�V����*��(U��%2c�l��>�~�$��a�Is^��s�Cm9	�?���Q�f��}�*d r<gZm3tDz�BF�SoS#�� ��L�03Id�M�w����TCy�u�K4#��`G8<J�)������B7A�%�-�8[���ٟ $g�r�5�v�1�$�^�S������o���ȇ�s���g�l'��.���2��K�;��s2���o�C��R��:Mٴ�nEr��`���5�c:I�^�:p�3����' �\�.�2T�ҀI�v
�'1�����U"Asx��a�{�����_Ny���6wdTeI�)Dݿ�:��Խ:z�q�&�Gͱ�RG�o��>�3�����c��h�P	D�����R���,�K����Q9c,�l���H���tfE،�'��1�n�������:�(%� ���`��qBUj�L�C|Qw"������]� ��څ;#�\"�Q�S�i�/:g��_�
�S�sȞ��F4��F�/c3�[_������ȡ�LU���!���T����`�ol>�p^���9�%�I�@V�Ot�⵷ʆǖ�ᔄ^��.u* �.�.��'���`S6��m���=��e�sa����q�c�Һ��e�x*�갭��i��Fu%��s�V>,�a',5F���A��N�+����m9���K`Ĩ!(�T�A�8��%]ú0�r��;�"���-�H-���M1*s��;�ˢ�$�/��Ý�VYco��M��v��d��<�O�f�Lh�{A	��,l%}Ԩɱ&��X�>��+�5`�xhx�X�/�ޠ�=��nª�};���Z���,�ME4a��\�-�W�f{F�Y�"r�}|�V���@����#�l)Ǜ�=�5˵%t;�V�f�=+wc&#���Q���feT+ �GÆ=�ҽ��q���	�ߋ^�u��N˕`t�*�=Kx���KW2��z�7�-��A�+r9��#&����Ip��8�^�gMlp�ά'�o�t�=��bH��p�P����	"> c���v~�u�?�t�6�h�ޯq^�w�U��o�4U���E���a�$��p�������x��q�[�w�.��
/�N}ܷ�޵s���-�ؙ�BՇ��f܀�ΐPG6oڻ�e�IID�K�E�܋^�MKb�����mL��.�Ы�}�x�t��GPa&m�5�Q�N�Tn+���/�v�팃YT����@7KZ�5��d�AJR@���ن�xۦ�}G���ا�e�E��7�N�ց��pxG�ճȨf��LC���A��``l9��@�/�|�A�2�=���s3}Wf��h���2l�:w�!�5Wě����1��4%K��� V�g8:>_&C�6W��P9YF^�� �Ǡʾ'TZ�w1�䎌엁n-[��:�	o�"��u��X㼦oe��3��֧"v���"m�o�b������P���FZ����p�|����zwv��ꥧo}��z�{�r�+SڑC��KPK�b\�7�Q�����K�k��̺���� s �-w�]�P<J�����?`�$���<h� �Hjv��q�)?������A�3��f�=�
���Ëe0_����3(+XP�zX�t���J�KQ�+tN�7�Sc��![(W>3�X.�^K��b��H�S�yx)��'��CΙ����n^� � >J�1���@�ט9�_�Yg��x�&[���Q0C�"�N� ��6k4$?��|�O�uyI�a*����總%��@���5Ş�ac{�x"�:�� Α�et�e� ����$�غ����MSͲ���I��r1�˳�!�s�^�is��m�G�c�;��uC�hzd>!`����]>Bd�w� @qy��Va�]�赆�K��N�ށ����3�����ˊ���2B�?HDS��/B��މΪ�����̴���<���H����H��"��hΐ��@�ڙ���Z�?��L��#�/��Z��uZ����3ΖOK#6�Q,R`!�B��_(�0�*8-Z��D�O�sU���!
�9�.\Anr�d?�h��f�9#X���,�ġ��7t-���a/���V�C�ԅ\Ɨ�����i�M��#�)�@<}��y�t#���B��G�v��@I�0��p#�������X^�P��dxB��'�[����C��EsRTao���;����������_�2��筽]|�Q�]c�V傥����Hh5��s0�2n�J�-��":�(���l��.���=���H$�8��2����
;�*W�e	AE��Ͼ
*:�����i&W{#���-���X莺^;WpO>1�"��r��	N�tZ3��5B����qw�K~|IB���:�Z/����L�n �du
'q�.�J]4�k�6[�>���#r9@�9�  pl2lگo.|�D��^���O?�Τ1!K��$�L��x1� 5�U��o2�LR���GYW#����'��]! v�w� ��WY��� ng�i]\�}8��������Qi����gy_/�~uz=��Fo�;-�@1Z�)?J�s-7Wɓ|pҾ��.��)6 s�p��=
s�~k��t\��Qp!`�I�I���
�F%�F�j��SWRB3����SC7����5�ǹ���c�g|p/k$�բ�*��0s�۝7���e:�	>΋\�2����H�e��|���x%X۴�mA���^�ٽRً%��l&@��k����)@�,EQ�
d���)����G�Wr}��M0�M�D�be���:=}d�$����L��"ВߦrYҎ�DCzz�q»PZ���z�5�a!� �ߴo��P,���  Apΰd����6Խ�!�%��'<�p!?�ҹ4�����)����� ��W�t;��yu�_/��ܳ]2�� X|ʼ�y=� 'P�d�V��dxN��b�9�`n8z�&8?!�<l�]��a,�yK����n(�<1=�n�a*�w���pn���F�x�
&hVc��/8o�����DH����_��@0��a2�_�7�[�Y�o'��+�4WL��t��w$�e�E�bY3�3#���L�'�@���ɍܧ�5�c<����������]0�� 	Yk8Wt9=n�Y�=�1�+��xA��VfVo�ϰ.�c���1"N=���Ō��;�"��� dc��%�.�د?�����9�BaL�W��RO�&
3�g�i�n����p���id�%wf\��MQ��9`s�|<?��h���h�;�u*���$E:G�E����Z�
@c�G���r�MO�[aU�a���ʨ��]��W'�e���/�N��	DTr6����o�f������@]r�ڝ��"���O{�Bu��	i�"K��-ρ�FuYh��w�_�j�gF|�n��`l�T��V��5B�ٔ�	b�o~ޗ%�a����C[���|�& &^�p���tۧ"��z���h�8�b�K��:�a�h����O&fYu�|���x�iM����O�qK|F��ȟW��'��A�C�Gܘ��A�pv�`"<�}�� �R�W�PH����tZpժ]����ޭ��1�Ŏi��Ԇ6�F��z\��H��"N�aM@�k;��=|���������pǇ���K=>�R0沎��*���^�s�1�Y1�,�ZizD&��=}~Ϳ�VҪ�mg�����MT8T�W��<��[�ԑ�_���: M�{�B�;��=�=u����DA��hK���+lo��C�4��j.1���+2��B����ވ�iT%�E�X� /��T�f�,<5�cb��,�L3J�}x����{�Ȫ@SOT��Й�y	�i~;|'ؘ�<)�R�չ�n�Ȗ-�@E]�M��U�'�A$�����g߶3��f�.�/��'�����(i�y#9C`ƚ�����v4�'T���y`�5v�!)W%�%��E??4rUNsXt��FG߃1�%e�I.���G�D�?o�=��б�;^-���xNبﷄ�N�K�´QdP�)&t�0@�^S"�WT����I��
 �̮݉6�4b$���!y0��8+tJ���Χ�����yq�P�꾊G�,��E�45v}￉đ+���a��^*��,�R6�|?���������|i��)��M]����C'+)T��8��M��vK;��b�1Ⱥ0,�}����%Tk�F�3쓃����c��5����k�0?+	P��@3g�K��0b�Ǚ��P�m9��/umk��C���\���Ό��
sv����:��̈́��5�7�X@�`���7��Mr�TC��}�|*bz�S�5����D� rѬ}��Ԑ;�R�Z����&�0�!�����Eh0�����Y�WyF�)�qt��w
���t��������;���!�k0��7��G�b�X�i�弛?4�Р�
uJ��d,��)K�mx�Ea��vz
v�c��k�B��y�ғ�VF����T|yӪv�`�T���h�츏ɥo��X��r��R��w�Ѣo��L͐ �
Q�u�����H�JM�O�p����I*r
��J���b�&�M��6���"J�ϥ�؅�~z�Շ�?�U�-�#Ot]h3�-�C�{��g��I/7�k��[��X�|���&* �Dx�����[�#�kؽ/�������z,�y��zd5r��R'K��M�mԮ��}{%�}��L��֍�J�������WF��y�g����v�>�X�U�$j�k��2��o�X��^_qմ^u�nk/��r��<�Y�v�M�;_��� �)�����eR�$ׅ,fq�'���"���A�PGE�K�,�5Rΐ����U�z��}�+;�����٦�*A`�c�)�^��E��U�,E�2]q�X�W����ݘ
9��r����dҎ?�k�a"�g܅>Pk0��M��l��ԧ*�����
td�xn�yt��i%@�L%4|������i��6Bg�O2P�#���SA ����b`F��1�\?���#|��g�\��<�9��9�Be��a|� *v6�߆t���h�3ٟ�e~�t��av�xz�-��ʞ2� �~�Z���E^f']Ft�z�Tρ4>����S?|�+&�NlNl,;����F:�x�8��R00�h�}�'�=�$����X�,�5�Z��F��dy�!I)�$L�sS[���<u������=�~�Kۤ<@D��&6�q<w�Yɞ�V �T!r]��������E�H�V�>eʹ���}Jgb;��Q��!�+�Z�Z�fۄ������*K
������+P�j�F���b�6�bL�D�ͻX�u�R�_.
C=������"�č����Nm4���^���_{C.Y]�~G�c�N;�R���=��l��HiQ����[��w�����Hi:ß'�dw쏚���%[/����^kX�j({�%�����>��
�}I��ӏ'�zȍ�z_�&�`'�
q��Ht[�R�0���c��B��Swl��N]G��	�~WX�_��Y.'�aóx-'x��\�:�МV}�KN���}LM��Ы�wV��*~JxL����"�wX_�ê�N����߸�a�	�WhHV�徶��b�R�Ҝ�Ծ"^��C 2}�pM�Y�H���Z�u7L�:�L���9�� ��w�;9�]U|�9��J$Q��s?��!���W�S�1f|������S3 ��[��ݑ���!�Pl���5y͔,�x6=z%ւ�yϤo��|8��WbDţ�˔׿i֟:�O��S^I �*X"9_3A���g�a.&$��d#��@mur,��շ0��j֯i��Y�����
�`��m��C���Sz��;)C+���#o�y�����t=P�SB��7���DfKH����
�[�f׭��Vn�X��^H��[�o#�f��z5F'j��n��]�"�[O���+|��V�yNb��q�U˫hKɑN� 7��BH�c�Aa�R9����$(�8��x���XEe%�J;5ci4�Eh��Т��|8V`j0�9�j��Sp�H� �CYA�M���xx(`uP��\@p+�k��r{yV��*c%S˖ܻTP��Y4�j8n/�ҧ0ơ�2Ÿ�(+�+���G��y5����eJG�]�vG� �(���vd�]�(�Jgց�2�����8L�����D�J����bJ�ύu�����^u�V�ԗ}���?��r�[�XC=�[Z8짹���z��=�J�L��R�����;<04��]i0i��ہ��D
����m����󹻾0xҒ4�����֚C���{۬��IPq����4�ӏ�1�m�f�+ԅ
~��f�Ha"�W �&P��n�G~�7G���$����gd���������Q���kkeU>�E��3�c�	�N��U��}@�p&��p�Kҁ0�f:����F�F�6Y��� ��+��q���9RN�댰�ppG6�N����J��/�u����h�@����������x8��_ޮ�����}2�HK^|�r3*L�i�6ٳ������]M:Γ���N#�t����ΗW�.��CG���|���Vv��`�|}^x:m"3U1�x ����OzM�Б$����Vl@�JD�ЀXM���Z�@²�`1�
�~"�1Q��N	q�C��U��r���k.���#bp�DK���&��$��B+3�l��l�9�-�|��\�~��B�d�.���K Ϳ�*�UT�|��&���<�)aw���� t8u'Z?zI0�� Ѻ��>���T��f�1����#�L���d��ke��y����I;�*����3�.q�=lVr�kZ'C_$Ԏ��7v`ؾ
�{�ҹ��D.c�8���n��$m��8����$Zd�9U9����1���z0HW\�|��<�^�F[$^ �3���C��Z�ʃڂ��@$�u2',!#�����pV�l]�8�%wMw���ٙѲd1�W���h ʑ"��W�^��	�I53A���%��I�'���[=�(vb�j�Ü�v�u��r��2`��jw�c#�C*V	���2�|���&��>�����q֎�Ǒ�b,p���x(��ID�f��/=��mس���<��I����N�v�>e��R	�%;&�6�3<�K��X�BzJ�9i��I�a��q!]7to�ȑ�&���z&��݀�B�+s$PVx�K�����I�+!d�iU�9�X[x���	���\S�����F}�6����m�i��z�7�B&�,N�Z�>��X��X�-L�`�򜢕�ku��I��DT<�ޝ�6�#T�$����M���X��%�R��q!6	rPT�y�/\k���D�X���J3��5�P�:+��dJO����c��rcD?���0���u3	���dC2=�둫]���-z"d��$�&K��X+I�]��6nP[���x1&�(Y����mg%�YS��`y��Y��E��>/���3>��쮎̌�b�_?K�/���Yh� |�i�^�4Ȅ�pq���֨P�~��$�=���M�i����ίZ�����(�e�x������g��P���^?���y�)uBĖ&��ꐤ�a�j��.���X�z�k&�'�A��A����\�z*[tb�3�s	[u�\cSpAG^�y�k��I�ƴ�f{~VU��rX:zD���I!Ypc�Fm�����et���T��U@䝇�Z��D��ͅ;��Yzͦ��t[Ժ����}Z�7��]rHG}	˥�HG(a5�9?�w���q\��{�~��mB؝��)pC��4��H�H�8\�u��TSq�4�0��IXe��DL�>ض�`�R��M���x�sy_j ��g��7����I�c	d	Y�[ة���-y�7SnO�</RI{ø1]��N�'�Ҡ����$#���$YD	WA�#���~|Ȣ���p7җ詭���8��~�P�u {!�3T�<�]���G�.'���|�t0�`R��}�:u>@���M%����0�c�z��f�N̠T��i�t���y^Rq���h����Ɛ�rx��¬�A���+���؍�`G�vfr��!gG��(13�,��^�Xy���ϧ�9+�_�h�A�VɘP����Ibu�ط�@�.J(WԬfeP4^v.�̎�#��ee�\5M/�b2��,��w�[]67^:.^E�����!Ԥ>F�8�r�z�b�Ѫ�	�f�GF--�wծ����$�W�t��͛�N�lH�A�v��\��<\��8�-Xr��+�(:'K#�w�Yg\)��4~������W&6W���V���U��)�����=­5�yX`/�L=Tl�t	rmuR�(��hgAH)���`1��& �[Dm�`��2�L4�ޛ��,�	�^8��2}��F���?�ɿ~����ͽu�k^。���#���*1T�D�M���� �1��qu��鰒/t�=�ԞŎ�k��]K���.��-Ͷ޷0T�s��^�,�tu*pR�CQj�w�n-�	|�
�����|X�=�p���e�A�H��œ_�ɑ��G(�!�Y�v�bK�_�����g�	�B���:�S5(���_XS� �����XV��>��4�XJ���� d.�d�6��Z�m��DA����z�"�K�Ǽ�B�*�R�����y�|_r�)�
�|?���p>e?���Q(W���&����[�gt�8I6�(�3�g�h��f�f�b�� 	��ݿ
�[�9�l�h�O���>0�j���"[NHJ��ݏ��#|M	����[Ëh�2���j�\�p����mB����b�T��"<�sK�9��A��p�=�ٱ5���C������K|���`��?w4V���nv@h1�?��`���^��~�!nf;K<�q�i�������L����Ή��C���k+K����9��l��$�g�K�:�n�b��/�Uc��໛��Z����R�v�2a��y3�w{#��d��rE?��r�;���W���(�~�1dy.�%�Y�M�g"��$��H\�@q�"��`0���6l$f���$�l�����\�#[b�{�G<��tk��sq ����U�
=.�W���L\WTR']�X���&���&⧝ DP�	�p��rq%Z�R�PY�{��!�P�S�M�	?���ê�P]��D�u��i���KX���[e�V�'�M��@KJV���?(�Ο"��qC��'Y`fJZ�^/p��3��\S�n}B?!�ӯ�1}N®��@5��/��s�����0ϙ�c ��:v��cI,�f4daCm�a�أ�:2�F0Ӹ�Մ7�3�!�`6o�0��6�"�Z��,i���j2�i#�G�K�����h`W�l�0Y���k�*�Q`/��SW�?��d�b��R��ˀ�nd9�嗥�\N��BnH���ǃ�6��Qs����DN�d�F�>{�k�l�԰�)�#q��˙�<YL"��&��N����#�K��&���Q�H;�ڲ����@U۵�ۆi����3Q��xc.}�h���1�OB������C�FJ��"�H����ܧS"oz|���
=�k�\T��b��tv@���{C�p�I3������Mu���^���L9�9?5���D�W������*��	0W�^���"%Q�%���$m`������v"Iri�W�{��v��[��<V�"-l��Wa/M�&W�0�[�%����zD���!�f�j&�m�B ��$k:W��{ͭZ���k�Ȩ+�"�w�n:�[��^�%�8��l�֎�0s!� �~@玨��n@
R�^"J����c)�8OǮz����Z�~Z�S�[ ��Ir��뇯>��X�y`��#��C��/N�x`�82i�f�S(`�ɀy�ԁ���B���L�w�	�}Y	�
��D~�!������ڟ�>$�41*y���я���v�t�Ob�]��z�����I 8oeb��%��ɠs�l ����}|K�е35Q����^]<�`�A��S�^�.�I��TS��ѐ�ϲ�h�T�e��kTO9�3��x\�zY	c�	����l�.�3��{M���^b���+����=vY����H��h]��L�<j�@v�ro}�F��b��e�~ݔO�&}�K*")��G��+�_ <@����ֻ݃9��9��u�M3�=$T�6�!�=�d���hfO�W�i{��~�}y��gVXPKr2�:2� �MHѷ�N�)D�oTkP,�D�\�S��"Ep�D�t����8a�\��ԸV���[���6P�~����7��u�A�4�	�Ye�$lC�����R����]&w�����G�y�&3��\�nh=~v��Q��=Ob�|dq�%��z:��;����?X�zޓ��:T��
E�9|�##e6GeI+;ЦÚ�ݼ�w&���2}Ȧ�;��y�Z��%��	��Ob��K�	M���ÛFh��v	~mCH�f���d��R@/�����j��Ũ��Gd��I�wSF�uh�i����Gљ �C���mro.�&㕣u�����Yg�}Xe4�Ҝ��z{Pߒ�f���|c��;��3�dR >�v3A3w��H�|ņ���LQoYR(c��	Q#��}�N1��I|	���?H�M�¼��E'E$[ٝļnX���-��䥌��g�,���ǰ>|�QV�d���k��I��� �po�����֟l�0�n�.��I��K ��1<`<CP���yU�u��ł_��¥X+��Fj3���\��6�@�s7\�p`'{v����31v7@f��fZx�=� �YMit�"H�8��<���%����[ױOW
t;���;-^�.3ޔ���O�1UI/�w׿&�JSrlu��ju��j���j��^1�Z�A�F�|��8��F�#�j%�I$Km{��c�F��q��}�%�ӑjM^~GăHm+��Xgͪ��_�	;�,��ica�	�1���
��b��܉�M��!�!C��W��N6���"�x�A"���"p��y�4���Љ�S�xMm��g<$��PfuP�M�.��⣨�[�a�˟�1=��"���)��jYҰ�e^�(\�T|;��;U�Y��-SR�<�ǀ�˴��N��LܷۭQО�GB4�=�c���v.��P>&�O�c)b�[.��­��v��+.[;���L��i?<���)I-��(�=���:�êb��x٪J�̜�u�����!��k�Yָ��c�´�4����H�BF�.�a|L0?�d�[�x��n��.l
r ���1YI� ��D���-��E�h��W*^[�%!��1��b�eARg�񟲑=a�y�b��I]���_���A-6�I~G��ڱ�o4����ˌD�&V�6��	/t@��-�և��`҄��e@	t�L��d���X�1enw��Q�	���X��� .��p�=���sZQ{ �1@�U�6��uIP��(���sg� ��Z����Ni���ry�:͍E���O'����_l��n0�0h������u廤���Ғ��J	pKyrg�`QA�ߑ
M�зN�2��&����_��AK@�k��/SZUL�.�طA�H��>�g;��d�i/�޺pda�>�x%xӺo���`:�\���e~$*W��G<7��pY�uo^�����Mb���@�����_����\y�d�;���v(�5W2��]��8���8������@���$�9�|J�ܻ�Y�a��#fp�f��&�Md16<�<����"|�D��Z���44�
���˕`�o�����wx�b�e�~:vrm�pFH6��~04���֨KEN���l;��5PGIhK����n����hr��[{���ܽ�L	+B_��Z�]��w�8čr2B�2�[҅s��0v��H%f��GX���n�P��K��z�R�[.�����K�7�#������eB8����-m��V����'�Of"���唴���^� 4Z��tH���0Ru�nѳ�r`�l���2�a��U<(d�5�,|Y���e/V�!ON1E3_5��=��l]������6��eSy>�n�}��3���wT7>�#�oE?JS��٠��G�%9gpM)ii���X��g$�#�:�/�� V����Ա���|�R΁[b�0q�ʫܡ@��Y�H����r3��s�Lw=#�VG$Χ,;,^��^�7����i�.p�.o��M����ػ	eT�&�Tc!w5�oxi�.�rzY��fL.�����M��tT���RG4�/�x�7�-��pŹa�Ȯ��̗�)�� ��_�;�AͲ������qn��W��2H�"	|槯�b��9���F��e���8z9���'�1�U.��4#��d	�&�C[)?��[9G�f�3:�8.�Z�����FK4�~�VE��g8�c)݄��	�Q�c���������>m�A���Y&��%�6V�#כ��x�dS�T��)�Ѥ�i�e�y��D�h����0#%%b6��o�.f;Gq���*�vǕ�����l\�=%W����q��3vٿԅ~S�*�m�t|�V�MR̫k<��2��y��t⼰J]����7��e�����.���H�,��_8X��M�S��Y��ί_1n���֩bA�ų��žʐ�4]j\$r��XwA(B<��������o�X�f��ZE+���^�fگ=r�g�b�PӲsБXs4)���*f�O���MRL�.3R?n�6��f�/ā��-J���u t.����2F���{<k���O��ROv��9�xx��,��D;��Ag��������0u�J�sm,��Nt����=���!�l(�VBp���Pi�?TN�)�VÚ�ǈ����%n�(F�ʳ���q�$b��s��T.�np�"�5����'��$,޾����M0�}�B��b}�m���U�����&Fgp�l��}�V���N�@N��*����)�uD���� pe�g��\f04LݖI���4(��TkQjt|��@����r�	D9���'5}�d�ʶ��O��It��#G�N���0=ֽF�����O!�aã�ր��,j|�+A�4� �L�>upV�-��鶓��(�2���C�3)߷@-��qEђχ��Ra	