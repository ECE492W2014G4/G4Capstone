��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�"��F9s�`&���a�oq���F�g�O�]�<ݲ����eCL��D���{�5��8̝DFI��Zp\m|Q��
�}�6C���UnF:<�jΈ�2�����<����sf�k��,jڙ�����2��X��Ss�HL��	�������+g?���N�Ż�����|�v7�{M��VNB
��Rs�゙�Ld\��X�'��R :�J���^�����kMkx�Q���3!P}�e���Z�Y?.�U{�RP	�)��lI{tI(S
7ZF8
���G��Gc�׸ ��C,�o�_JZ���"�u�[D����)��/��?��
ԓ�ٯ�*�1?���sX��n�w��tk���$D���q�˙B�^OS�7�����p�;,hav��^0�e+��6�P���^3�_�ĩ�ƒǽ*+�)f(��\��^���K�-JXߊ(foU�g�:����Y����saY�U5��<W�辕3%�A\�����YeC.�gO�j���b��C�@ NT(�r����L�̵��w1� G �e�ib���;xi���}��(���n��Β��~pFc�Ĥ��[ȩ\�"&A��W�~��60�Q^���l`y�æM��]�_�nF{+*�U��N�Z�S�w�DƌD�&���
�n3o�9��!�t?�_f�a�횿�=5Q#&��]�����	�̇�����9l�v��B/�,��K��	n�F�5Ze�U�|-�6�-,��mA�0F��/�ya-�ۃ���9��ǌ���Պ�,ji�x����M+�8��l�!�X���?�;�8�v�����Y��;���I�|�\$�(TVT9���C8�lw>��۞^V��y�wKI�/7��=��d�a��ʙo�伛5�}%b�I�g�X�)���8I���ǭ��v�]�U7,:��?��Vꐇ���[}3zA��@��d�E�Ex0̅��nI>G�7�pFl��?���}�	�������x^<DG��r�&Z����rq>��}�~��Y[�MKa�G��V��h�/S�۠�g�>���<'M=%����Y��Ln�ͤJ-��LkOCF�r3�c��L&)�qyw��wD�������z�>��)�F�Re��%u�ט���?�YB��8)��4%�����dr>�9{�z6&ZL�RfM"�G�X�}�׶�z�Jn��z���}*ͻ*?c���"x��X0�S��=O��&�h���2:���(�o�M�Y�ESY�2����<Q*?�n��&��
.����taF���b&��,�
��/eE\Q�Am$�v��p+��s�<3�ћ�^|��Z�!����n���P
�?<w)fA�j%�$^�Qj`��oi57�C4i�c`D}����\���`�K�K���j�"����7�� �	]:PԢ`$�:�04U~.��`7�t�n:��h��-�;��w�ظԥ��{ӯ!��Ƈ�d���x5W��a?0U*�g���؎�c�P��<��R\�U>[�U֕�yQs4�:yi�����zeZ��	��7�$̹0͂3�1�~.m�4N�m��ް
Bѻ�%��iP&_5�y;�)(+��l`��M�a���� '�D��ے�@1�V���*s�)�n���16O~[w�O����	[�� �	��]njj��7Ġt�z1}�A��8�>�j�@��j���R���������i�����ek����ik�懬u���'S�&
+��D��u���������Ҳ�E�F�i��ϲ	Q�C����Bc+0Ϫ$�X㚕���&���;C�>������s�i�^`��q��o����khͣ����\HvUXJJ�݆=�U�U��#���	��J���!nG���O��OJ�$� Qd�Jq�kx��ńu5i����y1�<
��`�Z�f����Z���5���"w_-Ѓ�V$1>�>��'|w���K\��h���J�Y9!x��#�R�M�i��N_�X��-kထ;Qd�;R.�N��Me<���A_P2�$�$B��R	���0�?)�p�ZX��cK#@���� u�|�]0g	F
_y ��Y�W�뫵q�C���;�K�v�������߽�*�8c�&$@��/}�5�'(�u�~�)�ޤ9�}������\�omP@Mj%�NYO̿Щ�_�<�ovf[��t
ph:޳}�瞄t!�������y�n��h���w�Uy.mǑ���g�M�-�Ǫ]�����{#u����L�fq���*���ݒ��.W�o�%n� ?-v�ILo���Հ��M��ݑ���g�K���J}��\��w���X�0]��I�B/´v�y��=���:��}SCٚ�{,���S&!E�|5k$y�ݫ�����!����r��4e�x05V�	#�g�'�x��+��j=���?��¾�c���?JBfb�f�����ρ�p)ǎ�U_t��o�?ʈ���&Hr��3Y^<+s��+�av�)��T�)7u�D�'p����P�v�qC`
��$[�U���(�U�O9�5Ǥd�!:7z9�@Rg�^Oe���4�Yv�3�-e��7@$^j���1�x�t*�  @�p�Y#٦i�<�_�%W|(d��l�i�UωOaP��O�{�j�X=�/���xO:�l��Q�l��c�w��q��9�e%�� st��n�Zj^��T����mܽ�\m�$���Y���~U�e\�%�m"�	�$*ރ�'�Oz��sS��!P���*]o��#��<iME4�OS��vR.��F�c^��R�zw#q��Z�z<S�0#�I��b�E>�_�����_q�Ї"�}X�5z�V���9~gT>�	��DN2W���_�Z��^CU��&����o��Am��X;4x<��P0�3���~���b�"AD��I�{�ڛ�O�
���t�^�?gU�n{��{���m8ɳ)���9���9[^j
]9`w�{��X�z���Yi�M��Z�&=<b��:)
�9[1q��Ͷ��M1b�Ͱ"
7Q�t[+��~���-Ǌ��UVF�Lѐ�K�-?��<C��������B����!�!AHf`�̳�����lHF7�wOQq۩�O���R鴼a��\'��ߧ4>��F��ڀ�Ә���N_�e�0�B3EP��k��Ov?$��Q�F+�I�`�W�ѕ/�!�&�Aꖖ��8�)�:�ň�pU˷��_����J^�[.`o��8� ��2LI�+�؏,
N�<4�҂ׁN2�I����"�v�����$�b��-������b�ʹg�UJ�'.:^�6�խ�w�ṳ�x�5!! s5/4o�8!�9�-T$;�/ l�ifW�	�^�#�ʶ.��V��j�d�i��T�F�\f�߭~���2�3y^�姨j���:��|�̥��?׍��ņL���>G��L+dX�L.:�����J��W1�}�A
��"�P��[ږv�1�;�%���'�B�5��r�zW�7LEq�3��p ȡ���o����Q�1h�)�_ò�I��+u�� �Y��{1:�jԓ���0*�:Ő�Pg�N��(�,���Q��|z%e�K����D}��һ����| ��.*��=lf�F��҄wn�0s��l�A�܆����K�YLG^`�}^[��E�H��B��yq	o�vp����;.����Qh��jut��s	)�=,�����m�le�Q�6G�{��>�s�{C�����#cWxhJ�? �����ai����8Y5��/��U�f��OQ�F-U�. �Ti4Q�~6g�:;���1�y�^F_m��m�0��U5+A�X�OF�|���)��[�x4!� ���YTG�	/��뾫�}�3^�Dx���x8�*7E�u�\z�QH�ⓞ��L�C�S���z�z��W�����$O'z�T�^ٝ��;���`�|�;�?�����%���9�s?�/'@T�P9a���9�hG3���͇>�@�D�lSMV�����:�n�XTT �8��k���
g�'}rK�H�W�ؒ���>J�X�s8��Er����n:Ě�nc������-�r��Vs���`�4H���L���|r-��	��6�s��#2GO
�����\�&ֿ;�9�*;8Dh�w�T4 h��@��:w�t�g�>��87󅨀?P�w9�"Km<�!�����<���!\lC4�99)$|Al�փ�����Kjn���BM��掂�?���.���^M�G�1����chò�$S%�T�7F�+�2ui{>do�H���"2F��/��5a����u%��|(�֟��ln�E�w�Q��F�C�[���0Bv���)�l��	'E���0f�"�Z��quG窝��f���v�.8a�V�G`R�+P�f�>�śF����=S�����snb������t^|�RR�'��އN'K��Y�y��!�ad�LY,��|2Ae��i��ę�X�W�Dc��v9��H5w�sXx��c^���C��]��&?�t�V5���M�hn������.������!�#M^e�v�⥂�tL��&�$̚G���
=- �W��c��-'�}�®�$���o�s��˺Z��|k���×[(xW�u�d��fw홳b�;���OS��?	lnP�K����k4p|�w{z?Kep��ՒV����D�ƜI�V�!��5����P�t{缐a����qOJaV����6��H�iU� `�I��d=W^P�M��H~��.5r��v7��Eς<r!�kL�q���z�cB��^&r��1�D 0,�55��T���U��/=�����A|5r]A���f|Q���9!���Ҹ�D�O2��>\0��J��V�A�� ��������l'�!�YB�o"�� \�U�}֑��ѳ�x��Y?��*a�qƖ~~~[��)�xo{���K2Z�p#�u<JzᲝ���g��"-�Pq�]A_�r��G�0�r�I�F��W�WsX	(��ɂm�N)\LE+X�7bG��;��֙[�nI;��e����|�q8����x�,��rvk��S��=�HnmM&}�F��Xk���S�#��J�·=.Dp��6�
�PV��au���L�!��Dx��"$���唲���6P�f�U��+F�#��ȷ�)���"��yq�pkm��7��]�S�s���-�=pv�����F���S�YG��T�Oy����NGe%�Ѡ�nA� ���k$X��Bb�1F��( G���H1�Q
��g��x~��~�FOW���u<��{ca N|�ȵ�2�Yū�-nM-���/����nǥ�Y��CB����Ug/7Qu�w�5'[h���;ꎸ/�H�֩5�ٟݯ	���`�SR}A..��ӲF�Ե#o{�1���`
fkJ/�+*kZX��V�Дρ=!�a�q
1Ѳ�$/:�Fk�-Mߝ4�D'�����;��	�əx��w�B�o$�po�9qύo��R-)@�g5ms=���� ���drL��{5��|y��0�W��T�n8֤T����H����yZ�8��篳-��8e�ڵ%4v7s�T���SfN޴�&	�saO���^�j0:���i��濄�q���)���H�om���֮�'l��)dW�M������,�t�.P����ۻVk+�'��R��Ķ�k�+UuQbM�1I)�P��P�{�Vƈ�b~�����y���!�h.�؈(d�nK��y��4�%�ϓ���Bj��C\ء0�d_D�榐貼
����2>L�Y��	�|����=�r��!r�"�ڴ�w��$S�_~K�F�e��C��9z�)L����r��{}��7�]_�۠ �B��!%Ul��b�ċC��z�����TA��Cl(��Z�&t���_o:g�d�4r�V����O�7<+�H���	�O�P��7�E�X�ln���ΕZ���Q[�gT���]p���\���w/�X����)\5�%�􍜈�W��ʆ�GI�.b�~��we؍����8�B�ɡe�����Th\�?K2��󽫜k;��:P��3�������̚�ƶ��(@�j��p���)�����mA9���(����N3�R��IE!��'�Zz(]�\�]h�@��?sro��/����Y+T��j��&Dc!Aa�f*����L�E�w祢/��1o��{�h,���˳�[���4��$Ԣ�^<��&]�~fMY"��x�NW��*?������tV�;���yN7���	�V��x�"t7�%�o�-�Ұ1QN�)��ڸ�4�;���&U&����k7�:�R�\��@0���Xga�k�!���E8�p^!���� ���@�&m���4=^颏�;m**�<I�O�w�F���T���/
D�]�if�7�}��� [�I<I�����rM7��x�r�J��$�4M��WYg���$J��#��ˆ�lV�z�2}e��ٓW�E��@��؃��.�p�B��K�N}�[7����JX��Y/��c��fM�Y�kl�!���	��z!�Ъ��1_v�B\`@���|�gw�H&�A��}YXq�s�}�E,��� Ө@+D� @ʦ��~UKΛgD\���;l�#�?�jL�'|��@���� >���ϖ���}+k�g_$60މ��y�5q�7˒PO�;/af9�f��]\�_��dI2����b��jP���}[� �w*��XTy
B���9��O8}Wļ����1���nK��6�.��T͟�������%��m�b��'�ϙ�Ѣ.lG�����j�S_���s�-P�?tx�
�êĮ�<�3·)�Y��[��)+�/nL�9�����0�ǅ�d�<voɣ�s>�ߍl�/;�����+V"�8ZָX�eKK _�v0�fsq�&�E���LJ�]�84��+�b0�EW��v�~.�ڭ'�Hh-��V"��R�1a��a�p����-��jfD��`=�|�w���lq0�FG/�d�f�7C�	Qͬ��с�s~J�2�K��y�J&�W��i~�1��]`����9����*�"��"���O���u;v)��+ˠ.�b�� ހ~nT�����a��d��9���z���EY��f����pYEC�����M�ك3�t�sŷD�]|nX��,GF��%�3>G�I=��o���1�C_��D*������o�����=�����mO;���z0>���Ŭ8�6_��y���V�~QK}���T���[�����
v��`�t�V:�I���X�z���%[2��i�IB"�8y� ���Ug���V�s[�6�V.B�ۋ[a�?���{�/{n/r��6�?tՖϘs�1����yx��y�l����u=E�n"�I��)�� ���I
��K5��R���@1��?錕+�wp������_x~�Ӻ�|�Y��c������r4,3�-IC,?�MST��p�U)K�O�*)��˨�<x����&�̨p�1�38M��9�6<�A ]��BX��8:���ATT���v��kI�v��J���݀㙶0�2Z���I��3.��9�G��k�(�c��1KJ�����Z~�v���)��YG9���!uh�/�N5��k��N�=��MZ�MU�@�:����]�c4�PDn��՟}��hc�Ȧ?ۼ�'>]��h�ep�d�n2
���vm�D����~���ٚ:�]����LZf����VE��Ox�5rG$0Ew팇��UD��EY���ⲟ� l�&�ȉ��J�"�#e]���$^�>�$�����j�Ǳ�y�� ����lD�%ڸK��*�|�ie35	��ӧ��#=�1{��|��*}3�(^Wk�l ��V��e	��QV.F����&@�z
��)�Av��E��7&+��V���Q�w��rk��=�^1�y��َ̣S9F��j�V��2�i��d��큩�48�^~M[��9:p�y�g{����OE٢�aZT����eaK�V� ��VKdmֽ^��9@P������*E�w"MiM�j��x��U����H�����A}C�V��>
�&ߦ�IJ��eXΙOdV�+��D(.w�o����[�M]��j5�dx���MT��z�/���?`ƆKCw�D�nQ�W������,6y��agE�鹢���fF?w�)7�`�BT廾�j;�`[[	����r�1�/4�n����O|��/�ܺ�\�(T׻.����%����S�P���3�Z=����y��I�v��G+�����D�y���'su:��(ToCQ*�u��v���_))!fa��(g�{	dx�jo���3�ѷ,���]@Pѣ��$y$��<��M�� �� hR@��e_"	^��<�sX`ʙ��e^���	�|�n7�/n|5g���gK�S�99w��Ixӱ	�+vxg��_���sA�x,`o[�+�u��i&�"�=�;r��L��Rڮ#
���iM����]����ғ�%�g������QD&j
fȚa��:5��z��22IH����8NA �S��+�V�ٽU)=�,�#���&�U(��e�3�S}�;� �lP7zTǻW��$ΊP;iPr��ֳ=�^�5��j?��Se���o�Ph���o	ӳ=�hj���B+����"E�OO���`6wa�3ِ�?����*G[e��`3i�B��~�G�Y���:�;);�D�8#��c���s>���6G�X�44QO�S��Z��IFC��C�(粘��d�9��kIn12X�q����f�����<G_���i����k����n��=q
� ���Y�%{|C�ǋ��b��N{����|?߆f�S���|��k���#,�H�J�^7���1P}��H�td���5$�ɽ����Z`q��8�8��y��'�I�mC6�Z�rs^����J��i�z���.�`d�H��N����h���O�㫞�'���-:-`�Ҷ! Jp2����Y-������6׶d�Cb�B�T�y�6��z�+gFj=������q�K	�=~�Wa�2��o��8$�Pћ�ѷ<)����R4 ����e������*���?�S_��슨n��?76a���{�tDU,Sʠz�=��n)�$�e�kpe�,vZ����[�?	��ےe�����	���J#���d�f�A��!�'�8�qnd��}717+�d�����`���z��X���4] ��a��,�e�X�/a���nzR����:�/O�|��I�j����P�r�X��G`U��i�1f}M/�Y�a�p�����'��^8f, J����&Ѩ�#���S�uU:$�O	�E�s x �ix�,#�˴C��
��
�,�?�6�I@��6��v�D�0��w�Œe�72���ϼi͜kx���)�h��厥��s Q���:��{<��w!���s�a�g�Ĳ!������g'=��{{~Ï���iB����M�u;�<�DdR���4g['��x&�}�����hK���;QG�V:��T�Md.���f�]���#��1����L��%���,{�X��t�q��5�5����`b������YU���/���Q���@�.:N��	��SX5��Bu��]%�W-���
����MY��N/�b̃�MUW�f�;��&g_�8H�cL�:�HDꟚO���8q�5#�}� Y?�� Eh
e��r�0B�|IF�
L��ؗ����i\���l+_�Gѩ�P�N��ظ�bb<4B�DŜQ�qEb��0�Y�;t2F�䋔\FV㛕�W$��n�Od��Ua��(F;�K0��Pu�|�6MZIP�]q��\D�ɉ�5�hl��D��{���S<L19d\�V1sU��,zɠ�j�VYG��ex�)�=���ͮ��!����L��.�U�/j[�����1�pB���D�gC��=��l�(��GC$����5���:B����&|}S��f������)=���)�N�G)��V'��m�E�ðI�̎+J����q0��H�5&qC<uF�Fn�S�p��7���9�O#�����α�W���9���=�q$�1=�b��zܰ���Hh�Y�L<�V��fMT�=C��)}
���5q�O�5��b-��g�-<C,N���6�`� �A��|mĮ�"���y��RΊ���#�2�y��myp<��/������|W-��8?t�II��93P8^g��>4�]pe�h7�f�!dzIw�F�bT��8��'�#����T����UҦ� 4���J{1�t�+��w�n�\UX�,c�6�v�F����v�1}���x Ꝍ(~
J����kp��o��I,8�5�/�w4�����'3pm���U���gD�mG�䖙��K	a������w��*X�����K'rv�j�S�,�*���vSN�J��I�ߣHΊ�Ɣ�u�"i_鐚>�dn��jQz��p6b�����ZKhN����²]q9" st,�`�_���9��*@�zW�%3A��>�Tv�ԕ�.zz3!�� d+�Fn����}"ʦ�­ V�K�嵬E���<SO��ww����l���?��Ќ$�$��SQ1�NK�T�R�':dT"���	ץ6�onS�ۘ��>�6�ސV}f�EX���ki��t�U�Z6�=�4pMJ�>,����a>�'�8t ahv:��sV�[q��NiJ~?�.�6��eB�,k/�E��bVe�CK)���\x��hQ�r[`�4"���@���F�36��<6������WnR���~C����t��	�RYps8�e�Q��{��Q��j<~gh��s&Z\޻�s
�ڔO��X�Aw�
�{�G6�H���W-O�BE��{�E\�"k*5nп�!s�f���Hf�װ���
-��и�����8����7k!�謸�	�k �z����h�Q�D� � ���*)�wVn?L��>y�ǯJ��[]��Ԣ�;9���t�b:�8�u#�EH�k���_Z��J����`"��R������l���Hɻw]�e��7| aʘ*虮�B/�P\j�ˁ�fP���X *}�o0��'�vs����O��(�U� �(E<6x�n��HO:"`V7:nWd�)f�NM-&�KҸ�ƀ���8#��k��ԍ� �B�9����U&1#;@'�d@1�Jq�,cW %pfl�<�x���W��Ԏ*e��D�(�Ǌ��7�e��ΡWe4��y�!�ZP0��ڤm���&�FҾ��i�m\�A}��+��Њ��?C�de�#���P���(Xn�ו����c ������S���I!�@�� ���&����@�D��CD�(��;���4(��BΑ,]����S=�i"�"ƊM5�R���ޞ��N���63Uyjә��	�ajB����g:�NR�*��p ���ZC��c��͞*ɮQ)I����07��[�z�]��}���}���ղ�RO�[I��'�瓸�>N�1QF�	,�{~��[$)kgi�о�w�v�.�c-�l ����N��`�+�m��&��3g���5�r-
x�w�/ �d��m���,�,@0�2�,k	��	<7j�����Xk��wrH{�ѐ�]tK�f��2-��p?�(����WɨAJ���?1�м�"vf�hA�^;��=����4(��%�gA��$�C��>o^2�nd��5������^�^�|���%�"��7��g��ז��݀�t�;��4�4�����<���X	�=�&��g��%��WQE���ݵ�r���EA3B�,?°�kh��=�N�JlF��.L�	�In�"ⳝ9��PJL*`����V�9��F7�����4��W������
=�y��j���,�s/�bk�s��1����C����̟�Q�\�)��3=�I@�69��J�f�7��᧮C=�Z�<���r��j����xTb_f�;��I�c�*t�'��R�1�b��F��q٬�Y/i��DL^���7��]\����ZJG>0`oF�&�$��m|���H�0������T�%q��e� �h*�W��X��a.��"�$Lo*9{7�I�+��q�q�ؤ��g e��g�M�p��I�,M�^���D#ܛ��<�yn(���a�r�-����h�3γ�� �1t�fg�&���=t����n�a��stۧ�t��Mߎu^�0 Ne��K�V��cu�&�F*Yxm
��o����z��H��f�Tb`�3��~�o��l�EM�@������-,3c�Ҷ\�@�q�@��L��c�@�p�Zs��Uť�BS��T��Ԟsf�Z�������e���@pG�԰e3�ɚ5��;5X��������4C��\*ѻ���|�q��I	o�˶��W#x�u��/:n���/EL���m"4�qP>��F�d�j�P}H�D\t⟼��6�nЖ��t�;#��p�"�cGi�/� 0�2�W���8jک$9�w����٩nm�U��m1�E�\�ˎ}c��^y�M��\շVE��tf��v�<td:[�E��&����Ԧ6���%������4�EZ��5X�6��]�Z��u�W1Z�~���T>�Sn��pVt�=
0a+��e)yX�(�{��Y�=_{��e݃�z�&ʂ#�K�EyG�*���0��}�#��
w9z���	���h����KYWW��&��e�
\�(�/A�V3��QI��<���K���}��G�)R��ջd|����~>ۊk���h�b����t�b$e��)�y>A����?:HYd�t��O�G��TO#B����]�m��_���ۗ��+����a3/\%�|*N��7��l'0�*7�����4�-�r��ʰ��n�Y�)v�p�gD2�p�m �
����q�{*�p���A�����f�@� �Q����>�i1�A���#���wWF2 n���M�w�[v��/�������\�k��_��a�����Y���ʹ(����i����Ra>	�4 ��g��T����b R�񤮘�ɔ�� �	���c��2	���r��<�����H��* C%��.u�ӠϨ4��cNa/1ԗ(s��#\�0!���%�a�+;�/������7�7�v=:@O�ldo犰��g!����ڄ^�.]��-�w�`�^7�C�!�]ֽ�9��o���f\���oA-(׍Kb̟X��*�ȚWui��l�^�ɾ3eG�}p����k}"��"es�qAQ�?�$�川�Z�'-6[;�H���θ9=��MS�Z�B��Z��)&�6���-/c�	6���ŶA���\�|;Òy��X���,�442�����6�SQ���;O��;>��W�@QeЗ9�v$͸h|)���It7��(P5Urh��8������A����PgUF�u'=����~%�U�3�)�6�2�Lp���~y�˧�^����Cu'��CH�.�ş �]��"��
K$�H0(?	�m�=��n
<�$+�u������+�t~��3�BN^@c�7�tC�̋������R�`�k	��i��j����l$iuTR �- �e�|n]��8E�]�/mp���6�4��+�$n"�!F3�i���۱������`q�E!����&�Ts-�]4j��mY����E���zeh�wU����\���%�&��0�����t�\F��I�!�����5֯* ������K��|*\'#I�F,.(�}�@{����[���p���Y�oۚ��e��/�-�x�	�7}"�H�ظp�E��:u��@�?�g��!�O�o����n��Q.C>�!7���r�;h��'��T�~����ܸυ������
)�/Y�k�t�9���j�R0�=8�Ҳ��yk����_p���X�Ս�Zo�p�c�tmV��K+kU���ZCK�L��ImW�y�K���A��w���`��A������x"#(�TC��?9�[ ��J���FIGK���P����T=����֝@ˀ�U]&u���B}�3qsD�ҙ�[D�rݯs�Z9���ө\R���[:�V���Oag%�;e���pE��Wf��z7-�K'��^�	T���O�l،l}�c2���*�z��D
�l��6��TV;�(L"�uW���Y�dIp�7����%cu�����~*E �_�G�yy�z+��/����)#V���9
s��fI���V�!��M�a�i��EJ�7��62���jp�'S�'^}~.E�/���#��Ob$]�\-c�`����㷏��VE��o�(�3$����?��1��F��J�\˔�����.w����?ƀ�A�N���>D��7d�~'X�4���4�t��>���xj	e���;ӎ����1ܩZ7b��\I)�PW&(i�f�N� A)<�;�p��ܟ1A @0q�v�����6�^���$ݠ�>g�E� �<�Xǣc?�}����,����}1���Lȓ��}�:�,P�4Ƃ���.�ߋO�V�8��4�_ble�[ �RR�j6�5!z/ٲv@FsF��u����̾���@�l�;�X���F�<��F��Л_�kϺ�ș͝2���u!�s��v�� G�g$�!L�^�����u��p��n��2�J:=T!z�X g�:�BGf���F4�y���fƔm��_h���b�E{���v��MU�7�m�L-ݚB	���F��ǚ�/n-�X�Q�N��<�e�`������?��z΄U��|��uQD�U$�z}~�`�~�⍅�YvYN�냸�|�!�e�Y����`�U�W�ֿ�}�jpc0�.	��rs�l���ݜ�RwXN>�Sp���OZ.({��;��'�mN�CI۟ ����䆭�"�xΜ1oS>[�9��m�Ș���]������c;[,�XJm��S���X/��B�f��/��u�Cf�0�]�h�j�t�^\�~��Z�E#L>����� s� �LhI𒈖�;���ts�&����M��:��;\��,�®X籓7ݿ��=w�L�G��i��w�(�B2����~�#�!��)�_��cЙ%���И}8{w��I$��9�U2���N]ad�=�{�hʣR�� u��X�8�������@v�vɧi�1�o��K�,:}k4o���,�RO\�����|k���q�͙��Pw5�m�ﺗ�I� ������`7a�mt;�t��m��a���w�R^2Ɖ��aDi��!�a��%���qJ$�Y��ֵ9��w k�f��t�!lNBh��)��p�T��W�F$v���x�]"�7�i�j-s�[X�-j�e�dM.�b�~bA�>��B�*4N�I�@����[ΪC�Nri������NSw~�W�&�l�h;�-�g�+ő�V�����0�:�ǖ�+�:�ϱ?�wU��<_�g�F�� ��`	 !��.F'e�~�q4���6 �╆�|?��X��5R�ӝq=��+�T��:N�L��0/"<;��	���~��5T���M�"�{h��e��F,�ߗs9�Ɣ-�e���I�4G��tc��B�G�����#8���z���t����w:	�ЅI{�f9��f�&b��R�b̓�hU�߾-X1�q"��k!�f�	!���'�=�hr�]ΰlXٚX�V��6V�@(4������E�����q����6C���C�1��F9�u`�#>V(���5�^8� �,��moW:��ֲԃCh�J&9ȷH0����"�%Yw��}uZ	G~�#j�п폚�F����avͼJx���y���,ˎ�m0#�id�D��$�Y��my�*�Q�
K�ģ��
�,����t�xI�-5��ڰ)!�.����o�%�=����H���� ��{
�s�����_ۯd���>0�@0��g}Š��X�탺�NB�M����Q�H��m�KɁ6��%f�s��f-h��9���*��̢�/5���ѳ�U|�)Wy=t�%Qg2����c�V؀���9�q�CX{��ѦŘs.�e��h��r���!Ą��q�ۅ���%���McC�G2Aa;�tǩ2PT��$������d��|����ωt��:O�
%�`q�/;O,�aW�헉F��;�m�)a�6]>��@*��p��NΣ���yLJWT`1XP$��9u�\�s*7«�$i���:bK�{Ψ�E4};^Y� )��e��1n�Z��7�FY��wU�8Ŭt&��چ���M���Y��MO%5�L�h6v�u�Pꋤ��]��~�����wjlg��ꈡE� g!�:`M~=J�nf��hB�����E��b����"V/�qR�X����}��Z��*:,��1w��,�L~��;DO���=�6�����j��u!�F����mKx`��l��"���ܾ(Q��¿���PP��	����h��mU�7KQ��l�Ј4�1+���ӄSń��'JHX���;�#��u�"���J��U���.��<z��k�.���n�{5�9\��H^%��V�İ;�5ǆ��I�E��^l[	��V^��������|�����9��+/�E�wX'�b��s$������/ޯ���~�S��� ���p�˿|�ڰ	<�~�O����0+�Yx�c5�	�tr?���.R�+�ɔ_F�M���*� >(�@@���_�D�>�oX.2��_�=�.�05�-��%MZ�P�X�cۑ��n^OVxD�yZ��}���>�������ݒ*PZ�)�-�86������66��I�vç^�t�$���e`=-.�_dO�Ϻ�}�'�ך�� ��L�Nn@>[�	�$Y�5�]����:,�_Eyy���Fw�mgG�(�Ģ��n
� �A�VQM�14�����m��霁/)��Q���dpi�kɖ�)���Ȍ�o}�N�;�ι������Ս+�����!%ۺ�=���\#��ṵ�Y�&��(��X�:��;���aS�a��U��G�$�;m;���p�A�7K�>`�]%��\F^1flz�����bFQ%������1�?v�����^Y��b�<Y�C���8��\ïm�~_��E�2��1��ڢD�X�Ŷ]�v	_?�֬�!����X��Zt6b�>L4�!���?x���v[y�QY�b&lA_����Q������4����1-Y�zQ�9O�%���?�Ӹ�(������bݔj!��^4.���-�^��k���e�����,kf���,�μ��ōKG�h4���=l��.�����r���<]cI�EL�0���խ/K.Cgŋ�t���X{Y�7k1�Se�Tx�	�ޖ 9C+橽�'��0�8ȅ�;Y���`�O]�Վ��)C�ܓ�o�K�	U���@�Ȅ7���FD�^H�%��A�"W"K���eKs�]���ݻ��o^m��j��〻|+�,��>��iw�����0i&.]��G%T����&�v�\k�^���;�bO�E�߳����%ml%\���%Y�{I�Y��3:*��ySl��M��Kx���4u��a��y.���_t'@�P��Q[h�~{v�H)�Z�2�k�{��KG�~�9��9v���V��}D�3]�F�ǘ�uH	��A,���F;,����{D=����{��s_go�4�f��+������1y���ND�*�����k��Vs�H����}H;3�&%���!��FZrO����q�5�(r�pg���� ���5���/���"G��T��_Z�Q!V�Sk.�B���L��R�)���u�"�����K�y�N��Y{"Ŝ%�"�b�N`Yܘ�X#��j;㛢�Ȗ���Ӈyt��C�ϲ��g��q����`ƾJ��Њ�i�Q������R2y� ^-����<�v6�I��U���<��U�M�����ۦF+C1�j�wo�o�]#s�Y����[��W��}�_{�9B�����M�EGAQe�{���rRԿ��=Q`���t�����jB?�2G�E��%w�M��a�,X�hy�on��_���}������/�{pF�~
��~Fa��Bf*�l�5h��&���a�1����:�X {���-��m�LΨl8��������K�7��RѴ0�5h�09�m�zHV��� W���-+>�:��Y:�C���t��@�	d��vۯbX?���B[�yo�9��g����u�V�څ�|���ř�q��;8�d�zy<肳�`p��E}�+c�ו��	٨T��9��P��K�+�T�o�mni*��n���^h�����wǆ���6�
�����3���m0{׻Ol��	��6\���u�=b>"1B�n���l��x��`��l��z���p�I�Iy5ly���/^O��'�&Iv�3�1��6[>|�f���,�=�MI�Z�$�V� @~M+�8�`"��Hڢ�sV��w�bR�3�Ϡ�4�=�rd4ۀ{6B^�JVZA�t*۩z��[9�Tu3pj�"����I��_����'�����ɼxPބuz��e�'�D�p�P�4W~X�v�us��:p�/ކV5i�X0	�W�Ga��%G���yN(R"�$M�Y*��mO���T���*.`3���io"�>!��W�� �_l�dp�:nB�h�H��U8���xɟ�/�s�"�����q�|v,��h��7/�c�=Ck�*�J������iD���d,��8�����\W�c��|:�>S<B�v�.�;��U똼���픈�jb��z{p��L]�Ioe�锳��Z�!:X����k�B��d���=���6j���[멕?����J~��s�1�2ZIto��"7�)�������5��v�!�*yP�S�Y�����v�3L�U�.sG�^�)K��#�s�U)���� E͢dE�N����e���}�������Ixh��5m�L�uߤw���$qO����N�lAEp�kvi�)X�(��D=d�R$�p���65�1�V]J���)LV�(0S�yd6k�"��%п[X����D�tz���<�1d���v�u���q�>�V'��{6�9c��F���\r{�si�m����2���&;A�,[)jP� ʴqBe��V�?�"`��r�d���A�ܿ�[6�w6l���4���U���[�ĸ;�O�����WT����n�� Y��l���� B�iL���~�9�{�K�"^�*����l�m��g]�F�EWL�lY`C13���1�&A�J3�+���W]��nB ��6*\=<��v���d#I��FT�f ;g�y���7q�]ɏAl|DEU�?�k�p�~�Wo�
�%ym��K�e*�6�X�ێHj�X2�t��rn��6p[=ޠ�窒- �T�6tS	�V�����=J/ �O�%�Ju�dv�t��XCG�q;�`���;��R{}#s�w�W�����X�����g�U"�tC�{Ȉ���nh��$�Q��?q��*$*6�S�G������WC;*'��Q�G;�x����K�v�ӹά/���i�mI�z^g�}V�s~r�������xcѩH��㚿�`�	-�e[c,Ȝ�� ��8�-�-uc�������~=*�s!��w�24I������M[�Y�����9��P*x{�����+рў{p(�[�vc9��K�L�6	�ci{	2�� N}��Ky��q����\�������ӽ�I�	�eiSgm�߈�@�!��b���k/��i;>���y7ݬ���̏��k�:�~�	�&�w�%�"m#���l�������3g��yWZ�[#�7�Yd�<鴏��M��J�?�K��0=���	s��Z+�^���B��M�;������Y{#od�wT���l%��6ɿ�5m[�M��yn�r�m�\G$��d����dy�����H�E*�*	=��>Gb�ؗ,ؙ�Q�H�R����,i�*�j�����`s��`Zi�n�aS���[�7U�C�qB�ՠI�e��<����3T}�_�M��$]Ÿ:}p�e@;�=���&�ѯ�g�I��<��j�b^
g�Rs�iJy��1:�9I㪋_B���'��pz�m�ʣx� #Ψ*_ygGܡD�<�k��as�k�Vp�W��Rzȅm�{8���U�B�{IX�%D&o&�]����PE�F�Ub�R����{Oy-�]���Z�������K�h�.�����Qމ	�M���R��J<�.�W�ǔ^����R6ᡛť.����E-�I3�����K�]�
�⇪�!!�͂f1�kI�.D�Q�ԛ~�!Ki�0����C�ٯ1�Xǿ/��%�;���F�X�e���7�5� �(>x6��L-�-�͡��t�G?WGj�8�7cxQ�;�ތ��}� j倔�%���U�����v�A>P�Z����ٌ	��>�dڐt��?Qո�I���s(��<�R}ā����Xy�k� �^��`��!�.+(6�P)WZ���;�$��.���3 ��"DhS��U�$τ��.r%( CD���פ�ƭ��iNk`����E�����B�ͅ$�>�[�5ap�	�����j����G�*m��)FaH�����=J���$�*h-[��ȫ��� �탃E����l��A��lu�	��q%y:YRΩ1���d�o�x�t6ۿ_|kl*ج�1	A���=�N��;�%N�{�辇���K�Y|-,ƞ)��l�g]7�?`PN4lİZfAP�_I�>a�!*A1�DF��ʓ4�7���N�i���X�Z�/�����gl��=�y����w������\�G�j�4��a�f�_|�( v�	$�m��=Dg|�Fo�ߝSj�P+�[��QPב��E��bJ�C��Hw���Ja�|1���vPO ~�ZcI�����������3�����ip��/e[B�!<BI>MRW���z�[p��i|i�zQ�!`Pgl�!6-@�����������o���pkU}2��ɶTITm;��J�[�:�(z�<[RZ	��������;�-�<S2��F��An���
D!xۚ�\z�aE��kx��]�}Y�K�~�N�4U�jE���Ut�03������zve��}~���X��I�$��1u���I3o��	W.������QPa�2 ��<�j�r����̦��/	�G$mH)���k�����l��VKmv�~�rW�K�fn�;�8	�0�Ur�6B/��$�4�9
$�sa^N�#9-��8�5��r�������a�_�e�< �Cd�/:0ӦƸ�$����N.���F�ZcOcbr���R<$�Ƽ>	Ɛ��{K��PЫ�-�\�ʛ��ZE�}��X��%�ݒ�V�QL����5�)�zr_��� ��E)8IBJ8{
�tg�r��(E4&=���@0�@����������[�)[�EK��zh[f���:�	Ś�g���댯篼�1��\�0U�-�,d���	���])	j��,0+�X�s+cp'�7]�=�a��6��4�/�������/�$�����G/��	&tֆ��aA@x�"��}{9���wmT�̮N 
l�ΰ+@��ņP��Mc0�\���"��/6�ή�с	pV��kIV�>��R�4��J��~�:��NvR�k��	�R�U�~�Ï���'���rs��lSUg��AÕ'�b�qy���K��G�c��*�g�}>�gX��w�hw������+Ä�/������
�%H�*sy][|�]�P�0ؼ��rS�'z*�
��Q	����(�v�!Ժy<�S�K�|e�uK{�����1�d.��m�[��z�F�⭶80�#�5K�]��E��ែ�?��7��v�N �w�5����,�r�$l��H@���'%���|��G�SK����:[O�^��#��Um����֡Ɲnf� f�i�BG��'P��z��N�(RL^WY!�[ tQ���'!��	��t�c)i^��~�GHq�PI�i](g\V�P�[�X�MC+e��1�|{���RG��>�#)
_u<�詪N������,Y�Ȱ&�{���� zB���gO^!c �Tq���>D�2ʯEm����+�������m�>��bb ��x�Jc�%[Sѧ��>���ß\�O�51�?����# +I��jet~�)�6ٽ(cYg�HzT�(*�i��e��-�^��\�q%��{h�D.������ԣ��hE`���������*��@�Y+���I����s�������C��� &�����Z���Fr�=8�q�I�?Q�U�*�XC��vj�*#�6�l�y\��Ч1��3bb��Ġ�ל������o�N��q@��G��ܸ,#����eC?1��n��W`C�p�旃DP+��)��5���Ο�	D�%��&�l;d�dzˎ�F3�LXA���^V���r`�<��G��� n�>�jž	k�?;��hЊ5d�(i��nB�m�s���T������^�PȊ��X?*fypf?�U'�)f�FN�x�׾m�
�A|% ��@A;eR�3N�ǁ�b�\/�v�,�a��)���p
�ځ �R�����
[K��FX�����ƫ����D��r��rg��RO"!5éZ�[�x��h8�(i@x�Fo��%��d�s =	#Oiq�;�`��Fp��%~�i��a3vC�� �':�:t�B
����(�^g� |�J��s����M�n�Gc]P,�"+�?��M�;^!*7�n�;j���M���&6:��x �}i��,se�QUF.ZU�x6��P�'�Nm��������)��������띠�4l���kv�f�G��ϋiM_�@F݃*������ӯѸc&S�~;�l"T1�������=f�/��u~bz��1}��0�0NH"�+��2.� �<I
��[FW��
ʨ���� ���`܇�Wh_��w+D��=�6ℇ�+�
էj��%uhkk����TI"�$�!�:�!�a9��p�Tb>oj+cL������6�@.�]0���7�5���8�c�9ģ[DA�㪉����x�i���8}��~�r�=r>����8Z=����/GM�t�*1R�ksa�k����ɦ;K4�*����ِl�r�*���,xȥe��$7��\�8�	.�M�9Ґ��Vz���}��?oϛp'�ڣ/%sp�E�PB�C<x)7m�\�K
����r����/����E� A�b���g�4n"$�L%oe%��c��l+�S"c<(C.=ɀ�Y�Gx�掫�d!6 `��8��{�dF &z�1ڏ���7.e�"��!^n`�� ��+�l?6��eDu�+�AT ���z3�����<��&B�����M.��>�"<[�s���j�a�����ǜ��+�ZfC�^�� ��ԓ%�S��s����!-|�9zdIoPb|�A��@Fa����R�v��˸���_:�᰿��ۮ�Y�$�?�nsSi�}9k�W7���;+��︃�� j�>	b��V�����5�[���Y��|���	��c�%�+cp������?l��L���B	�~��~n8��.F� :�5]�{5�����aN�O0Q���%�Y�-�<�J�G�Bǿ�c,b����ݖ�F��o�kBE��uh��f��Z�R��@.�
\��]ݡ?b5�h����W�m���`r��К8)U���f�=�����k�C��D��X���VT��Q�#k�J�չ�Ȏ�"R�����}k�]����Ja�D���ܓ2�c��x�w)�A_{;�&g����8tH���nI>�Z��#<m�\`8���{ԏQ��2V��D����'��N(l �7|i~���+�'a0��S�N�5̴���|Zc�r��F�Z���!! ?�k�:��a>�S������[�:|��v�K��
�3�Ld��:{iQ8��ў���؜�JP�D���G2��؛*�u����/N	#�k_53?
�a�us杼�,��A���8տ2�i�K�u����2�|������[���k�*�Ǝ
ZB
���ւL���N%N� �G~�{I$hO��]��g�/�j��*����\-	�"bWy���2ev���#�m��mt8-�-z^�#FR'�;8`>��@
�-='!G���v	sE�Y<�h#Of��Pq�I�$��#�sv�v#���9骕�a���nv�N�NPX�X��z���H��õS�V�: ����J���0v�ev�<"��_"���ݲ��Ei0��^�M�|�=��7��ub�dˉ�<��[FU��yH��he�ˇQ	s�3�B�2�ڭw��O0�S'Zrd��v!;�������)���t4���U���~IP��7�c��U�B�=E�����$�(�1���+9�d�^n3��^H�4-؉�ЪF?ґ��W.�2�g;��D�Dk��\61�����S=���:KՅ���X|�
���<�YT�#��;�4]]��X�\��+��o�Ӊ�P8�Т��I�Έ�%u��k�*֖ˎ�2�����٭�����s3�3�}�M�Wl\0�Z5X$����aw�Bb�zS�*;� 6QH�E�9�@�M�+�rWP.�b�0���^��������E��pV���u������Z���@4SS�8�ARI/��+]zHi�\A�7A�3�pL�In!{`�d�M��d�8�6'pAC�
����:u=�X��rj��Pĭ�,�%N���Z�m�SEʇ��c��m,,8͂�_D�<���Ͼ���w�����d�#���;���`���ZDi`��3�v��D5L�z��d~��;@�1�q�:�D��T[��-���qqA�n1Њ��RGꐫ.-.-?!��%��Tf�n4q�8�U|�n:X�[L:��-M��	Z�|���)�S���>���Rew֚3�c���:釈4�;���҆���!����Z�٩��)#�iG�b�q�8�_���1W�����v�y���0��G'x�J�,��}0����?&[S��؃��zfG����^(u�I��O$7��%�Z�9t��B�cC�;�Rύ��H��>���V�e���A2�dK�Y�4�A���W��ү��q�0�*=��O�o�!�
9p�i��{����2!~xk�v�v���V���1�\��?8�Q�Z�UÚL���D��B�V���%�M�%��o����LЯ&��������$-�h��cu��h]�S�����>��<���r�����%�[T��Nm���rDx֜(��}���ݳ�$Y�س=��L�*����[ہ�Z�3���9�e�!��� �P���%mc��k��)���M�N���lu���m����g[�*��^6&z�Z]����p��L��TE�˛Lo�u:�<}怏�Y�)�����Z2>�$Y��Y�\De��Y�h2/�n"�ݱ=��H!=�N���|f��M(R�x~ښ�=`����QC��)�3�o
�ԭ�;�=S�X�yvC}��*8t��R"j@'��d��s�౨��?�+���y�\WA#�U�s����5p�o�|��e�
�DZI��$��)B�����\pq精~[%?�d��h��v�(�]^m[���uhs?m������#�o$T��ٜ��˜��(�\�*�FGG�~7T���:M|_�# ��VJ���������!2��Bɀ����_�x��а�@�q�շO@�`����`�^�
�)"��9��B��y�m3~�~C�&�N�����5�x�������?�:q2v�^������̲�����@t�8�fi�r��E�Q��T�i���B�2������4�w��z&�I&����ǻZ%U&D6��w�̭��\_��8z� tN�'��x.��c�	r���o�S�t�'��PKG@8�T!��SPc8z��`>1��,�x�BY�.��ѤL�Y��Ϯ��j|v��֚W�^3'���e����
N���R <#w���]��M��vR����ky!l֜�|�Re��c���ͬ3Py���A��Qۭ`}��)��1Y�;��(��r!��0�&���8Xk�7�t�=�,��N>�E]�!vԤT
�qx��� �i��� q,n�f��d�q��-n�-�bkf@7�iq}�E�^���p��?�q��'TBC�r9����z���������A�M�y>�[�y�Z�:|Tw2�]���Q&6��O�5�Ip�����`��C����{���U��r���D����� �ȸI����t�(�k��[\���(��l�4w��ɗ�^,�2'U�a�ͬ�rjС���Gqr���U�| wI��$z��֮�5:�T^��f�ry	��^�Y�<_��L��bbz�Y���.T_h���l]��}?���+��7&���fȱ��c�$�� ��4��	/�W��0�՜�۩���\c���O�*��6AV���n�� ��WS�ՀQ���y�
㛻�8��	 P����1<�xWܵ��"�f��F���i��Aڕ|��7t�O� ��]��M�nI��%Nw#�|��:�e��8��p�(�}��{(��,W{w��]q��ZS���эH��NDS��8"Gl��Bџ�?��<q\�}�_�%�j�>��l����M3��V�g�S<Ղ�M������̟z݈D��?0:T�8R���0T6��y�&������|�95`��W\�\�i�5����j-���'�C!�� ��q��A��cso�Y�q�L��,��+�v�og]�eEU<E�V�u�H��<�r'��#L8��Jɘb����0�-��Z��-o�%�S��qmd{�er7B�B�/j@���0� ��ۗ�������p�Ą$& �tE�)>� &\(��\�Z�T�Uڈ�[�g��o�llD����%�d��@����{�)�y�T9�����������z�G�H�fN'�T_�t���E���.�E@xǤ>�߶��ʖ6!�P��9��r����1�g��0Vߢq��9hU��6��o}Z�a�����k+�('Ff�<C��w�T��V�Fuݹ����?Y/cA���h�$UU�W���ڣ���2S�ʝȴn�~qk���B�f��q$�%�8���VՊm��%ju�Q�dA�����������C=2��剛�yt��͏�9� e4�T�L�d�w�	S���x5�!��,���҅Z���lV�W1��{u�����K��a?e�~��^��栅���>��ܯr�e6@�����]}��eJ���.AQ�����JR���ݐ�e!�~��@w�*���s�	'Ϊe'*��U�Ѡ�Q��i�A�g���������6q>�����K�T,s(ID�'�ԐǠ���������{:DC��2�E+Uq��R_��� �u�A�~)�W��L}LT���u�ؽaB^�Ɨ�7;�у}�5�U�)�d��ʛ���4�]QS%�پ�c��;QfgV���^�'K7�D
77�]yk��5�
I��� �C��!�h�o����E$^;|Ʉ�e*��|5�q>XԦ*t}��p�њ����B�b~/w:��Z�ym��5���lqHz��]!o3<�ˣ|$��Y��=Y�OTr6f�c�`6mA���B�r)i����H�~���O��	x�`��(JG�2�� N⃆~b�H���u�D��l�0P�)!�)��|j`��@7��Q�p�)`Z�y������1��˔�Xq�Prn���Җ�����v�WK.{b�~�}���.��N��s�&}>j��b�z����S���'^3�Y��q�D�;!�\��W�j��N�h��'�v	��!}6�"�R������.[R�:[�&Ԁ����M3O��)4�r�7o��Fk�V̒�*�j4؞\W(���B׋�\N�\* ��H�N��˓j��G!7o�;�R�z9fb�gpH�AEi4ҧ��8l/��=_�(:��յ�#��x��_IK�';���:��^
$�< }e�,S�B�K��#2��b?<����`?�< ��K}
5��r�74�@��l��,�N��� �wK��e��<�N�L3��1�S�.Ҟ4��ҿW��Z2�rp0W �����̏�(K�0my
��s�QBF�	�eB%Ir6�,_�닆�l�8�o6DY�D��j�4� "�7_�<�2�*��|�Z��^��9Wy϶Y�a��Ϫ��`��Rb��V����&l� ��:ٱ��q�hќ��������#�"�s���f.,�Ӑ_�Cl�^�z��c�fX�" �_y��Ȏ,�&S4w����޵9+�/[Rˋ��ƥ��i>̥��C���Q�el9�2�(�a�j�M�󉱓��.�j 	G�}C�߮���vo��;~�23j�K���y��:�ː�G5�%��7 �ۓ���u��&;��T7�'��Ă��΢#��<�ԸK8��X�� c($�첎{�/}v��N�+H-w� M��Х�n�A<jM�Vݱ'��E������[�"�۽aN)�ٟ�yB��}*Ne�'����Yx{��KVNv��n�쐒Э�+�T�F�{i>�'42�Q����ҷx��wˠ��QGk�#�Msr;d��N`�n��2ݥ�������v��<@f�����Q��pR��lzuC�?7DV�@P4���y���&�Ӆ��R�^)�'#S!���j��Uȹ��ct
�\�e2�(?��(E�е�������A�8BlXşĎ����������r�L]�4x%�,�>���������W�A�FP�Rp�H؊��qU�7=���vi��"Hn�ukPK�R���o�Qn��c$�l��e3J�Iӧ�&��u�r��Xso��<`��f��<�`.�)b&}`w֎6��|���v*q1�Aʚ`�M��g@h֩���V�b�!)ӿ��h&c�ѯ4�(߳��=0Z�m�=�䣧J/�&x�-�Y���/�ª*���ďv�>��d��B�A��ΏҌ�=�5�_� �7^*��ˮ(�)ʡC�%b�%$%p�nk�f|�d'���1���G$!�h�ap�7s�2��@Ǘh�a�x�
��y����l���j�2v��?uH�_�n�� NY�/x�d-��_�i@�ǝgv�*ŀ�E��(�d7�V:����(���S�nv;�����V���8����^�30C#)S��{]�}/�nH�u���M����g��W��9v�\�*�~G���a�L�7���t3c�v�K��y�J����*�}���6t����%�ٯ��o��V��eu�@q�|X����1haLJx����* �}�`�f�[��6q5��S��W��9H�u�V1�06ѹ\&��`�[U��	<i���G�]�A�)��=��M��1���]��*��ۂV()���[406�g�:wq>���B���:�)2���H_� O; �8��k�{y9�>�&{)v�3ʖ�拏��@����.�wj����ɻ����	U���9�'�=�?׬�B�%:r�+�쮐�����z[����p�E���p���&�E�b��Ь��=�b�P���X��ى�"�t0<n�eU	Eu�W��ғg��9Uw`��/��?ἡlS������?�J P�VP�L��^=#8������qItC7�78�,��,0'?�t,�p��S|aRt6��$;LuNweBVajl���L�w�[)���pA�Qv\��9}���q���"LG9b��bR�Q�eٜ+�;��1�⦷�b�B}��;�	h�G%�����M)�2<h%�lz�62�6��vؤ
B�9g|�#'j'������������^���P�yۚ:������H7���k��C�Ѥ��6 ��6�����E�Yl��glT@Hh�U-���K�ۖ	��7"����Hv������&��po<�AQ��ߞ�c�hˡ�U(�o|�3b���#�3�JѶ�ж=��w�(�UF��\���w"�S��?��<H�y(�����j�D�Xg%�݋��9�/D�Y#�Eso��H�L��n�+M�Uo�df��:8��5�K���5JP� ���[/�A�	�/�!:%<���x.9ݱ�s�o��Ў�k˗G�4�X��c�Z��|i�A���W�>&���4�Hp�V,QwF�bX9�Ks�� ݆�|/�H#�>��:��o,����5y�y���R����b��UY���%i|쁇����"�G��|��W�+j��䞐~n��_�0[&�BA!z��*U	�ظr�w�l7�2�X�,�&���75$����A��G���u]�������+5��G�F����w��;����Wf
����`-��EJ�䙍����`2�"�.�]+�oz�����{]�XY�i��Dͺ�"�Io�W�2������!L� dy�EFƾ��U�n�gy`�@��(O�l��ŜH�{�On;�
-9�˃����]���چ.-�Mb��6k�l������,Q�خ*ff��%�&c� h��f�Ɔ��)�]�wg����kq��`8}�/��{��N��wGهƄ����vK�,Y�mm�@NA�����^Pj�V�Q!+����f���/�/��4V��K��A"�� 4c��/&-`"r�Q��a�o_2������?�8�uv��2���MR�TtX3�D�:.�k\�Խ�b�1���0��>e�d�(�˰�O"����oMD��@W.
p��g���n�k3�i��y�l.@�|T!��Q�.0����g��9�B؈x�'���l�]�ßrMR�n(��l�6���*FK�}���I��N�k�ܡ���U�Y��FP���V� `�`T���*Ж��z�R_�sGi��1�C9�Y4̄1z/���I�i3"RL��pRW�b���tlu�f�C�k�����~�x �LC�=ީ.A](G��{�ۑ0h�E�Vf ��zV��Ld4��JJ ��-��g�(	w�ԟ�ť�ѕ����
d���累�k�`�gpw�:�`���#}�/C�E����\��؆ai�#܃�<O��@H-r$� $�b�q��x����x�1�k��Y
�Mj.�t���c>'�5��z�Bp=@���=�"��J�`A���?�NsS�Eؖ�;�������v�naF�Ιn�b*1����I��7��/~q��{�u�W۾�{�1���1 \�6|ݒF�Gw�l�
�n7�;,, &!<� -f��;9
'Y4m���,A�Hp������[R���;s�K	QM(��q��4�:�X�L.�SN�r��~���\�F�C��e�7�`��_���@�$幻S9ө>]��D������]4�}'�<�W� |�!��	$�`՗�=�S1�5�l���>b7I6�3�^��%'��dc7���,#dɚ����H��g�	~z���4t"[�H!"P���}�-��QTs��J�7ߘ�o?]K��6Ԕ�=I���o,��@{An��}b5�/�b_��j�F��5T���I��=
�>mB�ͮ�в(��u��rF�ߑ+m,m����ӎ<���N��|%�;9W�Zk��w���G��ˀ�{�� kd8'7�\������Ϭ�¶~Q��;����d�Y��x��OKi� ��'vk�L`���+����/Vy�S[`�My�SG�:�b-*�±q����%)\�Խ�si8�SiG��M=�?w�B�����~���rF� �M�?,�;���_�`��T�|Ʋkǖ��C���`v�-wN�ÿY a�7Z�	\�����p��ҝQ�	X�Boǘ��q����-3���]`d��3J����@.�LE8y�O���^Ua�i-��yŰ�o��5u����U�/<EoW��a���]��Ћ�n�n������.��m��Ӵ�)+���\��Y�ŕo�V Р�*(B�7\i*BB�j��/��<zc�kH�{}Ѕ{�Of{{�� ���QlNp��.�=J�P]ƾ��*7����1,�{�yr!�{?�|3Ϸ����b� ������ނD���e�d��̊T�3d��0it��;+*9��5{�a2:h�b��	�Q
�.�`]��tw�C]�43���ۭz7�z��Ƅ�jDy�� 뤳���1Рv�ٔ<F���*8]>b��h�-6\�:,	�7\Մa;�ݮ}���Lv��iE���a@$c\��խ�������~%��IK���i8UL���I���k.*'*b��N<�Pux�Hv2|�g�~I4��yU�>��va�QY��/�=Ϻ	x��I�vQ�4-RB6��UG|*�KR�9i]H]n����U/cq	����STA?�����j��9�麑�=���U����~%�l1v~r�χc�s�Pde��6)�P��g����S>�Esse�d�{]]�b�[3w�z̫�{�h6J�z�f8�ȗ/{b�<����4�Z���m,�}u��Bpy�	��8���C�fC��vx}_�Bs����Kkh6�K�<�gG�_:^�w��[e:+��	��,�2�)�	(H�n\��J{��H�
_�����{͜9�̊�`�F�G��a���@1�>�F�Z��~<����y�m1� .yMX���c2�ed�R��hʟP�+w�)إ��A�l4���,D�9�� ml��4M�[����O�9�4�hH�?�db�?O��pD����3��!u����>!e�Z�^P�:��O��[&�����w���j ��	��g�o��j�`�c��$���bq���\#U�ZY���fRus��3��N�H����h���P>)�[��=�43���J���p��#������/���b���K� ��F�ǭ]i���z�x�y�8ѼNF.�f�Pb�ٸ�[ �GD����ĆT,�I�p(" 3�u���%n?���B8L�η%�l�1ˤl���_�#��+�L]��/ M�[��|A玢/�\��M3d��h�'>d�^4 �5�m�Bo6p��o��X�s�U�:�m�jCI=���
'X�OK�x��]
�Mo�ovbp����b�)su����3�74Qϕ��(�����9K!�xS�C^�C�$+:�A0:�Qs���>Btvr�R�¤p�vn����8S�z�$()3�Ma���ٴ{Z%���+�J��ĜfHM�h��e(X-Ǔї`įf�ࢾ�H��*���x*��������y�I���\�k<8��j1�m��(S���G�ʩ�f�H��E������Z���ε�`G���q>{H�#;��.Ӗ!F3(��tc�,F0Ҽ�Y�-�/��Q#��F;L3�3����O(��R�v���!�n��--���-��U��R5dr&K\�_r���c����aaD4�̗�d-�;[͙���<a�!c��*$�?�Ν?�,�ZR�ˑ/�P6z�GKeh{,ٻ/$``f%//콫'�Cr'��'?�W\��F �\�r�}N
0�.�����~��x�|�F��8�!�䮊J�Kj��#�<�s^��E4��.��K�D�[�,��f�!9�N)�["��)�~�jD{ ���"\/D>@��Ak���b��!-%��Uj|_�@&ۤe��N��৑\,KM�i�ޜ�a���:���4#��z�J�1�x���(e��H�5r:��'�n���OwϜ�aм}�J����&��e������#�R�������%]�ό�v6Cʀ:SA���7s.v9����a��f��P�B�t�e�VW	�1]~�m,�n�K�e��G��ēy���)���K�r��<:�k�a+Цqw���4�6+��^�j��0n4�;ɏ��j��Kv��'�����_죉��:7�D��@;X5���.q��Jtn:�lϾ�����(��Qk�0c<I���rtZSy򇪍���!�g�"4��I_!��� �磚�r�G�Y���k��ݡᣙc��U�[��[���|)L`�O�'���$�y�5��B�vPs����W6t�cT2�4b�#J`�b�BfѼ�2��LM���xBa>P�h�~�X.]T�+���nF_�;\c�8!�1@�,Do��p�[Pi@R!v5�^'�,!0=4�g�#�R�n39��5���	�f�=uVBp�67}[��p��?��='A�+v%m�w���l#�;��ܖ4��n��a�)�� ���b��"�K�s�w�Ƿq´� ��-��$^���fe��i��iK6��Hwխ�&��6���ӽ�h���a����U������'���k��:]�A�o���:���s�,j��)^������)����+J�d�
��-���0�u=;������h�{���]�V:Uv���)X�:��n�+)�&���e%��ҿ)녙We�K�SE��e=�	�'��Q{��5#7��m�?����hrK��!H�޲(>ϱë��K� Ǻ퟼�t��/@	���|��d6�]n|��XB[U&]uǌ���3^��;��n�x����m�6ļ��
�\��s˚n�y���K��mO.��τIr����_��*wc�	=���!Ǵ�x����#��F�~����`�8	�KT�I@#�,��~P��9 x �����H }��p[�醠�g����$�EZ_^N�s���"\�8�.��)����ry���W�U�_��y}��K�m�����e��H+Hf!o1�葤��΅7U>PZot���@?zJe[��,]��y��IGt]��_�I���b��r�,T�#��so��:2���I,��9��8h�j�ˡG���>�y�[O�Mٟ�
4[�q�ƻ�R<xn�����2��q4��Eqc����U�׬�ٗL�Q�}us�t6?J�P��U<��W�n9���p5���b�Ns!����jqJIk�jz���j���������}�@R�M}X^(�imJ�K�:JN]2���
 E�Z��ʅ�j��lt�]"�e�9���>������K�L]_���N���`��.}�P���z�v7��K��k�����)�թ�K��H��ס�0i��s=T�a�7��x��x��@8�W�0�]d��%�pv�;u��n>�o�������mҎ-�b�e��C����E����4�q{%�Ly?�gdmw騨�;�F٘�l���� �nEi��}�ep��WM���}=y��>�e查�&��n|�-����E���
:,p��S8��t�H��g�
��M�����j 	�VKO}����4�$Ĭ4���jW�P(����j�7�&v�]� �)>��D<���,�h�w��L�(�>����b�Y�p8���w�)T*U���	�3k(r���4U�l
͸��tD�D�5gА�����=��y��񢣭��b��:�_����\N�n8Z&��|�	[�C0nN��+�M�rY�ċs[�+���8M� D�V/a�=~^C�-%����o6ǫ� �ٓ�x�^�Gi�
�:!M��2C�'{#0@fD��B��@n�!�4,��:�0���J2$l�h_�튲�}Y//#��ؓ�/�݅I��-KC���9�}���g�xK�u��e�H�ۄ�!85bB��,6���/����m~�	��(�Fb�X]{�1���s;��v����!�wGG"��*��6�w���?�03��_)� �
�+Z  ��R��Y�F0-{L��]{��ܢ�����7!(#i��MuL҈��L3j�j�h�٥X�R'0ZYe�v���q�f��KH��/��ao�Q��&��
�W���t�n5��g��.�S:�lp��@�g�3j|��Һ{����.*WO9�檭`��Wh�N��?���+�:�2�|��n�H��X��
���@�0#�$�'�c���ܕ0��lu�C����}�&"�d��v�%�[�x��F�Ms��Ak�2�b�7[�����@�o%�t�d$��L�c�t`՗z�ZQ=�!5?���TQc��$-�9톨������_�[��)��R��������kF�BC¿n[��H$3=hfc�E��s�M��SF#�Ѡn�������,�n��
�]�M�=a��3vߙ<@|2rԛ��a>s���A��	\�G�`y��t�x��@��`ӗ�H4��D���t�"+G	��pIt��� Pp��x��y{��a�(�`������+6Vo��&v�]���rI��@��j����Qnϱ��豫�9�r����_���j}��#��U�Ĥ�v����n�ѱ�.z+(�u���c �x�q#�9�g��sre�4 �i���k��Rn}�?�z��t�W��+�Y)��p��wJ�d��Y�X��{ǿ�״���Ѥ� gHC��=g.r<��#����zN���Y8��w6�|V�z+�i�p �#���%��t�s��>?�v�R�o@��V�\+Z�>9�pb^��Dl��FR
�h�]�V[d��^�A��L'P�K�n?Q_���O8�[\��Lz�4jMB?�z
d�H9B7[���x��$������]��~�%���m�16;n�b���O$�[�ƙ/�j�2�㧬�*�{�kR�}x��k�
]c%�L~�ژ��j�J��Y?���\�㦧����:���UŴ�ګ�V>���oF�۪���#�����Q_n	�LjO^[
��ת�wv��*�%�T����M�oR��i�xk�p�e����`BAWߩ�����I����)�r\�����d�Oh!�3�3lR�x�>��%�#o��e�b���%:�-K��^iV� &���b�.�8���(ʬ?BJ�
c�sXJJN�:NJA\-�0Ec��J`��r25��`_�X�aZ�B��X,{��V�+U�d�q���_�Fx�ѯ�c������Y'�F��nq���',�d�6��'��0}��GŌ�$�z��A[uh\E������xI�ף�`��/��ښ�9{�Iٿ���(�A���2U�A��^�;fAC5K�����+�b��8rO �nI�m�p���ׯj	��J�Z�!��&�������#䥖��׺z��PT��?+M2���	d�^������׭�4&�~�Z�zB@�ԌJʛ�%�������V���P��$������^�Ǝb�k�*�fU���#�7i�O�*M+?r������Q�����;�v������ϊ x~��5v��a�߀��1ǹ����s�K���[�%<�1#M"N�| �"&���96T݊j��D(?��J�})��X���� g�4M#�T��:��[ ����Ut�1+��6���Ȱd%rNU>z�D*���w�7�y��L�f�����>�	)���ɶ��d��YN ��mX�%�I���8��1�ޕU�!�ξ�%�ȏ�vS��/S��揽|�8�%�"����� ��U�>#��!(=��ճ��?U�z'�~g�9�U6�K�GJ
�o���2��N �iD�����;y�C��� m���Hهǜ&f��N��=�����^չ��=�2��b�=&�q��[η���lN�c-q`�dd'�Y��ieS�h�㧐����ljD+Z�� wxN��kT.��Z�*�>8[X�z��n�9V����/⩏��O!�3[�Zk�6Od�9�£��3-�B�Y��Vj������� >�B�Y!����7�cOXBgi�K�k�M.4���U���*dSޅ�g+��2nS��O��-�~��>����?W�*2m���$��/nU�h'\��0E �@�F����n&ĘV6�S8"�z�pF�D>d�~��k��w$965�W٪�������o>�;(�@�l����;���� ���i2�k߱>�h���7�s�aum:�]7܂"x|��Iޯ�7m57�L[\�&Dq%��s��Xr#)�4�û ��O��Ѷ�{|X�m4䈜,+���c=��qR��XC��*_#
��A����gw��W��횊���;U:�,�ؖxQ�K0j��e�����t��e��;��*p｠x)@�u����O��|�͜�Qg)o��~	�s��U�_����e{��i�n�$�/��(��|: ��K5:����4�Sۚ�lSf�V��bKj�*|�����j�X��3���n�zE���P�p�\ ��xTx�$�Q���ͧ��$Thv9
w��>n0��!K%j=�Tw�~{WZkl�5����ҵ�dLs����,��/�Ɋ����W�N�e�ÙU�JV;��Pc~��HQFp��wD̵:��-��Ə���]E��:�����J���5K%��ha@PDM��qI��.tKE��]`��-��Qh�!��A���U �;N�׏;�/��V�^��ß���Z����>kPJ:)��O��$Ř�&�Dwz��qb"�v�����N�������>2P lp!e�|�a�sW�e���k�����H�ZC��T���/�J3���V{zDq�(�R�߄{W?_%_����>�������e���hk�}�ѹ�'��5�<�cM�й���f�w��'ʃ�A}�h&�å��f̩- ���yi�����r�H���vS����B#FA�d߁��krX{R�)st�¥���Ŀ�]Ae��2���`���6�f�x��qʁkiߟ��㺽������>�7��3'��}��j����B�l8�����O,����]3�7�?�~	v��v{����j���������?��,$ }'�׽yj���J})C��G�H�қ�Y�������ӎ�g�u��	asZa؈wd��fjPO���at�ej�� f�g@Lh�Λ���iɡ��q��\�p<U�ܧ;QU��XE�Q�}kq�l�����s�m�
?�MG�# ��w������(�l_Ҫ��r��ƹ���14��J����9���J��I9�"�"����z^n(M��g��r��p��f�^�@����HD��z�/ab�_5
���h	{>� {�ҁ�nyϺ�74��xB�ED������` �(�hK����R�I��;�Nr�[���8�9�pP��C	�Ŝ���d�G������ e30����s�oo��o��{��S�Rt�k�Q��^��<��8�A8����x��ER0��t��WzxG�62���0�������޶R\� �`Xʼ9tx��U�q4��F�W�e?=)67\]�M,/*R�p��&|c���ƌ�F��+���z)���#����@����~�à�!�Wު�'VN��hh0�;9�4pّ<�&��W�>��w������"����76�AD$�^a����INxH�jɟ��)�ĵ]W���Ô��h�v* �:�#5/��Ј���ҏ�����ۖ��aw/�Ru�p�14 ���K_F��������T��l�i���~Jq�Kx饇�<:�&D����|�=�e�b➷�p�X.�����].��@R��_.��\{`]Z^�vSj]~����
�\'#oj�.=��3#S�8C: ��$�!{ ��ΆЧZ�l��f�m���+;(E7�V6d8��>?��3�����3[P+M���2gs�!I��ZE�+ U��I#���ֺUT�o*�ђ�����߳�e�������Мߕ2f��ў�T!<��<��4����b�B�S�_�n!�>����yykP�Fi������b��Y쟭�cC���G���=�Rxº6)j9��ݑ[�%+�h��OW	�Ω���4����!"���>\mz���jFN�=zb�KCB��b;Y��̙���_���W_�lY�����6���M�L�
��ڷQ����>��*W�b`0Z�6�6���6QOS�`"wϋ/��,p�Z��4��%��i��4�t�S��>�7}#:�B� J�G���S�W�����1J�Ĳ)�]�1���3M�I��g��	ji��l��h0��������-c%`n ����#M$\Zx=��e������/H�ǈ�:i��
����b0CJ�~l���"vg\���5D����؊�{��G��@�,�e�M|#��B��By��8���3�̳K�V�E��Ț]��s�g�}WkI�xT��~L�v$�B
��H&�}�ϩ����I���ӻ�6EE�Q3���z��)�ܐ�6x����RN�i��谀��o$��.�:��|��;��%�i���8�;��P@�$д��Y2�
<,.�QI�KPay�=[�v��Ȼ�0�M�*nvO��`"��aҝ>��,������Y{�c9�[;ʲ
���I�w�Rz�0�B�m �[���;�Փ�,{��9j[��� G�n����X��@�7�n2آ������X/�r�c��?p$k{!G��S
l
F�$3n�{{����J�q�4����9샌o��lSR�կ ~���1آp�m�]� �@b��./!9�A���L�0A�I������
�[�Tp%��n��)u��`�E��$m����Ͼ|ŹL�2p ���%`$`oك}/��������m����*9]��-�CF������ʮ[kע��N�T0�~㶤�����?���[(ˎ|Mn����X��%��l���T���&Sh�}u�)f��T�v̭�����
 �ܙ�
S��=@�E>i��s�]��󪻵�H�oX��ZO���l�!��! �{䲌3a�,[�F2�'���\o���m����sOS�g�%��������q��4�e�
Jؐ照( �̰m+y#!\ȏ�"�j�}S�*�@��e��&�#.p�Y��@9��欦g[��=�ǲ��0M����ԻTChjڏ�W�4�f�cVv:�9m�G�*���{A_�=u~!��ؽ����� ň�l���^�t�T(s�a^坠:�iO�f���~�>B��򟩩?R�Sk3��-zwutLh� g���"h�V^��w��}������=�4{�ם~�I�l�#Y��u����W (e��_h�u�4�i�[��*ت�6�����0�a�\��̠x=�)Y��Nz��bQ���;(��t �ް���i,�p��0E*�q�6�b;�9_��/���6�5��R<L�C�~B>b�7[fRDZ ?�3�;R��3��/��1�+�	�"��/����� p^[g�RZ��$�����ҋ'�C����n�����b`m����أ�Q&Dԥ)�Agt��#+rhǿ�&��ލdgѲ� C:�=�M)ɕ�0�&�A.}6_��"���B~'�N��b	F�` _z�G<��.�H:��b�^59� -���)jEco�ؓ�ݛ�$a��m�v�T�Yz�Xo�a�
�4� ����c���l���1֟�#�0녷�sXV�դ�=i�Ԙո����1t�e�6�i.|=p������v�s�Dt�(�ǻ����)㌎�teɀ�2e�~Ko@}�'�{^v��r�#�t5b/�݆Q���'�@�\��鿈�u�b����@ը&�NU��'O<O/%�QxI������gL1g��A�u;V� W�7������5vy"�O��x�$��Y��I¨UE�� �iu���y9!��h���╯5X\i)D��[�,g��1*���eX�(��$9f����udw�>�d�� O�{K����!oA�Ҧ!�>cUk{�h�dQ�pB�P��+xN�K���"/�	.���T�~7P���Z\4���w�i؜CB�,����	=k[@d5P���;�7- n��@W赝���?�+C��r//8�������R��nc���^��؈sܣ�l��Rk�0~�T��w��!�3��g�h�����n|�I��ONJ�u��j�dHvQ��w6�S�e�I�Jk� t�<5��OEW�,��dA&������
)U�1��K*�;��>�Mh��������9FRQl�B��P�{��-��O�E�+8��G���+cͲr'rU���g,y���	-�={��"#��p���7@T��3"�C)�|mJT�7F���`�9sdd�_D>ʈ-A��a�T�(`�C��gu�4�E��ֹ5��R��]�[�����#q�@ܡx�(jP5t��V}�L���9 �[x8�H�w�x1�D�,��Iٹdbx��!#2�fb
���yNT2:r>�~W"�I��ʹ���M�'�=:N�T�\�:�e�OT��� a�'�"a?��>�K��8p+%*�@�
��l���';�����B0����lY��tP�a�<�ฝ�0Q�@�^�**�Ei�n��U�y��~��ATu ˦�%��S�OE�}�3�-\����.d�6�`���	,�H�[f��o3��a6�M&H�;����4��1o0�>Q+Y�!�SH��׸Fw�����Õ;A��	6����^��k��?W��.���[x��D�~�9ˤ�M�?I�g���ڻ�D�k�W��_���Hrn��
��YD�5���L��P��8�r�T���%zLihJ�_�Z����ul�d��i�@KrSL����\��	� �n'S��%�66{���3E~ �%{�A�?o�ښ��4tVzt�suH��GB��q^عd�4��6>�(�4��<T0���h_���6�����|}:9��nQ6��>T��A�ϛ���)�a��O���m�����w��v1Aː"�R�-#��v(�J�y1�t��BC����YE�3���ԱR�i'�)Gh��=q7E(�@+li��+��"#EX.�+%ݔ��J88?��@��j�N���ѱ�'�\_Ղ��D(��۵�D(�^��0�4��b�H86�`�m��v�nZ��\r������u�N�Z�����o!������}�Fh?�����P'���}�C�ǿ�:]�H:(|�B��"����G����/��*��:�&�Y{���Y�����\�;��B]+rK������\�	�����A5�'�4):�ʁ�E�g�;n'8q��E��u}Je'@�6�x4<���X��l���bƆ����'�X�siT�� Q:z���#2������R.vL�D��6��Q'����~��u�4�j����8SY�v�ੂ���7fL�#�I��:��F�sY���=.������ �,�8�&,8�s q�qЀ���L/��d���S���1��mE�6(m�	�,��k���%���H�bw�VT�>���>{���oV?&���َnR�-�b���{_��Y
������ Q���j��O��l�dly~�h�$�<^���*]�$fU�o�E�3���_�Z��J..G�^R��
S�����U�dY�.TȐ1`�r�c�E��J�1�"�	���u]݅�`Q-#Џ�<0��U�,��|4��Y�4��p`J��^��GG��W��to��!ʍh��WP��G������WO����&M���-�·�cn1�n:�P��
y�6$���I�c��-�2�0��̷�����1Ma#��u�Z�|Ҥ:���XLS"����8+݌��[���Qz��7��	EG6b�|#H�Ȍ1�#�1?�!���ۖ��1��[s���པBO����R������<
���<ܗ�ۙ� ���'T�WTA���� ���1&[G��1"Go�ƶÇ�b��x��yH\���r��W�!�����WL|�pP�@p��Yѹq��i&��9>7ݞ�S�W��Th v�n5z]�����5+
��DWLW�����~r�.;PK9$������9��vѢ�t
�xG���$�6rX	K�嶾�-۱=��H��!��IxdY��g��;~���ݓ8\Dڢ����ٻ��������+�>�G�5����)�B+������-~���p�bf�_J\P��g�`b��J#�4��Ď暌r�QZF�F����z3���.��«�Y`%$Z�=�tx��)���V��s9��|0�7��h{X̫bx�Ҧ���8��抙qxt��\�s�2}��?��L�`�_�Z}����׈>-�v9�|!L]�ev^z@zx*)8����������oP��3����Y����|"e�w|��>��~�̊�8G��3�[�br�����=|J�zA���x������d�{1T�,�W��Z���	iB��D���u��,*r�SH�E�=קբ� s��-r~�9���XbS&UO	�;��#��aж���3�]Ri���}GF�{OR&-\D�;�"�n��M�� ������G �z��;l6`���K\?����3Wo�����^�	nd�����[!��<�vv�	����h� �Z�
"�/T���x�ͤ���l<^/w��Ҫ��Æ+��xf�{��P��(,8�V/��6Y�.3q�cP�� �p�X�q��B�j8*�zݦɛ\�L;`��#?I��@8u9�Ή��WU�_ȨHow0�}��Gv
u���6��zl'/1?3��Z\��Z��s~ѐ�?�
�H��^n�J�Ebf���N�!��Y�I���c�98��4eMy�Y��<��SJ%	jZ�Q�a͑�j�H��yo~��H{��B�4�;��n�x�<y݆��b�ȋ�-�������{+�מh�!��c%�]}ҿ\��v>27��*c�X�w����*Uc�N�} ���X#%��f:�8r6���J8ܹ����P��{6�/��~*��Hո�GK���ny��R�N��v�F
V�q���CJz0�� �Y:��^��:Ց0��;���C ����q0E�^4��,bx7�&5�ml�y؃�9��������;�>�^4:� ��0�s��i�K4m%��g���u�e&B.9��[8=2�D|p��c��
F�$)i٘��!�,��
~ۃ6]����+�i���I�i�;�$z���t���.��+X���2��+Tn]�~�٪����4��sӀ�]�}���	��MЇ�Ywt!��y/5j$D[��i����C�eJٱ�� �(�I9ˇ��dH�������W�}.�	a��rPE�WJIeՎ��I@�~D�ȰE(\j����0�j���͉��U5��gwC��w7)4ܜ���ŗ�az�W>\V��eN��/�?WKS�O��5}%L��;ڢK�1g�Ԧ��#�Gk�Xhd�((_���}}�h󈳊�8׶�Ќnmx�\$��y���N�D��HNz�m�wh�$M9�U�%s��� �8u�W�-d�}���d�4x�&���·�^�.��;F4���f�r�hc\����7��͍&lӟUY��ξᥕ}���{�߆�?��a��\��GaW}-ah��>��k��_R��;Q���^�Q�ە����bB_QJ�*�cS!e�"M� ��v��	k�Q�2Mo/%�<:����eN��(A;^al=���e@��Yh��d��k����U0`�<{kG�bk��B��S���,��:\ N,��l~�LUh�CVC8ݝ4h~*�9�D��l���V�R��ݧ�g������l�fR{�=�O�:�c���zWww3Ӊ"G ����]U���
��(E��2���p\�`l��#��Ć�JG�� >��o�#k���"������G�8���)�XĮ~n_�z��,���1k�h��p>4~��L}����k��<u�cX��CV|��M��H�.�"t��Es���)�))U�3�K��j�hYP��}iR Ka��Q|��pz��m�ف"< G��ҠsA��"�Ke >�8 ��ͽ�{�
9���P� >|�ʥm� HM�F�k�TG�z�x)�����O���A#7d���v�U�t���w�O�/�L^$i.5��E�mS�f������^Caz���0�-��_>� �W�.]�(��46 �Ц5���E�ՌɁ�kט��V>�f=bhW��I�Z|v*z^�v_�_$�}JMa���G���sݠ���M��0d�	5�7'C��Ep�`{�#�]��t���G&��1����V��Dhy�V|��=�g�t_��f��j����4�V��t^������K�S��u͹�����Ke��Z��e�]��Q@�<Gr3h��RPK���62� eD
t �[��b�Y�wQ��&�L�N��Yy�B��b�c'i����1�Q��1������Е���	��	l�Ri��t!�3w����G[P�Nvs=��~��_j�A5���2�٘��Ŀ0�_�����|���E1z�N��:�>Lyx�&�#����Z�ee���M��&�E!(��5Y.
��9�+��C��Ce�!�1}�t���$�����?~������j��(U��� C],<?[cL"lWɹs���@`G��/Ws�a��G�ۇwfy	�̂��E$��ۅc�R��)[Y+��[>�]���r�����$C2}��� �cy6S�u�Dнe�[*TӃ[�z����ˎCMP��@�A�Jɠ�FKTv�~���8@�؃��q�	�;�n��~���]�i���Q{��Ț���^N�|�4'it�4iʎ6�f��<�����3�XVzR^���5��j��S���@��ε�����		T�!t{c?Pq��������mZOdyV�G��lV�Lm�l}��f.����=&a��Ã�ד7�d�XGq�,�kթ0�i�3��gӝ���]�Q$ M�p�L��D횓;T9����k�+���8)�bf�a���|{>V�>�z+�z�<�)���+�UG���"�ط�_���N���~�Gd�G�ֱ�k�M_�7�J>gD�,�Nm�+f�(]t��TV����l�*�;�,80/4i���P�9%2�V^[�����ICmҖq4��bC_��&8�E¶'[����zo�����w�o��~e6+:�(>pӏL� {����`�O�vg��(m��v.�C�0��dS*�>�9�Q�����&�ތ�9�%)V�a�(������������ڀ���'٦��ߧ)[+�y������ƽ:w?Q�0�Y�ɲ�~����ũ�ˊx�6� �osUr����7���P¹B����3���ĔF%[����Gc�]Q����ڂ��4�P6=�`eϿ���s;�11<��H"1��f�������H�q���H�A�5�� P�f�c̕���|����-�hA!�%c�LP�s�z�W�o�"O<��~������3"�2�@�L�!r�c�%1��õ�.C�Ē��͒�������J�o4x�
�ޣ��!���t�d���������_�!���ɍ�*��
ٿ�IPd�2`'���i$���d�Nu%PI�$���Q���HI5�������d�N����<��_���e�3>�������C���o6�o�&���地�rٙ%6�B��\��yˌ��p��,�?.����ZXF̷�������F�:Iƀ꾜Y���<̯�g��-�d�ׯ�#NT�|�uTN���ї'}L�!rÔ���tJ~Fl_F��0h$`D;i�&�:q	�$mp�E	{��L�Hmp(%xY�l��6�y��y�ܶ�d�W1�J@vLC�c�����J���V���A-�v��"Ox�����v��JC	�*OL!��U\g��d^����黊����(P$���2<Ɲ���rm�_Xz�Z�z����_OsbG;lư��d�UY,�ZN/a(���x%]�i�b��K����H*��) ,"���Y�K-����[��~�5��f%����v��|�O!�^X�:�106�~Yt�l%<!�,O�>
'
4߅�����S���^x��u�����������9`0��ҞQ$��0H�r��+�(K	�?��������.���v���ء����A�<�K%�����0�N���?�����L�q�M��WW��S��I(q8�����{�	�:m���K������;�p��J����_`�=<�i|_�%�y��]�:>�3{�)w!�0Ȣ�S5Ah���J���3�U�f/|Z��됍2��]�����43#��#a551�	j���o�$����CTbE˪{������h���Y$}2�i�򹩔nK��K��3 ��q�� ړ�6���<�|�E����bW`d�f�pw=D�� �#�"	<rN��#l��*����"�����
e�;:撎�0C"����p�ㇴ�o���f�өap�.9gW��tL)�P�d_vY%
r�D����� ����Q�~VP�u��C;��_0 
�ʎ0�]X������R����4�a_�f�]����� {���G$Q�����r�@E�0�`���
'{�yS�h����4Yl>�ś���Y�ܟg=VՃ�%!�ӆ ���ʯш�5��E��b́����c y����EtI=Bb:|P����XD+���~��B��,�/,	w��Td����is����}��oC=��5����~H=���Qj7��?Ux��X��6\�
L�㲉��)�2�B	�dIg�S��3����Ci$
���i-�3z����@<���3�8aϙ�&��MUp�&&}�cj�1*Uw�-��)��3Lpro6e�5��լx�0��*bgi(|����r�w-������o�bu��S ΀�����U�$�����M'{�}b$Gb9Y-�]=�������h���c�Ths=�B#�Y
� ���Y��t�狟�V�ɾ]�ch��/-����#�Ml��lX�@�J��(��=�kh���&��.^C��.��m��x���]Т���H,Úr�yX@���;�Ƣ@�l	L㥥8_���(_�a���p2e��W�@�x��x ~4�� �+��ٽߍ(L�����H>D��Uvg��c\�!��~��c���h}�!�2��~�ig� �/�(?~���x�� N��v���*��b.��\|7��"S$����-	���h	��0U�ob9���z��������n7��@���Zǁ��Þ�^���̌M���Q_&�t�� p'��.N#���a��kh�mf.v%s��z�P1M���]�-�+#>�R�[b��Y5@���s�����~TG,����W�z$�dmcù,�c�s����tE�o[߾X����Q�8�z��6"p��y��Y���6�Os��я�@���9ޤ;z�~��1���8��ʗC���e�?c��O=�ONG��D��8)��e�1����1�f�R&���,�)Q}�~f�?�ۦ��dG�e�j�y$�)T���>	�6�N��%i��H�$����|lp����@�K��gP������w �Pf�Dy�i����/��c?���=��N"�%�1W����	���z��>�)IO������+�^d�Q�!/���F��G$ė�<|�VZ��޼���Ͼ<��*ج���S�o����҈=@�W��)�:V_������fF��U��,�}W��C4k!)�Љ�S�*�9���k�l
6��	���w��(���U�)��Od1Do��03���$5��u��I�c���0Ǝ�	�|س:�����䄽�+�f�	^�����{7���u��״�?��|�U����e|9e���r7MY�*��fb�&[��l�"9=b�B�	���?���������x� 
�N��Ĭ�g��eH�e�~�!�1��A��0O�,��z
1�8�͞
j�8+ w��S6
ʓ&k���UK:�u��"3�� �=05�	&�b�_���I�U;$�,#�଎%T�j�̌?cqy�m8�����9�J��K��a�1U�m ��C�������Y�$�&��=��ۆ����F����z��a���&+��@f�c�p.���kpڑѦGek(�^��2�ߕ�֬��G���.��'�[tlV��<����l�Q�؝nBHި�E�?�B������U��?J�+���wT�Y�߮B��o�����已j��ӻ��DN�y@S[P̨+�^���g�@�̪��R�u'q��ڥ��M��"�B�L�F������}iC[�Cl&�i�%��H�`���O�[xw� ���H�.[�j�PY$���Yۗ6ћz_� Spz����-�u��KM�$�[�W���c��Wk P�S�r��0�1�:]1����������z�R
wj��0��-�G#z��d�#�Jn{`{tM1��e����c�e�
~L3�!�i9b��xS|eŁ�h���ӄ[���w���Z��*lh�)a�$��;=���Fr�� 1Q�fl�eiW-�V��L���S:Z��@����~�ŋ����Aq9;�O������M�(/Eޑ����+��@���U3w>w6�Nuno��«�}���ŉ�F�E*�[�%�h��4�K���̩�o�jOr�Nׇ�Q�f��l1�'ziQ�׀�>V��C��O�Ϟ�r�]�����DRxi��G���ښ��`e"�����a5j����	�ܙ�V�x���T������r��#`U�+�PaQ;*� s>�0��w��F���#:��#�'�ʥ��Ȼ�BSB���`	*b�sGԀ�O�TA�;���eӟ^�F ~4����<
�G�����_;[&��6R�]��G^)`#S$�R����ņ Y|�CAV㄂�[W�NLÔ��EO�D[-3��0I���\�u�Q3���\�6�`�w�dߊ�[�+�-66yE�B}��核hO݃���Zg���B毉t~>ʣ����y6F�>�iG~MzU�xS�Fw���FCl�Q��-�.X��S,�r�RI�mxu���Q~3�-��c�`4�a>i���<,F3��C��G�8F���pHT�/���3�?�Y	H��sg,%;��B�
�hX�)�d�W��>�3�ث��%)��ј$b5`�2�����b�A�=�^�H�l�{�c��sxNIrgx�B��_�F�x�V�����(�Z�io��;�2<X���Up43�p�x�, zȌ�� ٘j��:�#]إZ/4sѕ<��;*��[�`��j~�B;i��9��o�d�A?�#N�c�0H�wa=:V��"jF�V����=ʃ�[���_j'��|~�-���n>�?:�nb�F�(�^��'�:���w'|u�x="�x	����E��D��z������مbN�	]T�e�����mXɟEUn����Fr��(9��B�4�����C�����I	�	�P~��y1���h��>f1c�/���a���]	v6����|g�PǏ�N��k1`�����`��-v��3����6d1Ms��C��*�<�=���~��m|��g*ɴ˴t��c�` ���F����:g�(��Cؓ�4��\��mA��u9��p8�t�Zm]���ܨ����H�_.�T;�A�D�-R�a4#��@|���[&?��N� ��F�mr)�v���<$�K�o�{�J*Qi���$��mpG�!{ѹ ܩ��+i�n��Ō�(j,��'����"f�\m:3����	�Qy��I�w��o��o�6�/���q]��Ad�M���)U~�M���+HB�)���g�+�'x��r靬����0�\�Bc)xNM�?���Z30�	fSL�I��8�z4��9�N#	�b%����Z�ђ��ax�� ]�N�l�]�2�>a���w(�v�o���}���>Q�� �T�a��$�w����� $Yw����%�#�=��U��WR4�a!yxj_�!�7�H#�P������N
��:����t������k.�$��k��`A�O�8~A���^���b��:0Zې�im��͝:�e����.e*Ŏsi�X����iI��5
�uu)v��~��c���e�x}�	���v ��-F����,4��1��Ѐ�s����$��2�K}j�tsO��+�0��$�'6=ɗHu)S#����ӑar�TJΝ}�&������j��%1��e$8M���(}R��	���?�kd�ɝ��A8��S;���c�;h%��L 5F���>�(��D������.7�,i٧B�j��։Δ�l��k����RX�B�Ʋ6+K��40N�	i���/(�{�57+e�U"XVL�䬥0g$T�X,�CA`#o�hz|
��{������U��Z�p�~�I0�Wo�?��>��J���t*�͜iW<䴻� Q��� 'Oґ��*��j��m7W��x����)d��)��ՠ=� ��z`&�R۩���)�*�*�N�ͯ)m#kMtM�Y����)���8��h�W>��%˖��3��8*E�7���_Xg¸�������ެG�{멒Q*�|X��A��lM��x�kQ�n�	?��K�@("���)	{���G&[���?w���Vz�M�E����|����O�`T6 th2D��NJ�j���Xc�H�$��n��2�e�1@+^sK;YT�{��{������"=<�擸�(��*l��nz,zTK^O,6�(�n�*�Y�o�rK���B�R��%�����$�j�D��L��Э�Xw�vsO��7�@�T0��?9���^M����$mh�~Ω�lf3��0���� �_��m��S����$* S������DU|CFd��s�Ů@&n���,.�7�=�V���{%�1�~_�?4��ۊ��w��C�,A�� .�)m#�_O�@�S�3=�R���]
��~��}��`�����Ah��^�A�bН���TV�=�P���4���!+�ⓓAȢ��`wd�n%�&�����M��i�q׽<=�A��U�SS%����O��ħ�I1@x���܈��d��,8w����p�r��Ţ&{�*�?�R�>��>[!�R]g�}W�N���]�I�*`E��5�
�W�d%���S��S��C�V��pGSv�5�3+�Z�M���ͩD�^��gc6̩a4����-U���0!Ĺ��[���Q~����pw�g�e=��Q�g:�w�s�?����\ ��>�s�uuP	��!�iڗ�P��~z'N��y/Bf�|E�Z�.���D�p�YQ�����>�f�`u����G�D3?�`�ŋ%��C�m���4�`/�.�k�����
�q��8��yW[>�s���|/��tq�}�`�#��t���KS6�,���qv�$$IF�HW��+R�5ß?��]�m/ɟ:���U��hVǈ��zbsfV��*�ܜ�r3�Dm	��a�c����S�����~7������䯨5r$6�w�#���Ɣ09�i@m'{!���BGJH�����=>3A�&��C����h���[8c.���vzN�ǥ�7�u�h
�N^+:���s0�j��Wړ�bs4	 OH���8ѣ�c7~���J�V�iy�+����Fv�0պB]$NJO q��;SsHt�������_'M����Z�/	s�*on���y�O�Q}���g�M�C�8�0:Vx]�%G*Z��:��Rr�:�#�:��4ՠ]n��+���-s%X��!��K��i�V�� ckE|����W�2���y��g��w��3�B��}7˱��]�ԁ�a�4�哇__�o5������Q�l�� �;�?v��+Y&V�b�G.�iKr�^��MP�x9�2�W�[S:!p ƘI��1�K��?�et�[ɽ��3��\9y�q3�み����m���\+�ԭ�"�1!�QA�O�H��ߜ$�x/6L
�d��2��l���h^�3]�'�V�~l��⏆ޠ��e3Jvj�����*�������������� 5Y=�I�D��N�ϖqzf�Ual��[��6��9����:a*ش�	�d��hdh���]:~ErB�o�������9#���ܩ?����'v��P�é�vC���}�m���9��QK�e]���Kq�0�5c�a�a�S�����i��;p�S�{��z��!�]�ga��t�_=�������!�A�Qs��|GS|�+ �`���D��)�x��=*%-I��N��>�C�eR*�)ي��! ͐���?״��!$d˝r��%Q��-�d�i����;[v)�5 ���v`���!�B�w+L��������.6<���6,�)Ys��d� ��pY��,���Z��tn�{:���qO[��
��+�@K;��;?΅׵O�7��vٚ�D�����p���G��J'�b �橽��t�nF���\�ނ�w���S�[��~�WJ���x5�0|��Mǌ��fZ0݃<[���g@��'��?���R�K�������e6vAl�~?����^8�i�(4I�K�Rs����Xp�a��r�]��&�S�y�5,:��7�_��P��Q���������Ӱ�!�Q��Fš��{���������qD�� �܁��uG)�(��װ�~�5��(a��$�4��.� �`$���-�4P>�� �0H�n'7R�c
�e�6'�� c��~��%~m��TgEEsp�.�ع��'>�'�&���J�k�$z��>$Y����$
��vK �n}g�!&���.�m=J����ʴ�,��@9�����d�8��d����>j���E"��Z).#���`�Æ �) j�.���I�8�	9Gɣ�����;��a�Z�T/�@~�jj3��p;��4gz�n1A7B���o_ �����$?�Y��"���ai���D���}_>�u�~� ���H3���5�^����zg�l ��.\�:�����q�����' ���)������V���rF5��ɉ�-�9��o2ET8�)�JO+q��5�UnIMH7�'��WrǷ����6���<�s/G|G�o�-��o��#W��:+���S?��nM�z���G��E����%����m�nz���zf�;�y,aګ N���.�,�Nk���}.Ӻ�w1�6
�4ݓ�o(fS����V���{�
)���F+��k]�3��rt���2� Լ�G��S���٧G��E�fm��g����3�%��]j��۹-n�8�h�C.�#?�p��bb��y��G�-^��JɌs�� �롙�Ꮽ�q����G?�G�-mܳKKгv
�{��M!����#S����j��?H�/�L/KAc|�S� )�x	�.���׿Z��vW����8��m "ݔ��z��U�5��{�ɺ�Ѱȋ�X�7�ce�|Q/um_��US���9�~	'��`|0B� 6��A�Y���}�) J��s)���.��&N�q�s�=���~��c�Rգ��SfA+���;�7���<F�R{2��~�:9�-8%�_A�a��\qȴ�Sc3?��P�e���eW�6�~��LvAg�ʵ�K����,��-�^r�/��U�V���v����~�)1���I��G����n*~a�R�GSIjR�ºz��V �n0�L�Q���5K_Q7`l�5N.N���l��o��MȱQ����HH�G�:�xB��0���{�E� EYg�"h'��=T-�佥��X>�����2$�_��I�?�.ާ.��ԓrw���"*�*n5�ծ>F������\�֧FO4�~X�SE�����̀1��~[��	7�:�nㇾ�"~��Q�H�Q��7�-g�hW�h�Z�_��󍄇E���/��3��>�.�f�P梧�0D"�r���ul����_ڧ{`QΞ���4
�?�j�FfN�x�s�?��P]#�(�8H�ߍ�=V�}���!�[G ��e�D��o��XK���ae�_���qV�23\"´I��H^���˽5�#3��P�5�T%��r��������bM��d���}�b��Z}z��\�>up�}p	�(ѥ�6�v�3O��΁X���4[���f��0J�D���}!yM�s.�t`�hl����Y\/s��mA\=@χ��u�1	�$��(ɺ�Vn�~6�C����x[��ū��ܟ�� F*$��m�2O6�bd�0D���3�DuJ�g��5�"�	"޶��q�~�o������T��bEp�r�ϰL�V	"���Th:-�2{U~M�~$7+Z0��F����Z�7��S����Y�d|�8>߅�<����}9`��S@�%37��t�|�I�|�mF��I���8 K$����!iДc�&�Go�U+�ext��Ɛ��r�&l�t`���t�tF�88L5��۱,��O�T8ų���*b�uC����8w`���B��,*W���_��Bf�Ak�j�X��>v�4�m���4,q���Z��Ȝy�q�c��5��l�����n�X ڳ���^fu��Y���g(w�/�m���F#�R��m5��2GW����rRHǇám�~�Y��y0}|����k��465�s�t2���Ў��Y������?e
�mDem|}0��elN���90�B/��0xg�hڋӄ�-3�wH8�8F;L�g�J�Y来��i�2]Q�a6/�����Ű�_Ƙ�ӣ9G;x�f���$j��݅�:՚�1i�����
_���~[>�����T���1�g4�"K%-ƽ���)�6@�0��O�ǴZ����`���97��c�[!��G�RM�	�R�2Ԓ@gzf�����ڴ�T�qY�Γ8y�^L»�nMR�m���פ�:h��YF<�/� Ƚ/��|I���+��_�ւ����5�TD�7�	�7ZVo��e��a���lʹE 4J�!fo#@='��=��[��!��D)�ܹ�tYx�K��]��Y�*��8�=�33c��P��%hQX\J�YV�ΊK d(��i���	����N��܊kH���J�.^������U�3�R�;���.)�y9��U?�00HnI�'/�{͠� �E���i��%h:�R����'�Ґ�-0�^9i����~�����줌��akj3�"��,ZO�WT�����J��DM����n�9��-oC��N_`�U� ŉв�S�?x>8�cy��W緦�ȳ%�?�P�tY��F�5���&�TI�U	�p���,�n7u|����Vһ�GQ�	�+�K�c�5��_��w�a�s�E��1��FٚD��W���f&�w4�nv���s��-V���|�Dso�=ꎐC����7�H����+/�/lgG�֢��X��M-Lkț28�Zj��/!�W�8��
��g�۫��$����N} f�,��H/�aT�:+~���;93�d;a���N�Ly4fl��R����b�i]�)�yw�P����g�hT�$�2OGr@�ˢqB/#�Q��a�Fi1���-T�����eU=�z �g<�_�}o]KD�݃��l��Ja�O]ڐ�m5���z��y ��N]ܗ�{
hi9|*!���+x�Y?܃7u�����!�Ϫ�����@6�7�x   )��U�(�m!��wG�$;�c��e"����-���ߗ��1ym]��J����ٓ1i�>����V�a�%[��mQ7��<��W��	�ܵ�f���oĜ�v�!���4_`�{��v�;�*�A�	O�=0n�����Gۃ\��^r��sABFQ���lr��H0��K<7����r�;(���Sy�x��"n#�g���z�,D����m-�v*�Eb��iv��5	���a道��:�����.��=�3R��+��ԖS�nє�~�􀑫��U�B��}&A7��eT{�W�M"�}�����KǙ�����S�����c"c�2��E��q��J�y��S�7��Vz|)X��`I�}��-���aC#�}�.V��\����u��'@�!���5��.�����'kk s�~��<{b�aYJ:�1l���Rl�������_V��:Ǉ�#f��c�h���F��Q��F�&
��{lZR��_��綗�s?o�MYmG��
a�}�����*{t.t�����H/�&2W���er�pbhO�:hmr/�k�W�"��J�״O2^���T���U q\�&�^�]ф�z	�yCB?�sb��Ȟ�K{b���C_�_;���w���^���v"[F�:�寤ť�,��$��{>����#��yF<#z7�f�v�����������C�I��Ξ��jQͥ�X��|!!��{\���C�]#�O
^1Pw�}��܁�7�C��p* ��g!�+�&;Q� Y���-�{C����v? +�I�����J�߇�	1�b_����9ʧ������Y��ݔ���?�t��pp�K�W������>�r��'Α�VCg/��syH��렗�`F�r�4��RK��iq�YՌ�ơ,}�@X,�i�y��/AS�:��l���D�'[�e�k��i�����������/�|�����;G&��a�s>�	���α%)Y;��lM����ȵMT�}ε���� ����sz��~�x���6��=D���!�`�0.�i~M�
��ך�Ǯ�p���ķ����9J_��/c-G���g����hG*MN�jb�>��*(`�gaN�o\nX4F_�@��(����g�W9õ\���7��0q.��mTXf�Y�G��j4�%h7�i`�yA6.(�G
R�b.��ܥ�d��q��_8�#!��;�V�Is\�F`OU��|���}3�5�����(�R���0v�v�=4<��Q�I�E�l+�-�:z����*��4�_���&RFq�i5� ��?VU�.0G+�eB�=�x.��L?.P�l��W֪Y�\�T�:��^N��i &*6�g �R����2�Z�㹺�1㹱_a�����]�N@��C^4�`֢RՊs�"IX����<j�Q��t|sB��d���N�4]F��wX5b	=W�ƌ�%ƶ���}�U;�����5ڐ�ˠ�$������O"(G���= n7�VR��n`�u�74ĕ����y��1 E���X�E� b�h���)��)�DWϻ-A{�x���*�./�6!ٚ`9��f����@��קm�"���aR2r�������n]s�����A��)X0ʕ_�A�׺��=Ѫ'81�䔅���GDJ1[�2�s,r��L�,C�F��J��H���M1�'�;\���ʃ��G��`����\����S;�n��S�j��1>|?����h��>�o�;<�j��3m�JA G�T�n���2T-p�m��S����c�<��E-��ⲕ��~��3)I�4���l����z��x	7�{N�-!��Fi�^C�r9�,���!����u��N���;�<��:���q�q��-��9!$WU5�8?%����S��Mس��3A0��Fĩ�By �Nj�*/�����G��w��5F�-���%�fK��K>���cD_��%��G����(�e��>�ATi��讹�NOB���FЂ�������NQ�7���Od�Y>��Ԥ;hX�W�ՠ�C}��z�<����Tha r�H&sD^��<����Ā<�����@��D����̿���#�WૌW�?�I~�zD���@��HܘU'S��9�;�"�cT}�����Y�#s�������c7�@:Z�O|���C*"���\��;~o�!lt��:$�/C�Y]���z�V[����h��w4���CkJ�8������MT����\o�k:!�ഫE䟅�����d�)<��oȰ����1+�%��q��%y�؁U�0�Mu�E?�1��Ѷ�H~r���<l�	h�-�?=P&����Z�r7�,V��V���FEd�o(-P[���Fw��kb/D�Z$�Pߟ�Y>J1��{��d�ڥ��bn�����JmG�h"5��Q	���`�oI�L,W��zzS:�X�\�Ռ�4��k�b5P����8��_{8d���i�sTo��Dڭ�|����kq)����e�^��i���d.d��폫�>`J-�U�f��q`�f���2*�d� !.n
��u�%i�y��5����\{�� ���@ݻ3(�$u�Ͼ��%˧�Gv��$��qr�Y�[��3s��.]��Pز���ٶw�ڳ�����)��H�\�|���ʀqp
�D���e~��t-�qi��CC��c>M51�ؼ�.��SZ͖2mǅ��S�v���r� ,��� �Z�D7ޟ�]�_H�?��Sb��/_�ޏ���(2�bX����l2DK5)�nE!�n���&��7H<��27�й˨G,��Ԫ^mE7 .�Ou̞5���l]u�`�T�:�B*���H-Ԝ�K�A(�ŝP\�:@����J��f�q�"�aκ�#ա�$XŴd�wzKf��=�P�C��u��_eH�����x�/���T
�Щ��l[,���I{���qP��I�%����*��_���އP�2`�xBk�^p����z1W�Eۿƚ&�WY�p��C56��r�C���!��0"O�daޭ�*�Q�ᡸ#���Ŭ׍mؽ>�VE~7J��@�"�y����C�D=`r+����D։/0U����TQj���"謀���J�o3��e� Wy�t�tTT�͹��X�+_O^t�M�Τ��*u2����	�.4G���xP�X�B�q�;)� ����O��ݾ�;
��B�p�v�{	���|�M?+�C-+��I
ƎQڞ����"g\Gn:��f�*��g�d��)?�j�x�n.BAy��*L��Z!ܔ5W��w`�E�;�|�g�z��<�:�AL<c�#u��)W1��Ǜ=�=��ES�������z^�e>�0V�t�a���I�d�����^Yޘn�w�;m�"�o��hQg�����F!����S�Cˑy��?�Z��x�l�@�9π�O��E_�eܵ �m3�ޘA��E�Gg?�~�u���9r�[m�=K�ä����*�+V�#n��0����m��zH܁�qj���U�"�Ԕ�]z"�32�F�Z�Ϗ�ߎ�ۗX�M����h&s��M?�*%� �:9zɰd'{d�����N2�\�2�NF�F`S���@�%��U���y΢��=?N3��IVlN|��-5O�>&U�D���Rcs�!�6�)��Ϫhb!�|6�Ŭ�lqRA�c����^]������'0|H=��jA�Ċ��5��j���);����lF.?��� c��{S�41��.]�qt-�&8�\�/C��n���q�J���Dޗ�Ba�q���7�"�n�Q���F_�o?�h$��]o�>�����6�e'�r��ľNί[6��q8�_߮tIE�l*�AZvg��ґcq��+-.��9����^��l잟&�+��{=��H_t4q������x��J��-`'�2�0kb&l,�".�����H�չ��IrR�7�yM m$��/�ֱ%��bT�!�2d���h
j���-B(��b�E�[Ӑ*i�����4��"�S�X$Q��p.��=!�R�3'����&���b �Y���Q��R���^}�4��?
� yu���t z�сLPz[��o*zͽTty��Ïֻ>!���@[8}:s_f<XO<�ֈ*��"��'�m�5�S(W���l��#G�e��t�!�����A����4�� J�L��գ�R5�}F�+Գ���$&���Q�7u[0O����"Ol�I���r��Tsj-сA(�ϥ��ӻ��O�H�D��/1G�D��;֖S��B ���������Ȥ:��[1G�x�s��=�O[/b�R���p1-�ӗ�kc�VA��:^n]|f{�@ؤ	��o�����7Z0���\�l"� �G +�8l�Xы�^�4=tM�
�r<ΠJf�Z�Yq ���۪���4+poO�f-�U���V���ډ7S՟��b�2��;)���S���Ik9����Sh��|��-���l�*+b�7N �p�ڒ�{5���6��l G����/#�)&;f|ڦh/���}o��u��؛��d��B3@$7`���Q��4<2LS�P��v�5�&\�#��|�P���1\��Ņrh��b�gǛw�Y�>��)W��%��y&�|$�ӯ{/*O#:�t�"�8e��fy��t~��cH��� ��3�O~���簜A ��g�����$b�K��P$�~�Cf3m�Kd��t�W�5.l�!r��(�?��&�3�#V�|y�&���N� ��" Μ�c�'$uvu=��0��`��G�/�Q�7�d�-�G:�3Y}��	�E�j��{���������8�ݽ�]���>
H7���0�Ŵ�$�k�u��S4.�7�hˠY�Ȯ���O��]2��S�j�j#�hke����{�%%���,��T�ˍm^?�,�n�T�Y��m]3���R������Ue�Xa�&���c�)����)�d�TD�9,e�h�̗	�Rq�bY�â���B[����lU�X�}��h�R��;L�(W]�ϊ;���x�\6�:��ϡY]B�X��T>�����^���k
^>�4��u_7d_Q�J}�o�#��o'{�>��rTj:��К9��~|�1z��2�����|s�[v�^V%���L�^͊�%9�#��v܁,���~y~�H���+���)V5�y�XcJ����.L���ʎ�l^��	R.�<5�$�/���Ƴg���(qw{xKH�������-3-����� G_�{� qs@I��S)W5Zso��(~�������j��Y�}� ���A]gJp�{�m���R˜��بp��F�����g�p��`�y�E��ىQ��ӑQ��b�-f�����>����H�%w/����&���b|:��G�dk��!��\�A;UP��9�U�{�!䆣"٬l��H��Z����ޤ<L��?@W
4�P�آ��}���
hv:�BO}|�(C�#b�d�(vq�%��PN]�fQ�>?Ň�4%�Z��!��䜿���GC�� ^�]t����B��Qµ�#�ʰ+�օ�����'TJsw����1�Fx�A���ħy��z����Y��+?X�$�&�F�ժ�*�bW���b���/�K�躍[p��9d��k�m#�6n�,���(ɖ��@��Y�46|���ء�Gug1���u:X�Y��u��A��N��=��n�u¬e���B�gn�>���ZZTP�:�!}.���  ��d21~vVA�,J�Œ�>#��\]+��N%�ރ���K[�"եJ��1.��,�ok������o�h"=?� ,e��u��جVr��W�Ŵ ngԍ?I
�|��
v @qUY��1=������K����_��O�D�E�,�[*{�0�l\�e��9 -t��5F����;xgl���-��72�R�5�˵$5� 0} ~��T-F&�-��s
���#�� � ��:B�5C���W��J�Lu��]k_�
�#h!�?�����Mbqjf����3��/���u�����̲nI�k
����͛y���_������w�u���C@�ΔD��j�lJO?
؎���>��X�?rgp��g�:��J1���ǘ��]O�����'�$���\FP�Ey
x��	W*�g�`O	7����U�ͷC3خ8�!�
F��^�S�ַ��� sl�m5-%L��Ͻ���cdơ/�9qXa��$RO��lE6Py���N��	c�E*��1W�U��n˽�B.��o�SD���w����v�~`&!�	8��0��_[�􄔞�P�:��V��_W�G�8B���9Í'3D$d�[���hl�h#�Xg�p( A�{�9M2�k8���f���w�n�J<� d����;y����rC�%ñv�&!�N�d��>�r��:�b�`-+��R�)�˕�g�'	{%���i�4CRT����&���ӱ@�%�c4X��)u��K�F��ru����foh�|�a��?Ko<���3|z_�1<e��i	A΂FU�n�z	��I���򒾦D��V�d�����50�vn�f�T�f�Y���{MK��a{���r��)�U*=qxwv��L���w�"�04?�����\���(KJDm
�=Qn���Y���)��8�03�a
�= ���73���I+
.y_�O�?M�A�Z�Ʒu�E{ϲ���8P1]�4ݺ�JSKG_l���<݀�G:�S�}��!���|F^��6e`g5E��$@�����q�&_�s_��:��#�֑A&J��\wH�'r��G�6�@�p'��W?�^�Ë������D���I��f�+���	��=*B���<��=�
E�0j���i-��ܧ��i`���ȐI�&�L_!�5h�Q�x�A#�V�,2���	�8u�b	v��(����P���i�;��_"d�������pZ��Ҧ�'@��{XT*��T�A�-Jֽ�V��i .��W&�7���~p����Vi�ʢ���e����P�B��B~c�|��ayhW\j�zcF�x�7=���	�Û�Gx�u�`������f��C��F�g�q��s���DE�6�t�&\��d�8�?Nh�&[y���=9��j,�,�>��A�*��B��L�oR%���Z�,��Z�Ƒ�������K��0>����Ɵ#u��R�d�.�̾Š|Mz��u�8q�� �Jh( n��]��Q�'a2�Q�yІX�Q�x�:����<�6,��
R����+���:Oۉ��BN�\RaR�9�BJ��T�n����0�*4�Ql^I"EO�g��z)�H2Qk�}xt�2���2�mvo����4	���n�Γ*� "zֶ� ���j��Ƭ�@�b!�̥Q��<lZ�F�UI�Ʒ�]��``�Ύ�)�����8?a@�IN��R>�(*0g��&�^��bqHGX��%^�7��?��
{�a�"�
�#�Տ�>�����!(��O�~ �Mt^�E�=�$�dx���}�/�ʚ���=�k{�䎦�r�=�����U�#$ԙSR�e���H �: m�Y�8I�>�Hl� ڱ-v`1т��I&��i�uDS�0���;hׯ��������Q�����-g���`���)��,�4q��_��t�>�G-� �����U]hWCyM���@%2Y[�+>�s�Ϻ�����O�'�<޲�l�M�����:2�I�-iV��Y�z� tEU�3���T�.^�
��K9��\�d��ӕ�d�eg�(��'��FFF��9�.�F�����K���F�������(�ٜj�3A���< r.���;v���\��?�_p#���s��$�-O�WIpY����P�9�>���0͏�Ʀ�'u����;��u��;�����ȑ�s�}oQb �ߛ���T�,Q[���?;\��0�R��'���˪k�bX�T{���]�����is4E�������$EeH��Ւ*�Y��fK�M4�	�=�g�����}�hy���C±�MN0)u?t�`�tqG�����h�̱��1��� _�Zi�̩���EU�͆a���f:�Ǫ���}���*�~S`sG�F-<	9l��&�n�Y�Bl1�y)>��q�����bܪ.��`��
�y����t��ܞ��js���k�w���>FL��Y{~Pj~�J��>ţF�5E$yS���~�s�b SO����{FK�%4Z�`��;�'�����F+hw�?Ԃ�Sy��jHnj`ل���*���@:�ON7��d"�9n��q��A|�U�hc���i�{��J����tA��2"�O�)�ϒ��-3o��.�k�4#S�I���p�
I�}��oe�C�
���Sm�'Fm��g��	u�	��Ŕ/"R]nQ���L����g� ��^6���Q�ʃ���L�eް�:Ut#��Q�2^[Yb��b'�Wk�6�䟯� G�zsA��r�ap���7azX#��iz1?�;�A04r�]ތ8RDI#-�\js,L�e(�F�Ԁ︤�$S���]K�nW��H��?�hɑc%�F�����/2�{��8�~�¬�	v��㴹v��G���	i�Ǜ���=��ˬ��߭:�:A���,���}�2���D�I���.gWl��i��T�i5k���@Sѓ��-&�0
2Ύ�g��S(�8����p���Wj���lhț�`�8��9��"�7m*gN���x'����/��?�7S��0�j+
c��PCw�ߙ��.Έ{OeM0�t�>m��gPk`f�I�  0i��kJD)��Ek���=~K_S��%_l�^��b�L|}�Qr[
[�F����6�&�!'X�Ԩ}�_���ՠ��d[e�*՟b���:�:(<�����+zl�[�؟+�h�",yp�U�Q�
�^s!~/a�Κ�.*�a"mR�C�%�H�^n����w���$a$tH�u�$�i��9-8�s��8���N���M��)�!R�ч@�j������'�`J��b6v����W;U}��;��cJ�,��b�L���/�E���,8��5:�=l�g��M�T�Rm��&�t��9+�B9訇j��Z�%N ��~Uϭ����N^�a�*E����4G;!7)^B?�F1`B2Z�EX�U�8�o&�(��f��u��S-U�r���r,����iHӎ�u�y7��")�E��y�����
�:�hc�s�3=Z�y�6�9�	D1a?��3���&���λ�I�"p!`�MXr��>��� �!�V$��,_�2)ȝa`��ұ�n�����ߌ���i����?�����O�A|Q2��-]��1�eW��!���'�����.����߂.�	b�O�%\˛ F��b����rb�&H�����7k�$�	���޾��0.��}������+;�%s���|�1��?UB�]GG��s���]*D ��s�,3)���� ���\=�ng �RMΓ���aJm��e΀��h2�X��+.�k#�w���ƭti�R�zb�q�G˯ߍ�
��?(�e����-~�[/Ȁ7�r�R�4jTp��/Z�����6��(ȀY}�u�L2�E+�R+K���q�G����o�O4cGe#)���,�����J�K�J�Ȉ����7x���mO#�D7Mi�!�ʤ+�"FaGޥ�q^�]�%�z�Ge�p��l��[�ؖ�F�b|�up� Tv8�n'�ɑO����rn�+S��W��$�C�D���V�}!^�g0��씧��Tlo_"ovn��������E�A��"�]E�S�E`�L�uJQ �x}��UcF�7,��^kږ��V
ۚ�a��+���ׯ��x̌�=�qDB�#��6���N��H2�w?=�U�t��ټQaɔB8�v��9�x���%� �4/�S;��l�f�7fl��O����=��o�ch36h�<��}ꌓd��?���L���..����@�_� ��~_���B�r�x _��u$�������:��!�q�/P �~���|ɳ'����M��C{
�Ǥ"0Dmzs|_F�Z^�m~c`�kE<�m+��l�WHH}]3��['�J��(���[Ӵ��^���v,�<��"��͆�U����p�u�1�y���ն?�`�S�%#Z�`-hD��Y����$��kXD�tba����@���u���pW���h�I"̔̆u���]HX3����ʰN[Z�3�gI��Յ��&U!�'�W6�m;w 7�ڴ�i�� ��h�a�V��Bֻb�D�)�����7�@���l&d��P�2R�CՁ^K${ �3�'8Q��^�ע1 ��G��
���JmyQ�O_,��x��p^M�:�<�<�����d��Z;��L}�L�{WW���G`�2� �^���r�q�����@��
�&
[}A+��U[��8	�}���~;K�vy	�v�8�&��=k__�౏ׄJ�Hyҫ�ؾ���b��,��>����!2���qP�{,	a�|��[s	A��T&pȔo�ң4w����u�Q4R
�}w	�,�uA	EҵW݅�H	���e�f/��5�X�N6M"4�eF떹�ۆW�Aܩ�î�r-=r�H4�/9,NN65?�+x���L��!:�c�x��,E���O,��:h�;_&�'��W��e����Ǣg#c�g��<k7��IB}Y�qj���P�V�D�3
5��`iz�v3�����
z��4��Ó�u� j �c����u`A�4�[C�`|�9<N3;2����߁�����ar�����X�Kes#ne2������D'~y�L���,"P]+�Ɓ��Y�|	Y	��FX|wcv���N吻�����f_��'m���EN+�q��{:�d��}�W��4�j���& h�J���&/�WU�Y�wh5
�X�Ku����bRgs-A��hs��%��U%Z�[���f�����9�a#	:�f�>_�,���N^������skd;'���J
b�q졪�n�u��L���z��v#�=����4t�:��]I	�[:�=���2�����:������!뢥�lK�P&!orz�VTh������Z������<]��RM��#Bv�T˛DszG�}<�	�D"G�b�Ж�p�����gJyn}��m�6:��b�t&#4�$�#4��g�r����ZK�w!D㛱 �C<�6`#�"U*?�Z�c���z1�]�3XE+�=�R��kg����X�76�ITֵU��֢�tl)�f�,���G�����R�n%^������G3�u�E�:�o߹M3M(���F�r������I��y\t�Ņ8U%|���Q��x��1�m��D���М��9,T��S�6�q�O#��W
 �<��e����*x���	�t{�`��j��7�ӥ�E���
Ȃ��k ��#,m���!�h=u��D@x��.���͛u�'��6�`��N* ��_�?�+=� �I�\�%�<c<��de�z�mR�fŏl�e� =�=�ݦ�M�pON��G���V_�+��*&�6 �o9jңW��U߼+:�*��/q�g���=8�%Dg&��(.�ç�[��7�i��/ԓ9g|�����'�a4��F�"��7uXB_���!�f��~�M�x˨X�}u�.-�k��VwG�ޢ�䂒�{�5l(3�/}Vuk�VZ6��e�[w1��af6�u�f;~�&�'+�݊;�F��c�u�U�V�0�(� A�j�lۻ �YȚ%�T)(C��׵�V&�A��4�#�v^�Y��-�����S�x�թ�[��5���G~Y�E V�ϯ$<�7�НB
{��ϼ�]~�er��{��&��R~����2����^o��=�ݓ6���{�}x�0=�&����x������>���d	`1IIS1_��07�h3���+�q[L��P�rnAx�"�JӔ�k��v��Q��E��9b�b�����$6X�"�Z2N ����4����:��Lh�=C2O�o}�����Q2m�+�+��#Z�T�ݬO�ɷ4�^ģYA��;��r�W���9 pm��N1��ǻoGg{N�tZ�/^/��zc��1��q�<(n� `�#F�k||��a���<�|�pv���NH�r5�;������tZD�3!�yu~>�!	N��-_�����vY�ߓlɃ��[���b䥓V=#�,�|�$a�+�+�2"�7�)Vف4Dc�@��hb._`ۼ���n^�x�>Z�(y��g����g��EB��$'*g�8�yβA�p{�����w��"��%��11,�l/ ��	�(6��+^�ֱ��9q����2o;�k������RH�o��J�5�o����AO&��u|}>8n1�lf`���|�p?8w	
�<��z_}�?�A�F����5X�����S����
�F~*�ա���G�!ȀDqa&V�؟��%qR˗��%@bD�U\��C$q�A���>�zrm�Q���Z?j�a�����|�Q��td`��V��O ���w.d7�N���e5a��y�Чo���D�L�x�w�&�$RKw�$5ݴ>���Q"��Uʕ)@�߮R��=+��=�<�4i� ^Csk�K��Qk̶�B5Up�l<�~
��^�>)"3��Hh@���D���A��U��b�W�����;�B8.Mk�J�Q��`D	5�33�&ϤҶ_c�h�ڧ�����rS�</7�N�1U��TD%�r��	.���]�6ő�t���@�*�wԄV�ȑE�����#˵d�z}�:�e*t�7� uD��mHZOBܾ�}���Pנ��u+_���*q�H�	B�K����K4j���Y;�ߺ���4k���kZ<^�����uy��p0MgZ�̗�����F+:&B O�q
u�E�� +�5��>YƖzS�{��KR��a�&�^|a��}�In��R��c10�[Eq�>�^^�\V oc�wu�Y��U��,9�G+�ZKZ+.a��f�$�ɸ6��]fb�q>s�t��/�=WT�9���õ���M��Dp�	�I���sIJ3�;����G��:�r*ǚ�hiNf�ՉZ{��Ή��ɨ!)�]$�(��/�K|0����N�aOnW-ᩡ��_���V� mi/�Ý� �R �ro���D��w�:H���n��~�S)jXX.�ۛY�Bh��yk�ɘܧ����Z'��� �-�o��S�	�;�J�;E�%CZ��B��eo�y�"�|�k��ul��j�v����we�EL��~2߈����'z���fu�1�p�i@�b5��Q*�[�b0,�2Ra�3ޤ����`���W�{�c|��S��َ���?5�7<��z98��GpD�2����1Qp�3��6�����������=���n6\ب.شa{5���O��qg7�8��t�&[�쎄J*��^�7�%�v��ł���Җ7j�҄��^�5KF�I;����0��R��*��td.%�������J�^@�|�xǴ���7#;V��UFt9Z�֖hy� s��?�g�C�S,���6)�4��kݒK�vGY�Ke�`9T@�q�Og����|S��}	�?\ށ�lj�����~�_r#�Q=i�n���.�A~Z7i����k�yN�d<�g�c�\?Gg/�C��� ����B�Ǌܘcם.���#�Ƣ�l�ɣ�ߪ�:'@�4z5�����b�X_�!MTo�Mv��!UV��K�(����E��BRE��o E2_Ofa6(�?�.��|X��J8߇7e�r����S��:l�g�Ip�t[K��s��,?� ����]�i��5��%�ZᐝGu�����+���U��?j>p��ѣ�O4�U��ѝ�˝#|E�e�VLf��g��	�9T���K��{~|m���A�����tp��R��{�"����C�qwYC��`�ș��۝0M�0'��(E��w�~�:♲)7bX�s��F:%�$�|rYӞs����c ���;�`
]	 ��
�$y�.@�!ьJ@��#���Ȑ���Y0�(���k����p2�Ve�+�B�fF�3��h{\w��k�%��-h�ޫjM%���(w\4�&�ϊ٫f>@	��y�w3q�ݼ6��؀����ZK|R��,F�ם��_��u���C�S�f�W7�f2��Uo �N����#-#� �	=H��L�k���'`I�B�]#�
W����>��W�"�����ytf��M����R�:�*���@�������C�����m�8@Z�{�/�#Cݩ �ӽ�����d�O���W&��g���/���ڥ�C��a�Wk��� �Dh�}z�>��0m�z��@�Pc��]��g'd��_F���-)۩�[h��-�oǃ�����G�
q�L���x�k�lT�m�
*��^�G����g�_�V��C��YE_�����r���#��S�LL�Q�A�Eό�N���������/���=a�b*�y��[D(͞��l��1����o��R�������ZU����Xb���x�2_���d2i'$��**Iw�T�����>+����Z,���x�Q��>h�b�}rS�v�>�����N�d���Ҥ�W�Lw;����$���
�d�kX�$��pgFe��"=�0]����}�֟��S��ՑGg�I0Ηe��E��
k��������F�)������Qg?/�����{<n�M��t|��B!Ng2�cڶ��"��J:���Ș�+������|g� v��z�LX���80�ZqE������{ӘCz��Ƣ}�p�i嵞x޼�K�bJ�@g}8_4_�N�}z��:cL�}�J���_��sKy�P��e��#�E�A<_-�Q�eL/:Tc�6m��uӗ��.+rgg�7:����P���'�R�����:���7`��t�����;��$C=�T�-��� ~��ʁS�@d��i��"e$&�Z���|M_�����i)#��d,�?MF�h��}�b��ū�K6��qќ/���=�ѵb	��r~�SuHE>/��Wl��7e�|g�k�2�A��
���~U��Ob!��,D	�<!{tL,�9-�|�,&�.=X]��Q�`�\�-�i��"�9d�OTWh2��)��KX@��S�^gЕ�^��������f�f����g<�cwW�F�K"��u��\-�fǟί���ub���4׳9(�����7 ̠i�ؓb��	if�	�օ�N��[��yE��=�H�,{8��ː�1�[�0/��)}[����Iv�,�;�<���}�z߃�ӛT6��Y���>>s?�آ��A����>�C�3�E'�RH�a�����7�b9�C�Qhj�,6Ƶdj�%=Y�Tm�1�'D���񪷗l���=�����6�FPb��ۆ�$p�n�drf�2�I�^��y���O}'A�}�,�|zfEcG� g��w�w�p�V��uk�$��,Y�#�����[������]�6���%F\�A�d-��Y�Z��l�pc����ҳS��"�ɘ�ɦ%�Q�������>��za>Pp��i|�z�\�)^�d�IG� :�,��h�},�!�j�*Pk��ɠK�ۂ7lb���?(k+�NF � ��~���&G�[X�!��4�"�5�<��A�%*v���r�%YS�7�ٔ���Y(���*R�]��8�_��(�R�����4|\���0�'�)ۣ���f^����ik��.F�'ˬ�Տ�
P����.��eS��lp�ے��T��R ���3pO��l*˨�oޒ�#�Vc���?T|v>g�I� k�	ڤ5~nC�'�r Lax����jD�p��c�	�$`�������l$uw3��t�N�\&m����8S��v{�6�C���9���4����{��L��L�T�
�.�#�fw9j�	H�7Qۆ�i ��d���2�Qm��J��q
�P��,����,��w��	<LI�B�$k	M�/�j.�o���m �e�vݼ�* �J*ri7R���G~�0���ϋx�u�{�s
i#��bɇL#Ɖz�l�(J1��*��y�A�t6��UZ�.u6Ṋ�@ ������'J)���c5�U���xT�V���h���S��>c�b��s�B�w����Ш8�ͧF�1���,M�2�p|�E��*81�Hc�^��L�*�
��h�C��Z���w���Vt�0ޚG	@5ǐ�̀��1�6�d�z���n�Q/{�5�*b�W��p�Q)�O�;��D�C�[�[�MH�����ϝ+��֐XJs��L�.۔+<�	Ɂ�y}�u�K9�8�jb
�Z��ً�'W�X߀�]μmP��a�\�ף}�7>��sc;���q9{�:���g��y�"a�����x�gI6�W}0��P�^��*ʂ,�J0j?M'O)'��Mqmeud�^p���x�LX̹���`�	Z�n8��#=�3VEȭ�J<�;���
��;��0��݇H�:Y�5٤?Ĭ��}Wj��)�^u'޴₫2��,2���X����	7A�"ޮ0Z��<���"��vV�'[mK��N����f�K>����~g���re�O�����P4O��q_7CsC\_��

XVgۧG�ʌ*�D��+�.r@,��GK��$���>t0C��|`&�p�aͩ���@��]k�,p���~)]i\p$�s��c�{�H�&�� �T`�l��$�+C���'�ir�3iC���Ϙ۩��P $�.O�~������U�V��t~�����*4=W�^��<����83\=�cc��_��Z���_#V$|%�}�̖��|G���C��D��zRt�Ì#sHUă����CXF�牦O��F6b����T�(D+��xX;�x=���g����/ٮU[��ݨ�$Wo�<�X�a�s<ǘ������]>G��s˕�g0�y0ou&��|�����A�`��˻Fen	B6�0�|,긚
�Fa�%I���7��B��U��+Me�zH�d�N�휰!���Sε87T�o�ԙ�����U�lW*�������-b�N��
0 )�5v�]� (���VK����N���I�&��j,d��=��{��v�t!򽃕�Y�YHN��|$�U�'��e-������DM�ka��Zh?n\vK�^���/�4�N�.'�?d ;X��JoCi�2�3=E��L��wkn��-��W����{�}�_7��� uh�
$�������x�A����t��sZ�n�w
%�Kp�J/�T�藴:���fQJt��JVcj ��t�y��%��^H>c�7R��ܜ8��?����:�G2�F-lk�����L�����kW�� Z��H�?Ͷ�Y>`Xu��R��w]璗��2�ж�h1|������T�g��7��[��j� ;��fr凯�`:���8�aI���ON�f��o��Gy�����~�3!(Bg1�:��_O��5�ͮ;�*�9��26��>����}!�����F;{�Q�LЊ+��˔��Rs��o��=J��-��2�������|��([�g��F}`�o�cR���
p�'��|WIoE��`ds,��u3�0�0i1z��۾��WC�/�����q�y�H�s��3�r���
���F|�A���`1���sk�	{cE�~��h�B�.�5�b��$&a�iM��Fu{�( ^���D�@��=7�*u`�(kx禬�~�,m��cߠ���r�7\,x�u��aO������x��7G�$N�_�>~�����Ϭ?c̎[i��8m�7�B��궬-����D����\@7��ơ�]�^@m3S�ae�Y�؞�屐�S�(����L��|2m �Cͦ_���ʺЦ��:馭��e��EH�k�Լl�����U��}��Qq60���W�_�- Sն��Wy_F/���.d3FŦx����#j[�8O��["��)�!��M-M��5���:��p|Eo�Ө�<����RA����G(W�yw7�K,W9fxh�"�z	oG=l��JOh#ȞO{�)I�G~x�����4d6rf�&���;�6F�=6�2]!r"�<�"�k�.�p��'�F�w������=��"N��5�#�!�3ύ)�(� j��^4���Ǝ��|��q
���'�,�����!�A�P*G��S�b�zgV���S���U榨]X����#�������E�⋈h}�g�M��[����U��#a�5A^��Ud�s峍��~� ��?��B���rx�������ˇ<��
Z�uwgWq��:�+�$�9�V�ZɷRk\3�6��"�[qwaT�v�#�鑒�������2���S�ح�uN�VnsP8!;����*��i���jz�C��Ӛ���@az!���lͭ�E󱆢 A���Y{,�7�Pk���B��{@E�86b���x� ��a��D�$[�=�7���@K%���$6����5���R�g���?h�������z\�WE���1��Ȍ?����,a$²׉�<f��]�~qX��dy�\ۨ�s|pY�z��Ob�h�S��P+���-T����{� ��4o�����2:�9i?p�t�"9��O�j���ٍ��R��˟�.]"�(��n�S)��Z�nC��zn�I���x�Et��&	4q�Wð�hP���9C5*J>�oF~q���N�.�wo�0j�l�L,D�:3�򡏷�w) ���@��Y�}%��F�_�5ޯӥx��v>`j�U}����Ы���.�f����6�������d^�A������&%��J#b��e��NC���J��Du<�@�z��X��t.p�@�c��E���u�`����^�K2z\DA��Gw�jj�:��쓧��eu�0(/�����*��M㿖活���� ��*k����N�{訛+�H:W�E�vE��� @j�{�n�j3[SĒ���DB}p� �����|�=�����c���.Ϻٷ��19,�5�=XIJt��]��G�Ct�Ά��Kyh�^o
�_�
��G������wB��
�oa�<)���ߗ��:q\:�jdx�&zu~���x�莰�g8��/� k�Z��(Ȥ]�Yѭ�@E�`X_c��!�2�'me��B@}G�P�q�6E?d��P�0��^j��G�5å�j��l�kYC.I���67r�|���u�UG�ԷN�0�>�*���m��U�Qu��R0�_�=됢�^$�� �8��W[J��s"��5����Y$�` ��f��U'��"�0N@��Ց,�wS:ې�T�q*��-�и4H�_���v0���H��e}�f���{�f�*��V�
ol���Gu1I���1VHdE4U���_�^��/�%��91!�ЫXu��/��hj�V<�j�_�}�U<ɞ ���O����տ�|\8�p:#��Փ;�A�q³O@������n��+R
?���4𵦮�����3J�i4<-���>8~c2�D�1@�Ȃ-�-K�G�$��������;rC����#�&�р?��jIuc��,5%0����DB�3��!av���;���>�C��{�+�ԟ02d�"vX>s�I.�o�-*��e}�T0��e�_\����e�X�~ڃ#a���|�x@|�.�=�i�q`<IC<	ɹc����Iu���oՁ���ᮝ��q��
���'�;ͻU�R}�� �4��3F�4I��C��+���p�z���j�F������.�\���C�۪U2�8�g
��ߨY�jfR@G��|��;�����]��ۋPln�S9��W������F�o\SA�ŨH#q!Ϻ�
׆��C��j.��a�ｎ�_�����rS:���\�+ަxĸ�����_@�`ɓb{������Y����(�x�|���H^�P�.�j���T���P4a݇�K@"�g����"��z�AɗUK�� P�W��������K��W�n��ǋG���*���G~A�!I��ڱ�P�y��+@�9��gifr��w�:1lvzMF)���Z1>�\]Z�d�>�����q�KI@ٗ?���rg=���$w�~XM�R5AsmS�A`�!����GY�O���)R	���An�W 7���ѡX7��2#�Gy*H�
&rK�/QB����~��x9h_�ֈQ1�_4#0wm�#j��ɧ�1B�_�2�l�N�Jn�)l=��7�*���729q�y7��Z� ��U��Md{���r�y�oM��&<��V����F�Z+p~���'/vz
���o3�X5����Q��'��/��x�sr9�z��Q=[[FΨ��B
��:\��]m�r�#T*����"��y��p�2]3�±}�P�U)����g��ic���\3Y{����z3z5J��i/R\�ݦ�F,W�@�<[s�G>�^� QB��t� ���:Dg?~%�["��cG���/\Ά�m����.D������o�
A8�ٷ���e��6ґ���T�	ٔ�*v�S�l�6�1T�'wR�Va,�ϼ���=;q�{�;�緊ck�����T�77oucU�l[LdK8��)����d0�m�gT�S������� �4x�b[p�'Z�Pkׂ���оUsV�V��-�)��5���+A�N������b���Q�Fj.�"��2�&�qYE�;��p��n����#oY���P�p��͔�.�4�J�����m[k#o�Ŷ��&b�b�c���Pʯ/zĩ���]2;+��d/oۍF!�)ԡ"cB�9ouK�f8��F������������L��)�4�J2QN�S�.�zc�z;f���t����꒍�:��{��yؐ�=]����ژ֡\�ʹ��)���􄕉.V�H��Q�ÎՁ
�G����!���K�n<��.GI�ї�j
C�wCA�����/��^hG�#.k�O��=�c{ jh��~ �/=�Q_�?n��ۓ{��fR���A11�_F�ɺI�}�$\4z�����5�����Uy��>�J팰�����v۞����Q��NQ��J֤�b�0����~|�����u,���K����k0�"%�o��F>����;�I��O����8`}cH�i8��4�U�l0s�M׀ހ��L��w��r\d���>˂��\����׶O��[��&��T��#c=����.�-}���/��&�
ހH�L�Zϝ��9����v$bbډ�^|�ƃ&TƩ���G�>�n6O���0�1�%Ь	��D_� ]I�!D�@+B�˱P���d���{�p	P:�X��ZH԰��9�P�!�Wrz�1��+N#���3"-�jk込mD_ͨ�S�S����Dj�?��K;�B��&I�˾�~Ʉ3~4�!�z��o�
�^�1_k%��"��DAm�兰�Kz&�s$Zh@P는���=֬�øl��^mP�񁓆}�"GAǖ��Ԏ�V�����ׁ��t*9�A ��R)��.+�G�SS�5�آ��)2�ͷ���؈��_��$���5?�zK���o�/���Y��ؼ��(�Td���Q8-OO������Ҙ��ol �����s�F);g�&#`N1�
[�NC*���+�Q��a���HN�c��JU�
h,��WȖ�yA?�6(c!h�aT�%��!��~��d��%��C����v�2��آ3����ä��]�TT�m�|5�Kֈ���)i��J.)� .sŨ��x�PT�ҮT,�Y����/�k}>��rHz��T�������1��-#���� ���ۥ�lxL
�>R1N&�r�gH���+�����@B7~�~�E���A3�h��a�D��A·�J������?_������Ml��$�x��o�Rs�S}�������G5�s�n�ˋUl��,A.�� qJ���@[{��FS	�?:�����ّy���õ�}(��r�I���9�߅T�9�1X#���o@�(p�}oM<�1+��rk.���
6k��Y	0Ŧ%Ǌ���v!�C�6�ԍ�B����/��j��E��K�#>���?����6�ǻf�p ��+��*c�����0"��M�r��4C�+��K�f{���sF���F�<B�k�f�t?��Q8�i��Z��i��}/��e�oOd�}R�,�0�l3���S�RW� ��ѭŰ�C�ahԤ*���G�oX���9��a#���[>��=�p+�]8�6���eQ�OU������=�}��?�8h�=� 1������қ�4����0j7vi$��y X�Ҡ�u&��˛�~��MΜ��5;i�]�yq^yW$b�,��:rY�m��- /6D��?Ԍ�w�����VTH�\�<3��W3{%���;	�ޒ#V�w$�=+�=s�[@�.�&|^����;��;C�`ߎ�._�2.�o�+�Q�$�����E���,	+�A��c���c�ڙ%V[J>KsM:���f+�Fm8��O"v��H�ێ�Z�Tb��F>�����`��ol�Q��]�q7nUC����t�UP�~�ǘ='��1е���Z��G�(��{���|7��h�z�����`��x��q��1����6J���*rm�ÁSkg��>�5��"�b`t�HN�o_B�p! ���P$�͸z
f��i�v��z�q����s���oi�THJ� TX��:$%�}��$��T�kI�t�JSpΊ�S�H��������k��.��y�͔Q�+!��� �Ŭ؏+ñt��ia���7�s��t��l|?0���"%-,Ln#z�_6�x�������Ḵ6������v�s7_p�O1�~滅AQ�P�Anj�;���<QO��G�Wa��޺�+��x6ǂ�,5i�Im����@P��6�y��������Q��Y8�����߯�1X��Fݲ�	����^�5y/�����7'�aX���H��[�g�;�Cr�F��QxfnƱ$���z�&Ze��)��Y��~]-�Zv��`5>K	K�����^e��2�J*.��8&o�l�U*�$}��������h������q<����EPf�y���R�5� ���� �9�%��)�3��ž-��7m*-�f�Xܳ�
s��H5u�&%���D}��0�����p_9/%`���r6I9c�%W���|��x�hK&����Jp�8L!��+m2P����z���/��xgi�	�BnvR6�6�0�P��E��3��tK�`����9T���7�!j7S���ڊ���0���ǅ���X��l�5����ibH�>_�[�FGRV~���[*I��׮�y������8ȟ���s@c-���ڙu��
 �,��c˟���Y���ǁ���%��r�)�o&"J�,�~���
���;ƾp��焻[�ľ�|�r��Bdq�[]��_�'t������G�;���������a���� �,�'B�U�/ʠ�Ù��i�7U��5jx�])��FxFc�Rú' d�}݈L�܈xe�?�-A�Wvp)�MC���x���$eo�񱙽-�\r.�OSm}h�Ie#zي�!���	���N��h(b_զ�����i��_+�V������a<�S�!�:T]�l�-��4
����'p�~��X�t��m�ݛZĈ����o��v�>DJj�^r9�������7Z"\���N��z��QO(�����"+����j�3�j5��5-�-�[���%P�c�E���#�`,�5]��exd��?�K�	��C�>
�w���^,c���`a�ɂ�?0�h�%���Zg�|P`'�Y��%3��!�_A���P4pʂ�ⴾM�}�Dމ8�(".��~6�x����A���a>�� ���㖱2��S�i���/qj��,�[��Is Fb8�sL�*sY$����2>��4z�3�S;m
T=*��Tm�v);��U�����-�n�K��j�D���Uf-�k���PC彊�x���gxS= ���J�4�b�}F��4}a��w	4����A"2�OK*ݐ��lM2,�X�&�9�����bʦ�KX
��zEX���wb�.[��2tk�4߯y)9��w���(��s7�Z�)o��(�pO�mȻ��Kc�85�������
�Y��W�dDҏ����" @�XUݎ���m���e��7��#��/glSM��̭���^�Z�~���B��:���������o�����P��Jx٭=�)i�l�q��g��+�quyʶ�0�Ԑv�JېU�l�6가#؎��Tk
�'�O�T�ܹ��-W����,4��8	�T�)5HkvM����,d
9?�裯$ʧ�etc�2���P��S��y��K�h���۩���_�Z}��k��N�����|�`�n��OP�s�NV{�k�s���m��'@�� ���-䷂�۽��O
���es=�2����AV��/3V��9��B�d\�7d_-�Q�n�O��@J9u�BJ�-?�:w��c{�.�(<ŷK�0���`���&�����4�6�{g���m�^�܅�	��,K|2�׾i��X�?ӓ��?�3��Ԩ�x�(o)��2�W%�y5�_ۿ�ah�\�c�����Qd��n�1�x)bD^VҢf���N��N}��
M���۞u���)؛�m�X������tR�t��{�DC�,����NDt(�!���FE1-�O�i�rV"D��2)_���5��e�x�Σ�0�F�F����;�D����o,��d�>�:P�|��$�X����B2�5��`���g`�:�l��+lF�"� y� ��p}f҅�<j'!O���p��9�z����Ӣ^�{lMn�f�H�]��`1���C+�~0�i�L��r�(o�5]������9c<xs�% �2�9ԟV[�C��1�56���\E���:'9[;��^��m�q�p����+ɰo��<�Y��8�	j�v2l�C��c���J���e+�>�a�t�	��c`�i���^����C�
T��e��r�D�?�W0�DDq�[6�d|f^�Z���7�%�� C��zs����x�C4�n��T�f���C\<pe9��z�l���������n�����e`gV�vFJp�A���đ�^vc_�-'�"�=�	�f�R6��O��*��h��T׳_'�g�ʹw�
�$�݄\O�b�u�J�G���q$�~-���[o}�p���V5�W����舟p���mB�a�g:��&����,����Au5�0�����%�v��ȷ��?%�W�sV�i��Y�f��������V�7Tٸ&=d؃�kvV����IwS?%>���4��o��o�|(�S��	:�X��d�^��Iw?��g5��#H��}��O�'��Y���X񆚳pXQ�2�H�Х���,��Y��H�SG}]a��+�|�hM�h�^���Cm�7�:%�?Y6�1�(��m?���!.�?w��2Q7�*Q����&��
i�u����
k|Jfsd;&V�ގqZܝ���`��a������A�+0�����u�g��9X���Yi-y�;�É����d�(P7��9y��|���xoP�t�czDw�N��T�D��Y�}�nw���G���Ty�L٨��vdolXV`�n��Ծ���?Mr��˟�ͷ��f�w�
�hs��}��TE��E�;�:�@&C$TV�*s�*��`�����j";/�!G�Z�W�*��B���ٳ3���E���A��'���91�Ӏ 2� 5��l�ȵKfδ�HޏW�DժK��K�Ew ���9�3��̃�N^u�b���*ha?�x_��)�=4�r�L�E�b*���NKI�`v����#�CqԖ�+����yx���i��[ֺe���|3��T`��=�$L'�˦�mG�F��7c���i�$��7��&-]���H�p�3�-|j��ϔ*�v��c��z��^��^�����Z�QG����@rg�5@�
�V�-�1�H�9ĺ��{�6��v������\P��!2�z���QwO[��?	jpc�h���볊��n�2Y��o ��[����B6��#�iK�j�~j��$��E�MD E�{5G[���~�ZY_���)�u�-����XHG�����O����@+R�?��`%�E� (��ع��]�b	76e-��n����ko��'� $��ʀ�;���@U�evc|��m����9[Fנ蛼����1E�)hU=UW����'ɏ	��|�)n`g]IacM�2$_`r�`�`*�O'#�fK�֙q�>��'j4ɝc���e�Ra��{f��e#�:���Ò&� +%�?G�s��`OEn��{n~���>����������EF��|I��*�/�s�P�J�pYz�D��3� l�]^�
nZK��T5�;����������%��(���7�i�VIH�sɒ(���S�x%����L//�_]Q���.�&��"����+��e�W�bUpM�G������XI�aAt��<"��c��Fԟ��B8�Rx�<��s���� �j�>�[✆�m�~`ϒ�&�Y���$�?���h��+y�����JLS͈�4�Įy˯LO�M���^#8{T�'��_�� ���s4���F������YV�0�Cj�!���ؖ��W�]1�*Br�|��o���{S�>$����1�K|�Ơ��2��ֲ�.����]��h4�+��������J��	F�z����t���r����;�C]�5H#ϼ�m,�m��Jy�	l�0O���	iIb9�Dx��5��������X���ق�<k�,�v���(��(�ZT*�H��ʒ74)���ʴ�&ˬ0���ڻ�ۘƤPu�x&݃F��?-�;�D��6:��i�џ�*.i���X~�4y����#
�*�O��rMöIV�A�o�t89�7��k�>��q��ҖaWP�����d �*�\	I���0DkQvC@��1ҫ� �`�\���Е�4���-�B#�JwG��qk.LW:9;�N!��'\��Ԥo'` �4��z*��zIoɞ�����g��IE~(Q�TdAk�t|AR�=ʡr�q��#,�R�ް�:�`߳�5PV���0��(ʀ����~�FQ��˔n��=��JkqM��j�%��.wc��>�EJ�I��nU9Щ�v����8��h�{�oܸ��oD7�	2I���,Y�<�C��!tCN��U  x�������2݊����;�Ͱ'j�&sg�Ry�IɃ�в�5=����f���T�F*���7e|��"�i�_qx�U�VLr���YJ@�i�$������6�u�3�匋��&�)��V.��(�j���i�%��:�?~|�g[�*�"dȅ��Q(VwhG���HOXev�!;xi�P/��GK�45Q<3�I�/�l��� RvH1���,�Lm�]��R�~�*MT�eX?��Z��q����ٸϗ��\b�0�A`�1y�৖#[H��b����(���nu�,����wN�����}�t�w�J7�(������t�Fu�	��z"���8��w�˓���i�	����7w!dskT�a �0�a`lB���ȗ.�*��$~c�� /��j��E+�N�[�nb��F�|���q� O�s����|O݂Y��~nZ�x�M_����7��}MKY����
��KH|��#?dN���Bw�Qk���i�1u�`@R�1��ߧC�*��b(l��B�ᶀ��x�rF8ϟ|@�^������JAt*�3-������04q���*gXt��Z�1�P���� `���ca��&����P�]�MW<�N��M�+pEgD�\�v+��: B
Sn˕ց���� ��j��Z�<^�*�˹R�����Z�Jb�u�@��U�y>9�	�\%�����cE�<��i�;����.���sn?u^_��?���*Ed��P�<���l�,<@�&���r���[m�s�^��&���8��3����R6h`�$U�W"�.8�x��/�U����{�^��W�햪x��,���Tv3k�n�~k����w=}�&_S��hG"_E��]g����.a��q9֦�B�Օ.\|�,��-(k�kE����.�D(����V=�53b�cHiݵD����ʺ\DB��X�/�(��;Ω���}��;��f9͗"WQ������wkG0��H������x���%��W�<��5r��]�� )ܓ�F��k�b����|L�տ,�`�$�ڨ���͠��N�;�`d��9@�F�@YW�&<�X�q�C��-*L�u�rǪX.��3�O��|	u;q�M`��Z���b^z�-v�~���ET�.�Hŏ����'�,�JXg 5E�l$��aU�}�S]J��IB�ϸ�c+� �|��2��C��jWޒ\��ְ��T�e�BWM���_�M|@���=�u��K\<�'�q��H��׶OY(w�J�.wI�a�1vE�Ăx(�@��+m!\1��l��hM���;���{G>9S�׻5�p��;�{��pр7�h:�kz�����f�j��Ҭ�
{���6p�½��M=���Z=cyY���_u��Ut3	���Y���w������C�F�Dyڊ���hO��jx��zd�),s������B��7ï�:m�  t����� �9�<����S�і*��n(�=;��L��J�~��6,�8_�=DS�k���	X+��W?�i��崖'��t�9YC�uE�\���������D�S��`�ٺ�!#�'ޔHJ'2:*`�C�Y���+)b{hNޠ�lH��������t|�*�/�]��_�X����l�_�,{�����%�J��@�;a���jbn����bX�r+Y�g��9�>8%�Q�p&�aIk�$��-������|1Lq����q����Z����5�X��l�Q�hW5][���MM���� U�-c��;�X���%c�{��D�����>p�iP�epP�Z�����Џ��'Wm<�b�'��Q����b�v���7gV�ݖ�D���-���UAUziW1@���2�e8���
g�q��0D�rn�v ���w]���#�tܙ/�	R02_ :Ү���Uڲ��t�(�����x�m=�|���p�������}��};B1�n
-��f�C��RX�1�]K�Yn����KD:r����O����'K��dsq���s�����8!�ɭ@H]�		���g	��Hw���2��J�(�p!�y�"7�����\��#8�rꭕQ)&xF%KxXT�m���R����H��+{��L��(�U �ސ��
����"�*] ���4���O�J�ն�j�~�R��������H�.[��0L5���F����c�t��@e ����*��� 9zV�ue!cLbn"��X�.�:��0�b$������N� �*ڢ�Vę�"-��! �/�~�s�xP�ZT�A�G�~�:P������e]�K�_/�E���2�` 3nU��~��a~��PV�InlL�,m���F��K�
��crn��s�L��r��f�O�����oc��>Ơ��`F�NIىU`sX,���jF���Q#hP6���O O��$K���9Ӆ��k�A���Ԍ�3�kݐhe���d�Yp��nꜻЮ3�Rw�C,ё������.M݄�Iɦ�K)�����Ǒ��#��W�AvY���;��9_�".y[��L� ��c}˶�
6�>`���^�n���`��1�w�t����������<ws���/4� ����RSy��%g�)���kR�g�Z�*�^�2&�$��g��������
�U���������l�-�ܧ�i����.iA�iN�dزXp)"Q���{q���ડ�t��Ĕ�� ����ྵ?|;��#>d��=V�,�^����YF�!�
�	�gHQD(��lD�k�z0͈ࡆ2~,f@�����[��q��'�q����jнe<*��0�H���٥��z�22.�LH���|�0���6�6C�BQ����8!�2����6U��+����4]��+n�Q}�������5���}���FO�{:|��Y��dǐ�g�1�@���uG�Į�j��#)M3�Gڭ����L��F��^ߎWx�]��l�E�`O��;u���
h��5�O�Ua�O�s�\�A��e_�m^z�7Fy��̛�����NN�?��Ey�s3��p�b���I]�ƨZ٨B�#!A�����+�8ە
�	ܱwR�۩�R[�٠��7}2��%�ɥ,�Ÿ���Xzt�n��&4���IH���L�2�_R���N�U��A��ن���#���H��A�̖2���@�D��reN�N�lYǚ�8"�p�DEI�l���c�M���޹��),���BY3�4���2aN�ϔʨ~PG>�OMZA�6�~�uK��f�axno@��(��@uv�/���f�zD�)���T���Xۉ[�z'��. �����jnZZ!FKZ�B楲�o5�����$v�TY����D���5_d�c�a���,�&׀mV�Ҡ���S,�<���������f���o�p'r��x������|�hS4�?�����
Y.�|a�/��|����Ŧ= K߿�%4�H�EP�����q-�F�P֬���fK�>L��!�:6��-���W�[rX�sKSh��p�v3�]�\��_��<��T�ۢ�M�=<�V�CX���U14H:����y�
0��UC��H�SY���XA"=�;��C=���p�V�S��M�������;���h�d�?�9AB�ť^�綀�x��
�����^ukoɤ�66�ũ}0\����)@���>�'~ѵz���B��V��N���vt�q�}�M�3�ףbC�uC��l���S��hY���tAҥ���[G�<���|�Hz^���Pg9�$�E��A��'�U1�����o��Q�o���)s3�x�l��m�e�J�쇭r�V^�ǣi�g��������h��UJ��} �p/*3��t/�� \�m��K��Eå�%W���M��+�ʲ��QM)�Ä���&�a��d{!iړՀ�R���4F�|~l|�Nϯ+�����z���t�Ϋb���KQ�b&��|/H��ZUg�iq��)�2����ܫ?a1�+	���+�Fv/NT�K��f��T�<Iy�j0�g�.�`��^�P���㜴�� �p0ӻ�~�	���4G�:�'��sA�N,=�|[� c|��Aw��Vu �� �N嬝�
��LN5CI��""��@��SEp�R�d�m��h~۩���x#����tC6����\�＊:f����p��z�M3)R�Kg6!ىh��쬅�lk�S��w��8*���:�]�㓹�ܾSln 9V(��2�8�n������&��brty��3;���0����6.g�DT��ad[�k�j�nV���$C�]��C��)#
��^�0@�~����a?98���6��y�K�9��Ł�m��u��ي#H]IlE�O,[��{e�����YE�.I��Rb') #���oy��VZ3��G1�s�^M�#c� 
X\��bu�ɦW)E��Qp��s2g�U#���د���gK�|�p�c����h����`�۪u\�����M5|���j9����c��F5Nn���X�8�Չo��X�a� ���3
�_ZzRG!ֈ۽���Ҕ/�UT��Z���Г�����~����+E����L�/�_Z�&/��QQ��y��	P��� ���'C��P9�W����q��=v�ž�7�(��������y��a��|�?��l�k�\TY�	Z�� ���|�FzdACx����K�����·�V4F)O��7}�,�A��u}c�h��2e���⚉?�Ț4'G���a�Ь���U�N9�����k���(��-TJ�V�B�K��y���
���JF�P̆e~M�D
����ƴ�m�K��� E����_^�f�bP�|ʉ�ö�w����,휢a���e���k�O:|��E�_�	 JU�)8M�S)�B5l�&�yJ��C�ޛ��^W��q�k�j�)���jeWOr� &�\se�,��oO��'���:	j]�$9 ��HF�f�b���M6�X|� ��6�(A8�e���"�����ʿ8��Bu��Ka�2BoBf%� ���r���/��1-���.��X�kx�f���pJj>@¹�s}I�Z8�i��U�CGҮe=e�)8H�!�7�6��0�.��"rN=5���Z���`[q�ڎ�����d��\���\��n�Q�[�������S�R��E���/WT������O����b��YO\n��>9�^XD���g�9�0�2~"�w�6@+c�9xMk;�s���>���8i�'̥�e��C#P�1���"4NJa�(,\7���/!�����C�p��U?�����iĕL.�ePHѡ�l"���$dggm�qYL)x��.ou%R'���
Yut�0p��\�%r"�@����O�*%AXX��$| *W2Qq����d�<�L;XIϫ[���6j8���r����5<t�˦����x�+���8�Snji_^��g�ve ������\�?Ҽ?�;�e�������.�/tC��O[W�
���%�.��zM�J�썱c���ܭ�崞�[v���8A^'"	NB�m��B�:h{[��2�M���|F��H-*,�9�c����}��w`4�<�a�O�gyӮk��yos� Ζ�[�$=����'�ZaP��e���=��I}\ƏMK��T`x�a�� �K�{ :z�a&\��ݩ�༕�>хz�)���?h��'��V�W�ɨ��t��Vk7u��f�b99>�h�a���ߵ!�d'ͳ>>���?E���!�pO�E���
��7���p�;�gƔ�s�{���3�e�0����m�I���̓r�"n�D6ؓ{��%O�r��w��)m�o�l�T/ �X5�.��P9/����Etq ��N2[+7�2d�y�2�:�^�S�t���T��FZ�������4F>t���bl�Yަ�S��� �6���z�#��7h��$�5��*:��}oO�����#q�<&��LUz6f<L[K0��t��\S���q %>#���_�59v�x������͓�J�$~�K����I�����9��+�-�(W��\�}�]�����	cՅض��5�.7�S�����w�yu�!/�0ਠ��Z�TB��*�Z�;��]W
��_f��}�jո���k����嗿(ŵ�c���46׭>MG�j�YN��2�s2���m�O�|a��wg����!"�����ƾ`ݥ,�/�}�D��K���?���39���k��3�؟Iq���$�Z�7 �6�����W��m,�g��1�n�rN<f9�=rR��-��!;�;cL������	�=P$�	�͓u�l9�����m��8Xi��)�w���uJ�C�P�7~���"�X�x�j%P`)��J�X�YPP�_���+?qB�_�� ����v0����z�Ǝ���M�9Tn��}�+[�s�$�ص���P�f�V*�O�x�~~\O�(�	���ʌ�'GR�$��H�d���@�؁F"�W}p��JA��wOMr��.9ӑ�>@\do=J��R3�����[�!�l��(m���hK��WԵ�b.�Q�L���v�_a���b���&�/�m�4�1̳f���Tg��2�%�fӿ/D1-����+Rܯ�[��V�Nlj+�X�4[���":bM(2��l���w�
�)���k��Fٟ�c�+f!}���,��.����/#��b
5Ѿ	�f�B�z���Q	<� �Uw&�?_��*�z�7j���0��׌T P��%��w�w�լ0xS�/#��	4u�h��J����J���h�,N��ΪT��tBe�4��|��H��+DvA������?o\	0_ ���9C`\(�e�&\?�QO��f�m{m��]�������������߸FN��]J4�(c) �[*C
BA�װm:�A��������XW:���<��5�2� �5Mj0x�s-���CWr2��м�������tR}�J����zʠ@@1���Ox��_�uAA�/�(�B��5�6�u��C�ێc6ɧ]*N���:��x7��� O���S���m����J�pu!<��z?=����H��O�p��� Ob�� /q{C$�Y����(�F`�,��g��Yk���������7#���x����ED�+�r�#��3J�X g����ӄ�ut��~�@��j�t������
�D���TQs���v�;K.�	�Q{�b\�ÎŬl�7�J|�
�e��ӫ�ıT�A�>јqե��;�L/�ק���'v��1��2��-����~n+�������û�@WT�W����ķ�2t�N���ݶg�%��:�L�>�m|�%dr���-���@�~2 {6G:��o.�q`�bE�r'.�V��;�9���+���z�е[ِ�;H�Y1��Ye�Az�Qt�0�|{�>n��@W
�^�vlqiq�?M]E�;��� ��"k���1�Zh��xDp���ʋ�p�ً;��]>&�'�4����5.Q'Y_�4�n��|���v[�+
ҙ#���r�H��2ƙ;�&y�}�W3o����9��nXd=��4ۑn��F�x�h@�Z�7�ؗ2l��c�ڤ���BW�؋]]0��1Ƞ���}����@b�+onD=�5rBc�z_Ζ�����(j��r?v�{;) Y)Z8�����b��KJ
���"ҷ�0��7�[3������n�p=�������c�_���qQ>e���j['� {/��E��I9BV݊���t��>*�!&agj����]�E�/��a�6���w<������c���r�����N۱��\?;�aD�r�T���Wa8�n1R1d��կZR�|����p	?w��l�{��^e }���lX��(�#���Y���?mR���+&gdq�:}�I?z,k�U�B�	���~�)�<�ZVJa�5�� �=����/RQ��?�h'~�!�Rm�!��t$�cĵ��jĞt.���3�'� b����H�9���W��#>��?���k4{��!z�:��wq�;�8~cu�p�����_
E�8��R��U!�H^���p��'~wr�����=7IP�zܬ��;f9jK�o��^��؃C�S���0k)uE�&]�YÝ�(μ��M831I춠qnʵ�&�k�F����Vk�F���9f1�g���;�IX?v��o�������w�#���b��˟% ��J(Y��S���6 ��ЅǄB��D��Bw(<�Y%1�]�k�0h˰�)��b9��l4wJ�J� ���P�����]`��G`r.���,E�%f����20
=���Ӈ��Jj�,AL�%��G�ʵ�O"W�ŷ������uN�	/h�HG�+njY/�q >}�o$\m��ݴ�pŚ,�)�i &*	�dq�$�� ��)���j]�n�U���������c.���?v~��d�������GD��v��o.R����Ub�y�x}��я0� tA��)�ZD�{\�L�5*p����B�i��.h��TҸ6�:�������j�:�q�v���&�k��^ɰ��>��U.��9	TP�\6"�+��k1=��;���A�d�D�ngK;���KBp��P��ʮ\���XԂ Gǰl��{��)J1I�A�We��>ua6�O4C}�70wb���֢:"�
5�i?E=���]���4u�����zS�?"�Y6��Д8�zfp7Wn�<�&K���U9N
��H�d�B#xG�#�n&���4��S �����N��s��H$S��C��(��m�[�6=�Wh#��PpR��$r̒���E������
�x��Ɩx���;�h�ק2��K]%n�LG��f2~�V�-o�e-�0t�P�h�S���xQ-C1�֤k>��V<��lČh���3�?�բ��}�̦�B5�TX��框�lVh�mU����ϡ�uCi͇Opٻ*Fm���q΀����J���x��\/���mw�	z*ebk�6^V�U1��8љ��˙�Kؗ��H�[�Dy�~�M���^J�)�`P�E����"�����C�ޯ�S��?��W��Y	�������;N��3j�����⛾���d)������(+J>���o�_�D�a��3{��F$J׎��d	�e���"MEmj�u'g��k;@Ҩ��j`}p�d T�5TLǴ�S?�GY�.�^ˁYtH�m!�Ъ5F������ج0��iɧ�I�9Y�q�H�]��]�P�%��z�~�١�1�o�@���^�%٘���f\ �K�K��EY��P� ]2(A.���vq�[q���6嘵�7r�ƅ�������T �4�@� �-�>�5�4>eM�c��GJ�PQ��zeEü��"������"����4ܣ�>��D��"�k�m
ot`� 6�I�E��ՙ	L��R���(S�K Lܧr�x�� (%�}����]w�u���xz�ދ�SJ��H=>`��7U�d�N�	4����8�%�vQQ;�6˞������1�*�4�H�����jBx!d�5����FΫ����!�;sjSt����U/�eh´e�Y��[֕���Nq$�]s�`x�3�� H�%�Z8�EZ���x�X�jtp�GX��t՚�_>.��Zd Y�>�3ӿ�H�.8����k�΂~�-m� i�	��؟��Zp�c����C)U�_�k��/��p�۾�c�+e#c�'(��^޿y������YrV�ޥz��('�+7�e\���������R�}૤�A8�?��=�؉=��
哼ZCN uz�ըD�����T����re��釈�G�o��~���n$@K���q$�� 	��l^�Xm�.=\^Õ��FQa�M����O$:OW�OJ�����־�_5	A��׏��0��Z����'��pB��^ÖS����Ʒ�d��^���%�;�����w)�3w௵�~���|�K�N�ĦeS�v�X��3�A�ӭ&�$��(��e|��.b���6]u�0-��|�]�!�6+���f�7S��	0���󾟆��K�2��s��X�g�,(�ȸ5�d[9f����y?����{���b�E<"tˣϢ����L��3�?���;�@�����n�L߈)�B	�{�(��1�C�dΎ��iQ����;h��-��{a�V�Q4����0wq�-�b1o��ظ8^��?��(E2�EE��E���ij�2�y�yǒ�`��[ ��?���%TX:���TW'D�{J^��&����\c|��_�ԃ�9 V1�f8DM��ŀ�ת�MR�d�m��<���8��(�y�G=D=op3��4��l�<(tE�fј�Ge}�/p�0��f܅��m.��f���nu/*�ǼDq�8SΏ��1�"I"�؜'
��-���CM;;ؘ>����Xڟ�U�_�>��=@�?6g2�,�}A&q�m㙩��{�D)�����9JJ�uTbrR~�ጣ����a��@�K�8f���J��T�L�����[�և��3���'��� �i��c�'�]�(�;̥���
<��`R��c��d9���,Sg7�v��>�e8{gQR���~L�p%�4"��s��7��馢�?��8�xy��nZ��n\��"�&ɸv����`�i��l0hٴ��<����,����nt�=��y[B�ɲ5`��P�qQ��;3�b����"�7�%T�����ѫDDD)D �]����%%�P\���٨Eʔ�
���{��!�`��S�l+�d�v70�����(a�"'��/+���M�Wt9V.�t���ZR:��i�Lj�_�+��p=�������	��Hl���RgKT���Y��U
	GF�cf�l	���׬d��@mZ�K��N����WP��&��Hȸ@߻�f�W�ԥ:턀���ڭ��0]�"N&4��$��r�zF�w����c��)N7�.���T��	3�F�vU>�/.�˸�5�#ߑ�P�0��N�T~i�����'��u_���oL2���*��jG�$5/I���_Z���QR/V�u[G�/a��ƽQ���Ś��{���j�4JB�8��,��
!	�;��쪜HJ7u�2[h�IV�PF���	�j ����oz`O3�����k������K��>��$��(X�悂0>�k��u-U���(*UQ�e+�����Q�=/-�h��7���!�ɱ'��N�[�V(V�L2�%��v�`�]�D�B;�.e�N\O���ٜ�a]7���t�n�(�L`Z��@3�7���0�;*�Y�P;��F �w��EPNѥ�#@��X�&L9�xwOq(s��C�P_~�V�͝��5�P=�ʹ[>����y�q3��s]}!��[h�a�����A?J���$I%4R���f��tE��:7�'�,G����ہ�n�\���C<I*L��`+�i�i��d��5_XҴ��H_�E{=��Wf�}�A9C�z��b�����@>N�Ƒ~���m0���(h���� �)pY_��qwc�4;-�0��m �d;���ii����kX�� А �S:�Ǆ���2�
gq��f� ��z��{��ϵB��3DFt��G\��}��z1	���n�`�~��U�u^�_��k��"��5`�¿��\�>�V4JD{���훐(�AE>T�4o~g��LE�__
���J�/��~,�̈淨Gh����wت'ԕA�1�'�3ǘ�.\h����j}�)�
�i���yJ�o>��jz'M_���1�`��Z��Kom�b�-\*��%��i�1��CjJP�����X(��L�����O����Yԋ�3kwp�#2���)��X�>^��i���h�������˭�u��7Y���BcU���}5����5O��u�D�{l��!et�'%0)i�qu������pF�A�Z��p���³بŇ���� uV,"8�=�/W��%8�f\
�0{���#F��5�F�����az{��WF��#f�p�i�[���Hd�;���������;�U�
�Y�X�]���sٯ�t�1��!-�*���� 
71��KQ\�Pf$��#e'3�o�8f�^|�0M�.�u��.�7���
ߙ���r��O=۴b����JSʥ�\nғe�����p'hu.���ے-A%�j�m�F���	����S-͏]?�un�-�0���
���i�@XE��.�]��XK����>1�F�7����Cfؼ�w=`[��}n
�I:ޛ�9C�QAɲ��n:.�on�F�6"�;?b	6��"���%��ɞi�GLt����܃�����&&��fG��r@:DæЏ�}7�hu�KJB��@`��5���;Z� ⥀�5���W|����%�-p.� �N�@��}q���E������C�a�Í4/�>q}>���tҦИ95��c��,2Ά��cy;^�6��$.#b�r1�h"P���<�%}N_� &.KC9Q��
EtH�"kL��By,�Vۓʱ����"��s�%S�'�ГO�*��g�'[6�&u�����i�lg}�*���Ǻd[���&�zɬp �`��w.�}�F	s�ct �F*�zy�qEz�٫�"��5sþJ�n��@�*`��UI��BܼU�0� �öpm�VO\��P�"t�e	gLq�@兺�lj��%}r:���ê�J�V�|�l�f�ְ�G�'�R��&aK����Ϋ�o���"�)����k�h��	�$S�J��B����v�*��'3ƩJ��n�v������u��ó_��D��Tt�o7[�}ǆ@r�7�ҫ/N��� �5�+cL�2>@+\׭l��s#�X��н�B_��&�ɷ��������{LV�$�wM۵a��o��j���ʊ1ی`��EoDI�i����և�k�#Re=���q󗪐
l���<�!JN�Z�W.�e�@���'y�����.3��`6Pd�v��~�L��;�^(�N�I�����y'����/�,�� �6�����Dk
w����oƬ���jRaw��&LG���'3sҞz� ���w`e~�޻G����:����_A�����Ai�,!|_'��L���݌�u%���>�$Vާ���=�Rj����{�Y��a2nk=��0m��M^x�o�W��&A��X��ou��wG�Q
���g�����Q�)�ֹ�_>Г�a�^@�@��{"�q˜����(�o��c\_-����!E?[���phqj�<�N[R�@S�r�F[ۆY���9:�����嚊�����g�5m?<��!��ǋ�ہ�4�?1\c����Q��@����/�l�]C�]L�4VY���4S�[�J�,{ԑ7���1W���7o��{|ڗ��;�R��������ɒ�-�chW��}��gd�I�N��w��k��Y��Tp��ݔI
h���!�nZ׈Nu�����6^���EU'�!�ۮŊ}6~*��q���^�9w���R}�di}�QVɴ��q!7�ۉ�$��͉Т�n���p���eV������3�1����i��o�K�	,��8�)UK5��貨��o!d��Ac���Dx�/��}�����8\�C���mæoW�YQ�b�T�s9��H�~���������ݍ���ި �W������� ;�H+#��?�M�%N4�<\0K�(I>�$^�7�;�c�ac�N8)b�;A������m-�"���1�`�R�a�����źBŝ�
���Z�V��-<oB�n$���s���79fS��gA<�Q�x��A��Pd)	y TO���V���ucH��P������������n:��d��n�	"8?�)���M���{��v��spAK+F	�ە��E7~P�(ԶMr����!�gZ�!"���PT�]�%�!vݑ� ��M�Cn!1j���+���L����#��6砑�n(f�z�E��-��)T��X��Z+&����`F��B�����Պ e&��}����I��~��NAn�s-y�]��̻�]���7v�ہ�6����s��ˣ^?�3�긔������0�*�|�Z�ZIH�%��FnPNd�[W��ܸ:�a�]���&��Шhˁ�E�y�d��c�W�{��"-�$���It�1��}�� �K�]!q��JK-d[Ig��o�����^�����F`E�r���07��gg�
�'����3�7b0��<�w$��u��Nx�ʜs��>~������[ɛo�~��� �~N���n�S���m�]&Ƣ0��z2/A=5�b��5]��g�/��Q�H'ZT��X�Q����}r��tU�l!���W�RW� DA�*�0
��-hx��;	�_��Α?)��>fև��>�C�߁+|?��S�w��ٕ!�^@�ۄ^��h��z�;�k��5>�N,]~��d��Q�o�Z�@�5ֿ��Z�玷�>�Z��@UB�G���h-��f�&��ճ��в���fdC�������o��d�@V!=�97/��2�`�.9e����Y���j�&��cz�_!����2�L���%.8��*uh̸b�&�x�*�缡k��s�{�V���DKx��,R�Ჽ	�����/T�u��_�릹��9p�-2WOf�#���g+MT��=�m�S����%��gM�欈F�s�+w�E�0����NT���7���O�+�X|��?���H�$:��$�"���3�Ѱ� ��l�i���3Դ467N'E 	]�+r��Od��:2��u&A�FrQԼ�P��/:<�ia����=����V�m���@�5
J^��ٱ��`�����*l�Xr���̹/�#��3��p�<jU+i�%7`v~RШ�$�"I�	+T�E!���s�K; �����o��xE�[>j3ۢ0V1I*��w�-�`�X4�̧e�1t�,�3��܃Bo�j��}
��X���1Uq_!�@��@���V�ݫ�g�tsZ�>1�,F-(D�O,�VƯ?xg1P��,7ēY�(�\�
V�4#��x��[裉�ߞs�F ����ҡe��/\!�8@tL���P�A��G�����?��ip�ϱ�[��"�(�����m�]�PG�T�='a_�@F{��ެT[vF�������Y����t�O�#"��`e��f�o���)�|�S
����b�������:ه!;c���8� cAB��%1@Rvͦ+�M�GJ��#3O'q
�
�u{TЃ�/	���P�	���}<c�dqn�!��ޱ��!~�䶗?H~�$n�r1���boJ4EpT��;:�*���#'y����?$8��BL(T��Q.p�w��-���T3|2�YSs[�K�Du��=�QJ���++�R��Ȑ�yۮY��L�<�ߪNtr�3�筲�c�K3����c�i8^�݂�pù��"�|���������,.ܜ�_������.�
�r$bA�0�_u�z�Jfa�Ιd9�5��SM�g���\|y/���k2n��4eF�`U������%�}/Sa�*�'��'��M�ٌ7���?1�v[-8��&�x���W�F�0���)�0:q��y����I�1�����b���p�����*o;
�r��cv��#Q���R1j!�i@���0-uk��'�B=��ļ�����x� '����:wO�!��I�;���O7�c��?�&;�G�iE�+��f˘.+�6Q�i��Y����Q�<%�\#+�p��(u�}��&L�EΪ�p|�}��� wj �.MI�Dz��p-mS��� ���C�bL`4���ޭc�V��8����=B�� ���D�K�,ĬA�!	߶eS7 h,W{9���ۣ�t�CD��iH�����\��,��X��f������C�O̕�
Ӎ`[�}j�F�C$��ި���w��(G��jX���9U#��L�C�P�,��ɒp%���n�Q_�`A���t���h%7��!���(u�sO�<U~p�R4(qZ��-6{�]5_���-�G�غ��x����`�-��&�bzw`��*�
Iw �u6���Ц�Ȩ5��B��4�-FK5�T�]˜�3&���@��jׯ����ڂ�X�d�>Ɣ�po톊�:rj�U�*q	�l	n�u<���p+J��p�ţ��6���3���ˏZ��C�6�]i������7�����*�!�K	��f('R�xP�~ϰ/�r�c���Ե���X1ϫ�'�yN�R���}?�"�,�*G� ���&��D�X��p����.���%��Wofhaơ<��K�9��y��&*}C|�������yr���/�7�6'a�,��K�N�/,����|�����l��G��� Y�:k�6��7����lş�F�ws�r��^�5���;/*`�������˽s17��6i��{�iMZ����b9?6g�xɊ�����	<�X�޹��Ҽ\'����~sUn?J�V�lQ��������;H�������r1XM�.`���!iP�l�m#`����h �C��Q@
5� ٙ��Ї�I��#W�c6�2�o�QM�{��ϋ1�	Wz�������:x��%��#c�F�2�4���Q��g㽽�!��X�I`qS��<�(P����G�$�A�4��<���(a��z
=v�n5'���-i���A��G"%zj��1Y1�W�i{��k�$f�2���B�g��1b���J��ג||�eH��m��h�&E
�oriQ�5yy0���;Z{�^�jp�	u��S��is�<D���{_�E%��$�⧺�O��g��2��K2ކ!&^�x�;��ign�QO���Gat�_E�4���<}p����j�\��ǂ�W��.�BuX�u����X�>YU8,l���"��w}��.
ΏI����A�t�z�� d	���K�	y+FLKѳ<��*�\~=m��Ѳ�ڇ>
R{���w�[�e$s{�0�J�r������:��H-��B5�;.-��a��&��L!�΁♳0POs�f��QJ�\�s%��q�%o��0���h�f=o43Z�T�"TqU���S���D.6�j�.�9
u��Bt�M�$���+��ci�'�t�o_!�R��/Z��Y�����í��EJ.)��cȷw�֞�N#�a�*x��x����A����}WZ������=�:'���c�4Rl�Š�$(��>5�]�n�h�?g_��H�^�'�2�E��*U`"��e�m�-�JKG�,r����M�̦�)r@z,��D���
����'����"���Y����+�Q��E�M=�`�<M+�8ǭp�V�3D3Ȇ�7m��)��!��dԮO*@�����A��E��W1#MIU2�������4`L]��g���d��
�k���$��g솽�k�������;���l��!3�۠]>���g0@��RW��<� ���,z��re��|h��r� Du7���eS����~2]۬�>]w����<5�
F��o�W�.�u�� $���Z9 n[�FX�4j�:�ј6�!���˰0�xkV�� E�jC�\c�T�vwT2[�`r�
���I$弬�)>����9:Y@�g�R��pgv���+���l�rdOHM�@�&�e��_6�z�'�?�[�V�-��<Z�P���P�2���l;��S��sLdl�7d[C�s&�/�_Xme��-s��Y����o�R�u�/1@p�t�I�O
��s�~��2D�I邼�^~�2U���ͦ\K�s<솫(�a���bӱ�%���2nr�5[�/N-IJ�|��,,r����p�5Q�j���O>r�P�2����+�x1���4����V2�dk���k{j7�گ?6�L�Ӓ���\d�:��"�s��k��'��`���0���Y�C$ʶ�C�f�����q�x����a�?@���SPj���-�~eB��[}�K�l*,mQNؒ	y��b��mIT��W���ȋ�����ʪϽ �tA�vA��=�$�FX�Z����X��"yd-�)Dt���䤶�O9�<8q�a��T�u���s��_�:k�Z��Q�x��	��KI���-H��
�G��P���G��ƀe�e�d��ېy�8�cŗ4��xC�i��&V�"�ß���	ͨ=���)�Pg����l�%�\,�!5<}��r����<m@ O�����+�f*���fH�n�'ei����'C����h��S.(�
,y��7���>�S����Y����Xz���T�5�Hh�a�~vn�DG!���m�scN�$c�қ�q�xD$.��=������*o7�w�2�ެH�#���2bSL�@��j[�im>D(�b��^y�	g\��fJ�&�q5b>%��i�M�i� �m¦�z�2�:�ߕ덙��nȁ|��L�I/���ۦI{v���K�K��7[��k�O��m�78�H<���tb�"Y?yy&�&==�v�?VY>����-��:ET�_��.��:.Um~֐�����/i�%�� c������3m�j'?��8�	ǷM;!���,��
��ү��� �q�����c���YQ���#�FI:��B��\� �-c����5�������e:���r1�R��Y� +�����c�f�&��j��s=�U!���N�3ާ-���A{��e�hn��'�sDyD�OmL���>�ͭ�5��y��[}	��?̿�Q|1_W^�x~/J�V�sRWu�H��N���ea�<kٛ�񤆴죟w��4�>a|MG�(b�\ُ���Q9.	z�_F�|�dK��[TP!q=
�o���Ku����]�^�����+��9T2�'�c�;
��}�%�y�k1��
��Bh)wv H��n%: �YA����<.�?Y�ެs�p�d�\+�7�ͽ�5�`�������~c{��X��� �������=uP��p�:���s����E�j�p��]��U)haDH[�d��.�����<�~π%V�i���K�+0_���mm)c��y�
!��#�I�
��!}٩�-PO��.ͻFF|5�	4���;��{����.;�����c����F�|��<<�� �'s�E�f?RB�����n�ۊ�-��:�x��!�'a�[3�Q��͹T�T�rݙLC��J���d>�|y�Y�J`{�=>kĖz�ps�樑2vs��`��?3N�L�q8��k)�'�hunKc<]1i�WF�<���T�b��*�v/��_�P��X�W�4҇x���F�!�S��8d^�09���Ⲯ���M2@�6D�ݾ-�5 /ߋ�x�J�W-��0"G�F���ۨr՞V�Ub;������Ɲ�h��U5�>#o`>�|>�4�D�]������5Q	lબ<���$Ÿ�K�N��e{��*g<��M���)U�6������6��%! ~�mI���Q�)�gK?�E�����	a��b�Յ��}`"[!d��>�OUy� S�,1⓪Ԗ�k��h~ =&s�cX ��(z� ��[�$���%���Xq��YB0·�<�Ned`�jA֎X�<�=���*ZI�L�ϟϝ��GWۊX �e]6L:r]�uS�d���κ�Ryt��58o����MB�����C�γ�z���n�����B�s�
��� ?� ����[���Q�>�3@��ֿ,��|���h���܂�Ĝ"w��b��p�T����f̎�<���g�*�1�F�*���A��$�3�*�8g��$\~У�=����Q������bC$"s��)��!�D�����xD܆;Sw���;�����X+%�~�f�=񄈔��(�T~��k��	ӧc��C������o�������q�����0=�\�d�I�l�zZ?���Y�(�:M���Ioڂ�_�#�;Ђ�����F ���[�o��!g5ȼ�}�q0'౱�2n�ö��3��K�ֿ�j醹� g��)��a����n&�Eר#�8l.�p!�t��������=��5� �	��@�Ạhk�/�U��$������{�_a�U�O2�t�M����ҷ�|�'�(#�	�<v�@��n�7��b��?�%���h����x��!ǃ�[�%��X��dG�0	'��m�ʖ73�w�J������C�����\� ��%��%L�'	�W�l,�d�`��#����V�e)�'�l�'1��w��]������/�1`+����~u�]Sv �Ʃ=}_�]�8�Ğ5f�}[E�5 j��:�AX���-:��	��fjk����x9bE����(����� �k���l���&ǒ����Ae���>9Cn�b=J^���߶���{<�w+S�1q>b�|V�Ӕe$\wa��Pn�3�5�y>���y�n�v�`�pԡ��+R�E6���~0�/�m1��e�WǳR�(��2��R.�]����#8��@Gy����'V��	$��H!o1��<���v��fޅA"9lT�����4c?�k�}p}���	_:���]�/�:9����-^�B#eHa/���]�h��b�9��������sK�Ǘ�շ��������0d�EDܬl�XH2�/�D��x�~�Ҩ�-jK�P��!��v��a�*�C瑯�G-����6q�F�x�m�")����3�p��Kh��Rw�d�Hݧ�/!�M21�lR�V�b�������L��V���t�(�t�&\�+vW���N�#�d�RV�g2���?��e�9��NW��P#N�����4|zPF�Ln��w@��U�oT.A�v���>i���%Q�3�QK C]��,��� �3K�\A���f��O�{�A���X����y�^�Ow�T��--���!"2R)d���ݫrҶ������m��YJ<�4��U�#C���ڌ�,1�9�U�&��":���}��=��&�e�����(h܈���P^~o��t�#w���6C�m��rp{p��%0�O��pB���?���?Ř9�Z ��G�PZ��4Y~�@����T�Egq�k�1�dB���m��i=-�q䫧��j^F���rLT����V��V���Vnw�U��Q������E:.0�KݘOģ��N��?��^�
�4h�'P˜b�n�-B�j���^!�!:Zi�EI��E�d'{).#z]�jB�n4�YL3��A,I�J������T�>*��S`�������T�ܴ������2�0 ��sh��P��a�hUxв�~E#z�%͌�>�����2h��nl��p� Q�
tWK\*x�xrX�U{hXT���Q����<�;��w���t>�� ������-��57�p�&r�P@I�
})8J�T�w|��/��֪��?��ņ�@�����$�6O�c������!�^����[U���Ր�3n��0ژ�0b_�� $���B��I��� ��)�H숷��V���D���^!O\��>�cr��6'nW��30D������a���P��C��[U������x4�{ٯ'`	Mg�!|�QK��x����E�&`}���C>�_��Aw�k2,�k1��x,����9�[���r���[!d�O�����6�x�2���c &O�ŗ[䲙�P4������U���WnV"G�J�b0��4bGh.�;I��@8bAn%�?�������S�o�i�N@V|3��/�x7*��w0�qbIr�`��Uv�CN�V�򮝋�NK#�&a��t�J����	4?G"��j�̈́y��VL�����R���<����B��Y� �%�C~�֊v�W�aeO,�#�l)ֽ@�3U�%������2�s�m_�z���9���`�^u�z�(Pnq��;�Q����[���,�B����O�ij0��"l���:c�惍�+֊Kj�=dˀ=��v;'>����h/�D-�
��®'tF��Y���}Շ��~�����KW��J��ĝ?�,1�o��ފ`II]�f�����F��)�RO�p�[��8l�Dh/�2��iڇ�ޏ��V�$��L���^V����U��V�����@vD����E���x��Gh����Wc�0���T��`w��Q��w��5�cT8y.$�ÇuB+(��F/k����Ҁ>���!��H$�� ���1��*�Y��H!������V�%�<{����s���h�x˖������qg�u�RA�� -m��C�nS��{}d�$W9�����W����/�n�\H2h��xAY����3���f��:t�q�o��ߟ�|(N:�OX��I���`�P, ��wnM�O~��x,"��J�����;������i�){$"k�=����/7g�D����_�O���M6>�c_�u�&{��G��L��n8�ߏM��3Δ�q8�iqaT瘰��<T2*8�D���A
$įs�ڍ�[S���K��R��E�+)�S�yN�R����Y0� S*�
�aqe6uG�K�[8뀈��N7���m_��L`5;��ɛ�L�t���nX6�ǉN��
|���D}�Y�I�,�Z	4Z$�豵�����(��^CxØN��F�X&�E	��Ǳ�7~�����ׯ��yX�����Ae�*rQ��x��%�LgN����!�
{�����R
�Ş��L�b�kƯ�fl�%I�90v�z ������P�"[|L�1s���'^Jة�EH�#*P��������Z� ��������Hb�-^hę�z� ���/x3���}����i@���VC�S�7x�h�#1��dP�[�Ioo��0���h؈1#������s�l�]w��qn���Լ4<��=�̞ aHoC��7J����K��0�D�,��������8�}���]򙏧;h��U>�+=���|���x����R82�.	sឬٵ+��$�2��2�c<�2����@	���2��k#Jk�$u>-#�{O� �p̦�y��N����5����;r�Q���<׿�\�CmZ�{������c���^�����{f��`�rk	���Մ)��y�:
�&�\�Xw�^�k/a�N���QǦ���ǽ{��N�J��#�/|��rN��7�y������e��#�1[5P�1�R �y��c������I�.La�^A�;���^!{��fs��U��������ȶL�5��C���=��
(����.xv�¸#�9�.��$
�~�����>n_-T�¹�EW:H>=���k�O�-37r�%�Z���邏��Vm.Äh��^*=uK`H�HA�~�䖛�u}� �u�
Y,Cc�'����!J;�O�#����vib`x&��<�nP�ť�9fK��\u�����Z��G�M��'��ձ�k��2��+2�hW���d�S;�$��	0j����?�|�BO�I֘�P#I�OR�,ז(�5(�\ ���l�(��N�&W�r�4Y�/d'������D��Hh��%���|d8���K�i��􇖞��\c���d���5Ox!�H����J,�m�Xwa�]N�h}S�.��/CԒ���o[���5ӗ��0	Գ�)��{�D�B1�?���F�ϕ߽�Ȱ��%�e$���q��g� 4Gäo�g�jS��t��6�tj"Tog�������|��`ʂ��8k "�%������>��hZؓ("�OI�O���"�=��>)��N*N�A^�૵0s �22fy�񝸍�;�}��l�iW�^�T�:v�&��Q�����QN$Vʽi�?9��sf-���ZB�N������u��#Ui�*���;�WY)[Xz������9.��J/hӜ�CN��������x�i�Wh"rP�hs��9S�w�*Z�R��і�N�q*=�S�����
e���!cO���xR �U�����Z[?6��O��:��GYpe	z �`x��"�.��h�D�D��%�1W��w\~2xZ{O|nu�iZq�f�kq	���YyM�p���q�#�A>��m�|���2�*Վ(W'�Q�
�
���턻��Sl�W������4�r�.