��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>��`HX����5a8Sjf\�|Vv <��Ɣ�����hd��� *~b�<��G4�aY�M�z31�5s�Ԑ�s��
:���j���w�BĠ�9f�i��?!�B,�PAuO2ua�a�{��m	RK��̓��<��e?�2��ֺ��^��}J� 0-C�"��h%��p�V�}yKn�A�C��%ꠢ<���xL{���41����N�|Y"r�k.����d�M�tK �Qx�Vqx���6(��1&lS�?⽽Ol�}1����$D�tҏ�fĉ�x����=���7뎍3��-�Ua|�q0�mWG�|�t�� +:�P��ěD�	h��w0�Yv#%;M��y�@�#ʧ
����``�ѥ}q�:m��vW$!߬�`7{z�O�1�P9�s)ߧS�i�mrZ)ܔ�!H.�r��ٶ�2�ej���D�}4���y݃(gJ�̋�Ǿ��i1��/��/0�`�ZR�lx�N�
R�[g�(T�;����"��(���P!Զ_�Y�7��.\�<qY�|�����s�R�����I�o�RO�[3(L_��p��#�����}V��ut�>�`Ν��<��`�b�ӝ�-��)WV��P�I(L��|��N�D��;������؉W�G��A���Q�����n���
x]��{�en"�ˁ�߸�91�=ﴙ�u�-���FcX�y��.󍭵(UM[��[���,�l��=�btDJJC$AO�)��q!k'��iT�@f�\ 	��G������h�J(��r��5���F��O�s'��ML9-qH�T���w3�q��1��9�i��L-��Q�D�.��ZZֶK��S
O��9��j�A���0��G~u���A&y<��|
���\Ʀc�-�����!vQ<G�4㵪(�ћCJ�4|���5{�8wR��q��B:x��זJ>���kf����C:1�O���3�o�j�,jp_�}�>ړ w���P*x���C�6����	,&#+��۫6�����>5эS����-@~0�Gj�ko�R<�/J��*Ĉr�9�-�p���g܊�7;�){�\o8�:�)`tD�����ZeD�j��"���ʢIG��Ь>�WTz�@��ֱ%�)�{�9O��[�׋p��3����w��]�("ؙ���o�t��e����IV�W����q�K�SMd,�yv�k� !���Q�W�q]�����j�l{Dd2v���S6�z���lb߷gU��r-*�(��حM���0�rd�=dz��޾�MQ���J?Ou�(�S*���j�b�5�M �cr��C�|�-s�5�Oٟ�����A��o��p��n<L ^Ʌ�׶#Y�l��ચs��٨�DL���{����V@��n�x͍t��iYc.���"��
�W�|:�Vf���"h`
w�Pz��%;I=?�6��OFz�Ŗ-+�@o���;=��H�L����2��w����ޅ,G�,Q���ľ�,@l��xt���*��~T��Gb�o��d��\@���l�L���%��ܸq�a����Xl�P�V�&.fc�*�v���tS��Ც[������f0��TՒ;,��nkLfz�,ʺ���B&���p�v}�I�܊�*O�v�5l�!Uc-����Z�7���R�+hg�G�YL`��+B�\�W���1\�b� Y�$�.O�G�pMkA�g_�] �����5U|�p� �;�	���C{��XV�ÙWR{!�Ĺ%6
P`/z�n��;��.O�S�W� VOլ�����?09�^�	%x�w�5�v���S� <��Y��Bf��F�-ï��b0:�/龪 �X�{g��ˍ�3�	s-aM�5����Jy}�-�lǟ��<�u���4jG��g���zI��v���p�MeSW��f[Z*�5�[��.!ڬX|A�+E$>V�����H��O�PW�B>u!��,�]$:97�Z;�p(�-|���{%�� �v0�Z�T�z-��#�<r����*�)��#��,��eUB1K��j)�LV)�ƴd@KW'�;���9�4&��)�W*�3���j���M�9��s�E.��Ή�_ٺ������0#����dt}�=y�W��y*cjSC_��̐	�^)��m�#�2��V�(}H�Fӣ��s�9��5_<�5�vy8��n��GeL�f�����ʨ��*M���n��e	�Ct�V�0�``��I�����Xy��0zx��,F�]��x���#����RH��~J<ݤ���9q��G����o�i���<�9Y+4�����D��k�7�BUL�*	��������y'�]��;��*��]Ak2m�����v)�Z,�[�W!܊G�}����"K��c��]��v�O� e�8�H7�˄F���4h��ϱ쁊�W�#gh�4�r�F<4	��Ƣ^�ǆ��j��F���o^����AN��4���ȶ7A^|q�S�hX���q2��;e/E�Ү��Gm��ɺ�':�(������]�N��njVyv�����+MY�z�n�7u�ݾ�v��~U����0ݴ��R���2��z�Wr��a'EqfΓ���Q> ;���'����	_������V��!�0�3���l�3jI�-dDŊ� ф �T�!T��(uT��6�<���6e��@ܴ��!�D_nlSd�.F���!e��Z;��  �}��N�*:"&-�k����xBn��jj�4�[�Y�?7���`F��U�V�d��)#z�����"$� .���QHbT���&��|!ECw��}#�ry�x��guP�g0|��s�r�+K���[ŤWD-e��9�94�H��7�Sm2�z!���=8U��V�B��Z�]be�,�����^���_��j��	C5�<���K��XE>F$Bx��7��̠߄[C�)�ӿP�z)�d���Ҍ����`g�kҥq�z1�ZY��ׂ�����s$8?�;��7��5�_[	��!�ͩ��S蜈�ڹ���qVh_8m�nO����ų�@;#����>�e���h��y�p5�čr��&N��JÒ�~��W��g!��)I�}2#ŴSJ8��,3�,¦*�OdlRb�=%���8),(s�>��b�U����d_�U���HX�_��а7c�m�ӻ�V������hf
��i)�B-�_ּ����@*��*������C�DHI�f��Ɔ���xKHD��H��p2�F�E���"�`����8>������c��@:��[#�`�������˵�0'��T��A�jM��p90���eL�PF�/�v.Ԇ�N���G���52���%Sjh�>��%�3�;\{�u�)1m��I���1;Z�O��+���S'��V�(����+c��ax�K�jS�c� ��'��	Z���X��@���E*��(;��M����ă[��4���Vx���?������ߕ�Fd�r;��)k&]�7$ɷ�9����Ε� Rއ7��f���ZH��?�o1�	��n;O�ɦ��0	���T�nx�o˴�K��5$ӥJ�J&���>���{$���G���E�53|�����L\���.Y\w��}������+�?�4OP��b)�:�VY7ص �=�����L	l\��������Θ�T�~�P27�LѨu[�bxA�����]
���C�#T����>_�6�wY��[��Y��QK�8��	��C��J�UT�Ʃ-dVC�Ɩ�3E=��沒y��+�w9ǳ�i�mE���>����[Qmz�<#�r-�w�;�A��"LR�wgd�ڌ����D�KSRL}�4
+́Aq N+99~=�c���#�X�M>��<P����H��Ns�6�Φ�j���߂7�k`}5���J���?�Ѩ��e�F1C�Vh��K�x���!~܋���u���=�k���)��6~���VJ�"�K�ޤ��=��ԧǣ̵�`��Rر��7����jU��5|�au�^�Kd2Z���8�M����в��	^0���D##;F�f=�Pg����;ݚ�4����/⴬�U,<J� 1��yz����y�qB2�Q9[R�M������W�_����	�#�[�n�M�|����{�u���0�R��l�N�ӿ���E�a\̀��,�G#�Y��Q���sR�Ə� ��癍���m[�2�y9�F�	���niB�k}��-���O
 �e��נ���mr	B��>\a��}�2²�=�o-;�浄���Ï''z����&O��$���=.����;�+�)L�O�Y����%��Ms����iLhJp�Ǟ>Ya֘g�(��{F��WJ�c����7K>�z7��~PSd@�J�W�~�+��G�"���x�Sr�A㎶�0������a�^�����5Ongb\���j۴xRn���y
���M�P�l���>hc{!��FN�-�ŀ�Vɚ`��O�%�ө⿾�R��l+�}�IV�k��ϱ�$Jd���$Mg�,B�Bpu��B/a�X?��o�,9�.��3v���q`��6���'�g�;�6�A_���<�/5�:������luz0��uWz��sH�'g�Ǵ���y�=<A}<����-UU�'(>E0�8���qb��� �t E�������*�i{�R�$��>f�����Z���,�d�8ģڗ��3�m��ěr��Z��Զ�R�5v�@���3����Zx��`+�[M���g�8��rO(� 4Q��7W-�3dP���~�����;�����1_K��.���;j����dy�$!���%z��S�I��+�L4ke>�Ն\��9_)��w:��+�U�����>m�fo�9�^��;�E\��EX]�g�s��K�*-y���>���D�x�rQ|�#���Q��7��YO�XٹG#t����7�p��u��(�0���v� �z��y�1o�0\e���Ũp���:�h�1�āo�C���_��lZ��	_�
$N���9��A��0�k�fx��;`=��v��縘�;�3(��Z��gH�.���N��>�K����X
Aʣ���U3��ۗ6���:��k �	��0�=��jm��,DB���Y��tM�mhUm\B+�]`���2Ԛ���pL�E4t�I���F�1����!u��rE���9%O�_\�y��D�*�|o ��i��,��V,uw�˺t`�"��ѐs�䉭s�u��swzjή��Zޏ���7�,n�����ޓL�������E;�h�n�3h�mFs�!FGF)����Rը5E�qJ�h"q�O�G��?�����o7���;�(I36y�O���?���b&<҂Yc� �}�ܢ�pc��sC�EO���>Q�P�C��|7�$(����*�s�wd�>Y��"����YRMh+�̏z��T�=�q�����}d%�d����<�wL��gV�W�*Z���Z
?@�m��
�n�Db�9���LKDˉSd���#����=�}�Y�~�k:�l����t�E����Nζ��
�^ ��C:��c�I]�)�Y���'��}��I=���*m3���f]�>���c�4����a?���a��%�r ���r���r�I��P�^w�U9Z�F/���ÉP���`!Љ{"<��G�ڰ�P��ʺ���pd��5h\�)�?BQ�7�"-��'�|]R�E��ܔ=^��5젺���%kE���"w�;��lv�h���p�I�a�yN����`�PH�����#�m�m��#Ɲ�c�f�j�d���௨ x��%�M�ߣ'�^q���7�d�.�������g<ń�J��L�Єfn�|��\���C���}�4���Ja��e/��#��$���,��C��;~Ԕ�����(��o�^��q��΋�_إ5�x|o?�-�E<V�Pm�^��H��!�cv}�r]�0a6�5���)���|}3v����P�X4�~;gO_H��.���+�%�+�9Q���V�|���?�.�jF�O�UY1�W�n��8T�ͅ���V�͵�a6�	R�E��B{�3�cx��A����5�O/ߙ��p�7�(�O�	l�0'�a�Q�Z�b���|����ra�qnL�d'��� ٭��n3X�;���U��đ:/a�갋��n�($$n�Qa#^�#�d'��e�Cx ��GK�����P��M+?�7�Jtn�$U$<ͭ�/(N���"4�H�����I.�s��i�˩�B���K��]G��4g j��(��u�O*@��%Y����J��!�i��"��d&$D�p��~�69��ܤ{#�a�L	��J��e�S\��,N9����
��̒�����cd2ؑUf�;:?�+��I���f��IWv�72\H�@�ކ�̝M-
I����n�-2o�6\7���US�n;�	���ǞF#��9W�EI���+��_�7���Q�IU�u�.�s�3 
�M�{װ��2��9�l�ߥ�!vG��M	��%�Aj��%<�8KB1�v<���J���$��*Xtٴ�|m#�(T�J�躃k�|o)��͡�dU���W�@଍�d���?�&�w��H�e�YP/�(�b�+�ϪO�x"��A)6� L����mz���
fe�53o����N��+��5�߂�o�*�H���
�t�FQ��6K����2�S�af%��A[;Hٝa�zv���x̀͘W3q��ȋ����l/]:WJ/��k'�5����7̗�[�k�Ѵ�_�eD�l��.%�CD6zn�"�ܠ�2pJ�T�!��ӺѺz��^�$r-,��:�<X��%a�9���q��������n���2��p*#�A��<\�6�񱢜f��B�nf�t�d=��oy����J&n��#R(�ut8��11�e������d:�K-�`��i@���u�@����'C\�V|�,�MCȎR}�H*��8~h��).��Ut!ʪ�����~�����F=~@D��N��v�N�z]r��O&#���x����¦��}�bX�f��*���z*�5���\
��S]�E�'�g���vˉh�LX�b�˦��7	J}��<�A���&�T~��c�\h�R|��Iae<U��6XJӰ����<у���'��D�<$�$��_c�+��JiȚ�6��;�%��m��?9����(��b`�i��1�8���l(�B��M�0'�)���G"���`4��d�`�?3�K�4mC��U]��?��9���(_'15�z���#LT����m�,�'��v���}\F����}���Wb����F�lJ�ՠG��~��v�����D��`lǈ�獜��Hoxq3��@���_�9�Б�����R��
�<U�G4��\��0��ϗ�(z�C;�,�K��}�I<���OT��)��m��:^^�YG�ϝ�77�_�'?	�t.����C���8sޗ�"6?���>�*��߁�*ߋQ."��Y�<��:#�y�E�q=���ǟ��u�IO�na�ޖ���s.4�݈�!%5[l�W^$����;�us�ML��9���chpD��+�!gp�(=m� �ʤ��;�"������V8#]����,��7
�����`5@����g�_�E�f�;q}���I�>�,x�Z��qe��b���CV��?!e,��7O���~y��9NF'�� Q����Zen� �I���Ѽ�E&��([��?���^���ѩ8�%��-7[��N���ۙ�f��~�#S�����`��؈~�UX���R�2k�`��Hܰ*����W�P#G�̷��vL��?�8�?K�9~���gt���V�=�I���g� �}�_yH�m�yfV��1���*v��h�4}�X�����v7�~��q��%�b�&3��fc���V�l.��}���� ޻�b�#��hW6"#�飠����@�=�-�i�ǦH�w�x�<�m@�(��A�a��N-ÿ�}{�Ck%Ҁ�8�sMk�zt����;�jd1��6u^��J��0Rr��!���A��^HU�w���?�f
��R��^�-�H�wy���ɗF{�C��BGՊP$lG�XbԐ-�٪���0��-�O��$�Ѵ+�	hd�l���Qs��>����T�3*�M/�/��>����")����E="|�'l=K�9�����SB
H���շػ`��(m�vj����Ǫ���xZD*��$��f�إ�9�ߏz�h�	�o�*����1�+��6`���e����߰���O(կj�z�9ü�:�l�{�����4�7�6l����R�t�Cq�#��s�5rܥۻ���isԭKX'�f��aAq8Mt�<Dә�jj��b;��U4sl����E4=a.�KA��~F]�X��޹��Pe�f5T������=������f�Q"
�hƒ��f_��A
˚���� p�oI�VA�^��[9��|z��_F2 #���������?"���o����:b�Rݨ�f�Ӿ����W�b�Z���v�Mm@t��y�ȳ�U�G�Y6�� ����,u�Q8u^�A0(Sz��<�$Ko�JC�XÙa�`tEe=����="�4���]��:�7��Ϋ�;.�iUļ�n�~k���M�as��jyaC�?to���Eq������2L�S��l�"��5�F�.s*m�nE���T���q��FZ-�:Y�C�G�,V;���d��>v�&��:a@M�؛�;�;v��z�2�Ea�@�v��,��@K���\����-7�щ8NsTk#&�Moό8��p���C�qɯ�U���A⽖)�Fu����vZSv�β�%�?��ٰ���e$ϪeIXO�l_�[~�?�A`>�)��S 6M?!Z�y���K��B����Sg-dn�f��a���_5�d[�y�=�pa�x���hxc��L̀}^��W�%���ܯ��t��?o��о����l�朁�� ��e�c�x��U�N&C+(jl�/%i_r���/��L�snX��u�^r�	����6��p����߯q����0�<����.�Q�EP�e�,�<'p�f^�������r]���sO]��O%��8Qt�J1�O���{D�c���&tޥ�^�i�р�� ��݄��?��{��՘	��2;z?�b�%\t�^)�$�7���~ ���v?@�C#uއ��|�~��It�K��q�T-��w�(��l��h���T����@ԙ�cV������4�����V�����4�}N|�򦈹����}e�z�n*z������<Wo��Te3�(m��/K��ճ��	��Vx"ʉ���;�`T����fV ��f�PR�����e�+!'���ܦ��� Y	`�:� �l���1A^ӗ��5�3�5ǈ;"y�l��G�¢�^��La2:�����<0|�>�a�ɡp���$!��JEj��T���1u�-�V��5��x�������z��F��2��0\��J�h�:��⛩e�sf����V�Z0�j���0�� �?*�ل��+N�d�5s���*,��TxZu� �$	P��y�kU^��'�RJ��L]w�>�ӳH�՗WV�}���7"��qR��2���^>w�l٬ۤ8-d�(k�֪�cPV�j�H�f4y��W,�'P�ZA�f'���u�Ğ��.D� ��`g�e�-���	To��Z��#�=�9���y7~3N�}gjq��:L�9ٲ=������f�n��$��U�u�Z��6�2B���Hf����ENNGD+��("Y���X��x��`���I� :?�D�O���hUVA�a ���5������t��r3�zVh�AM��fE������kv�4�"��!�|W���!��Ǹ���+'�z�Pʈ�����;������~�-����-G\�e���U#C��67n��J0� $��^����gHA-�]����SK��1�I=�^�!���;ِy���3j-_8-����[D+*�O���
�e�&�F�c���B�+�z�a�2KLM�Қ]�l�p�p�/*��PU�ä���Q�d t%<���?*�಻e�fr�^��[�G5�����a&�L�8�͡���a�
n	�4�[ݬcn¨������fOpp�oK�����*XQR���������b ��'H8s���+�;,�V����� ���&�L�u�{��Z�Xu���m/� �-M�����y��x�nG��oc����nw�����zYp�i[y�~I{��t��Z�������i�o�����y�,7q}I�Ʃ��w�8nK��K$����O-��A�P2�_83�r��$w��p4�_��;��(A1�����a�3(h2���]F��~��X��*÷d�c�.8 c���%v��)�T��^)#�;ls��id7
`ݼR,���øj���,`�	-�g5��Z�(��W��X�Y�)<�0��R��������>VS�;T�ӟ��$,�U�� ]����
�%���uR�h���nk!��!>��ۉ���!�#r�i����E[�ʍw��og{/k@���y�����h���톏����4��YO@�x��G m�R}�~�	U������b��:���[�5������mwtƘ\*bC�}!��S�F�f������Hw���:�E5���l�:�N"����x'�}�,L�I�"{�¦ѳ
��Ee��Hoõf1I\h/�{�9&�����j��(�3m�O�$P��/� ج�w���Z]7�b��:m�7��=5�9��a͚7�a0���/ED3"��r&@�d5Ί��W�j������� �dP̀�جf"�%�@[�*Έ3@�0��^Og)3<��(!��+=�����y~0Xa|R��i�M�^�%i�3 <�)�I5��WΑ#��Qp��ۂ�{��a~0���m~ ꈮ��H�v�^�]����`w;��W�I��U�֍�v< C��{ɇ��3g�YW���l�&+w�- f*sj%�=	�Б��D�5hX	 ��|GU]L��wJ�jqv���Jx�UՉ����D\�(ј΁�8�.	ݠ�#�������-�tP�6��E�ۮ�-��}���a��x�&��{���DG����xBy9W}�����p�3d���%�Q��`�׵��(�W��]�
t`���y�"[ڒ��m�|W��w"�{#�t��-C���S��_��?�Y�]mXu���.��K[5�Om��FQ2A������M*�p�@���k�l�z���c3Ҵt�wD��/��1��**�$���s3��Q*�x�Bn/S����]&�/.���0`L���'�l\���86�U�=3֟R�{.��.�Ph%�ZhqNd��ˤF�^�lN�7����+�JN�u��N�Pj�2� �?��9����!��#�,Rb;y�uh7�}��MW����D@��.XP2DD&��g���y�����\�w�sqi�c�g�B�nB_T�f�obj�	%|�>+�h@�=�� �%CsG��U*�\0���U���a�ƈQ��6z\|a-RSHĻU9^)�����E�X�B�2�ŠZf�~m���`"��l2�Fqg뛁�����a�iƝS�4yi;ߎ��K�G
�~w3���x~�BU�O�if���Ir��*�v�}1�I}֎�I�0+�s���2��i|.iG�fQ���F���#��T��@��F��{e�f�%���a0/�A�G=O�"hQ؄F���|�ն��~X/�����v��ݨ|t���$�x��ڴ�9"UˡtB�� �7p�2�kf���\k@��T�g�S6{��sbYPI���n쩌���Ut�IF���(m�>��t���̙���4�H�6�.���כB�;����3u�&����*��3�
���Q�y��s��_�Ф���HӢ�*���2A�TR�"4|�թ�I2�ϕ���I�`���}�n�bU�������0���(�-B��x�jE:$���x��� Mנ��e���l<3��=�ͷ�����oz�	7�V��u��7�ԩ���.j�K����K���Y�oQÆ�̷�1�;���t���8�d.h����u��w���r/�@��ORμ�[e���Wʿy��w:B�)H�2�!X�s�&�,�U��SS>�]�ӆ��'��,	1�JO}Y$��� �<�����|�a�p�e��V�%.$��4����zM4�.<��mZ�������b�|TLl�I���6=ʩ4�:(Jjl�j󜜷�oӊ�r�y;�f�3�:b!B2�Ӱ|������ll"l�n�V��`�0<:d�ب]Ie��`w,��7F�-V��\��&bF� %�?
/�ݷ�+����"{���p�����~x�:�ӝ>����@>�;��@��.{�Htal��?9���TR 3z<Y�-+��2��CM$�P>D�{���C��&2?U����*" xy4�e��,�_�&|C��ȴ��7� ���#5�x��� W����gW���9tK@� ����*x;�bP�e<��ۃ?�x����Hњ�%՗�Cd����Ұya8�s�X��?w�g�-,�A��l�(�p�
���l�U+c'��Ӆ3�C��!x�^?/;�T$��SX�vc����Ѡ�$>��H]
������x}���N�)eqR�����ύa-�C�}��^�4��6jI�b=>�H�*�����_��s�ŷ�ln`n�^{�7ᵙ�ր�6�'����>�p=� �y�(�3�?�=��B`^ID�/|$L5Ы��
�0":7��j�_G�qr�����V�[@c
��2���c�����=�0#�j��W��@&R � �uW��w��^gq�R9v��6��9Mi��n�g3���1J���,k[�ImT�5��T��:<԰f���U��$!� ��V����Vqs`�J7����L�)B���e���-����O�L���5��m�s~e�KrFӒ��Dv[�mQ�y�!��j��h�����ghl�>�s6�ױy�A��;)w
��z=�~��]��~;����>�����c-Q��Y�*�̫g����OY6�f#�H��+=�"�k�K'��jU��N�Q�_�T�S-�<��P��{Y&ׇ�����H����%�[�'���Y���B�Ȁ��Lb���>�EVٯ���;*����D�T�6��ZոE��C���G"���X
�V��T�7�7�%k��3�Lw�*0]Ѫ���"����J�͉�ګ=O��<{⨈��R��iJ]���Ma�_��B2̧��*'�c����	��_+�	����[���Vb6�3�zE^]nL*�Dg�i��|*V���k��H�W	����]װ�%��������d/��ޤf���"��Fl�ge<��%��ʃ{x��? ?���s�cV���(���
��v�Ds����6L���#OXcn��Mv��)R�wI)�N�����]�y�z�h[��X�^-^ȸ�'���c��GU�a��\�@:@���h��+d{�0�`��'��Cr7�D���J[u��S3Q?O���?����3���}�!���7���k8���g��%�%�HA��3���`j}�J͚���
sΏ��9H}K�5��ۣ��)�K�_���U��>�/u�m[��9/�!y��!�e�h�)���=y}6���l�S	�R��kH�>���3�ѵ�GN�K';#�G��[E
YqK��v��T�����;�����T߲�F}�e~kx��5��행Z��C)�RI�_���K�nR��=�$����X#h�tѶ�e�XTa�w�N���Y��7	f��QB��+�-���(tOߩ�뎠�x{����������j�(9k	7�>6`3ֽ�h���R���H�B��\��瞛�b�3��}�<R��ŰR�bVs���|��n�p ���7�����M�Wf�M�uǧ�̧\����c���O�c��=S��A2f��f�+h�[�3��nҴ,M����wܾo�>��l�?ˋ��:T������:�h��!��ߩ�wK�i����$�6�0�	�hT��+���OV6�� ��ys��ȿN!ۦ=��p����O�J/ҁ�1����R�j�=���h�i Fi�i�2}�zMP��Xu���>��2�5�úk�c�V�����r�\~��%@���us�^Z{�ۈ���� �>��Sv!��U��\�[���3�2�xL?��e��z[<�.�aw��dtu�u=�� �p�6�\ڣnY��B
�ᚮ��e+[!f���@G�� ���?`y��@����������q�zC�+��[P��`��7N�NH�&J�MbZ~S�i�D@r�ީ@��,�����ۄߠ������ޝxt_���&�|���
��ەuLo'A�O�`��-}k��تOV�D�˼���ǀ�E/b�<��N�\�n�!긟Ē���q9�E���e�lX�|q�EGYH�n���N�Uw
�#�=#�ȝ1`��*�6t sҵ�U��d&z��oM�Ww=��o��~ İ��-Q�2��+��c7��7�R����NE���C4�ODHs�� �l�(�� ��*D�G4���f)�uM�����p�� iN1�W�=��{��V�N�<@��(��)}�O�P�1XC�Q5��	��2xE,,�_��d�j��o�+H�`"�1��<w�}O�%�45dV���P���tޒM��N�ۗ��-�p��>V�8�{������>�i��pߑ�~�ɖ� ����{��&]�Y��E2<�Ĕۄ�Fc>r#kw�jJPXe�5�ך��y�����E���*@h�lX���g-ۯtDv�$�r�˞�}&�f+y���ʬa`U.�rjo��}����*���&̎���TU�H:�Ev�q
��y�H��~ٌзޱ��z�n"����*u.֙��i�ԫPD��~��R?&)�Tq���6�<�6a�`����҂[���S 6l����;v�N�mM'~[\��!�s�?��ڤ�OV���j! �	�H�T/mT�vZ�iǧ���G��lu�9j�u:�6�-z��Q}zVt:Go+y|�z&F)3AF�\]&\l����,i��j_3�z?u�š��]Pz��X!@B,RU�j�e�����(�2��ٿ��8�:'Jx�9���ݰ�8�L�1�K�t ���.���u�&����M� g����~�ˇ��N�D�L�����t�u�}!D1�N��9t��D�ʏ<��j�I]P��}U6��n51�b�f�!��2�|�>]E�V���@C1-HG��d̑��mGA����yGɤM�)�����"�5�+&u	8O �K�.SR4\Em�u� :����D ���(�ae��g4�;�*ʹH�
�����C9�r�qWSa|c��w܆3���E?������Y�ittR��3V����~uTAҴ϶q(�~n��G���d��$�(���x��giL=dHO[�
���[Q��l�VA5W:�r_��4�����:Ԋ<��fs����V}��Yf\��b�.ƨ�k���$������&�׊�Č��ҫmԃ_:�t��f�^�[��IO��n�y���HmWJ|s9�˪A}��:.�	�����B�߲|
�!�)*G�zPSg�O֡n��F���R�2���I�t�?8����oA;M��f7��C~7eYg��f�~��@�,V7�,��J�,��|"V���ʏ&\ʾ����hb�I����P{y'd��710l��duS���.�%�n�U�W�pj�h�]�;뿲IC^����M�D�G�/q�3�5K� �:#���bTs�tf�e�tX6�{�a���bJ.=���V��lv�68c'2(��I���&������w�e�7o�l�c:��ԥ�4�i2���7	q�5E[cl�1����k���Ě�vv'�X�Px�X"�F�T�|g8��� #=nK)1f�g��b4��P佅��y��A������д�X�(��/8���7J���\��>[�B��3\�G�:n9H̊"��֫cF	�i� �%�iTk�ʿ�|��c�E|9"�x`0x����!w����8��g ��z�R�/L��X�<-p��̤����ʄsķ�1�!P˖�N�	�a9ꈻ��t�He���%�1%15F
��iq��J�\�0� }8�'�b�,�)a��G����=��zR��E|p��h�~΂n�B�̠8�wc)r�|��cQF+��/�:0<�m���SQ{�!����HUXI��{�r�ݠ��1�rhAz�����&��(M��A����1L7�\�O }�qG�?���̸3���($�kN}U�57( �7��U�ƫ9��ۏ��;�I<��Xs��\�@o���y�	�6�6QLN�<<�����*�h\n��y�J`�G�W��Np�8S�����K�5 �Q�u��(���Ƣg�(��; ��o[�X�)�3�I_�nA��� ���噠\�	4~�T��8��K��sUY!V��U%nu0=�����u��q�}�v�w����X�q�x���<f�@���a�>��/������d���/#Q�� R��p">�l��:�J���"�QGK����M�c��פ

�`f����WS3������:1R0���a��}��$#1~�BL�8Jm�瀀�Px��]� {ɕj�d��ךɝ���� w�q�ofG���3���X{!�f!�
	N��g">F�+Z9�0��2���?��!��04Q�*䨬�~�y��d������޿��*�XT|�o:�`֠GBn��p��)��G�QIc���'�/��L�eⅸ\�N�W��aF�3������C2&�o�������Uŧ/*I"�f����"\��}=	��f���9"��|n��KoSz���V�m�O�����J=��ZQ���'8x7ߨ�F�*_ݫ��b�T�<w�q͘p����씈w�������I�d�8h1r!�C���"��~&�Q*q���#�F�fx����z��7�kGI�5$��JA �ΨtU���ci֎?�:")�LNb��QC:�	[�a��a%�UT �񨴋�/�'pW��5PS��~��F-�NJ������C��oT�t���N^v1&�p5���������ٛ����S�:;��y!!�ȭ�n���y���|铙mv)�m@>Y�ŀ��S")O�wB�w_�p�,���,�����(����QF-�BPJ���.6➗f�LIx�/�8�j���+@O�]q#��:��,���C��~;�ޔ&`b-�}��e�S�gN|�
�2�\� D��`�0T���W;�df�P�&��^[o�[/ߠ���O��
�t���F`B�`r��p8��%��?��
��Y$8��L;��>t6���l���)����"װͮ�������ZX+�f��o���$��<�����O�<p����b�K~�"���؟b:Ք�{�"�h]���`���$�p����
��·�Ѿ	x����jD�(${$����)/ (�w�2���X�ZV�X�����2�kA��y��6�W5�}e��Ն��Y�"�-�8�I?f�hFnSQO���a��f�6nw7��CȮ�{r'�-w�U��V�s�y�3lɑ�L�c#��U(W�����&��}@�K����n��>�s �R�����:���6�颎��W�z�����^��o5�N@Ńc�z���k[B�uK5�v�K�ġe�d��Am�w
�V���&(h�����^�o�����--��Y�(*Uh�cr�&9���kiP���վ:�W��5Kڊ�ɱ}Y��n�<���u�I��i7]\�"��9��r����o����O��DI#�~U-��P�櫒G;jʯk���*�sx��x �Ck%25"d���Q	��s@�.�x|9�Z�_��#�=�hSKC�`A'��>��GeiU��f3cap.�[F���f1����v�.y���<8��iMzS#�~�q�|���cz�4�?�s/#��Q������l1S�t��X��ʧ`�0���U*�Ov�y�j?Ǜwe����J0�˳.D7U�I�t��#_9�&<��M��pF3�
>��8��P�La^<��^�;x;i���r���6�7�\���G� ������&�t�N���]���N�'���kT?}��l�6/����\�z��z{�o�1755�B*{[6|n����|T���d�l�ɓ�':�:f��F�e��4Wӊt��({=a�O�:9��>l�a;S�g}�����3ߕ�[*��\����hݪ2ӵ��_�#��녁�C�.p ɏ_�uȕT��*�F!����;�g"7����=6Q��HH�4-^�-*x��ǞM���3.�(HT�Q�y�G��\���[���a��HV:X�ށ�vk��J�l��ȸqt�A�p�cڄ���6]%���^�[��!�zz��^����|M�S�Z�������5ư���N�}MB�����������%��d'�r�х���>WV_X4q�~�*��}cpR��chq:vu����@D��::CD,�'�n���{��!���>qm~�K1�tB��L��#��x�z�d�4����G,A�-��B)�Ho]w�a���\'�tl��6��N��'�:$'ȫ?B�*��6 �v㓇�ڲ�Ҟ@c��[�/�a�c�=��#��l���	�gv�;Ϸ-'Tso�"� �%ϔt}Cz/����T_�����^]Uʰ��gY(L��l��t�5I`���1�N
m �#�#s�aA��*�9���-5�7�<o�J�?���BvͲRA� ���=�kצ~}>g/,4Ui�i��t�u,����)D��������l��>v}	������ޚ0�����?
Cv&��R�"#k!?�d���	���,@m�)Y\B��r�n*���L�m4�A	��6��9���z��Q��?�������h�>:�I��t�-m,�K���;���p1�1]3'�t�v6+��܆����v������5����o�oE�3C�!�vj���Aц@�11�	�y�����<�5a�2��ho�m�+V���T��%��fM]ʄ��ij���B�D���}Ϣ�F�n���R�=�n���P��A�� ����oA��"������g�T��jh.GG�E�m�R�)�.��\e�4��;���~P��,�o�(Mh�>�@7�O:0��#�=���[����Xp��{9��� _��A�N�H�"O���~mrS�����q���[���%�����:B��kGF	��9ڀ?ᩌ���E���m��Hݠ��	��Uݶ$�!�6��^�/QA։�'N7a1?�(B���*V{�QL2_c�D�<�e/��+�Gx]_�:�>��z�'��ˡi�{(�ZC�J���E?�^�H���sl0��y`DD�>����vjv4�O�P|���(J$�!#��)nƦ	�\&�)�K\_㴖W oz���U88w��C�o(x��v�혐w�ݭ]�7Ar�[\D����������J2ZynS�
B�c �p�3���	I�A B�%1�:`��g'�/L�V��m\"h�Z�`��*�U͛����N.Z�!8	�9�쎒��'6�5��Ǘ:NŅ��u��E#l�^�Z9��%�r1�1,P�f��� (�0�N1 g���rU�l���� �MA��$�+
o�K{�7Ǚ����0\�⇻���!@{�S�������*�X杖Q�H�:�����%:��aa_D*'��D����a���-m��q�~�
 q '�فws<љM�_C �$=�t�nei�^�Uzf�(��?����)b��{�І5s�oV�^%$B�hOO�Iya�#x�~�� p�  e��6=9�6~�>�����l�G
�![�RY�5�:ay�_I� �ɃR뀆�������E�[txy�K5��BB?�!C�4#]�-G��!&����Қ#��}��ͱ�t��Q�<�i\!o�ӄ�MW��/�#��G6�;IaXw�jګ@7��ŶxD�_uH軈�~ȡ �]2(�w�q��MF���Tf�~H�..�{�j�K��w��uM��kx"ߐe�4l_xsib(�Ծgr&�L�`V��}�8����I��F{ӁK����,t��P��!�Vw��X�p�1�AV@��q�i��X�O���9�����RH[l	�nl"nU�ӷc���V��Gd������NuqdI��w�-��dn��o�/�\��vi�P�,��✛V�_�R?v�}�h���ٷ,�0����k�¦2��3
�m���P ���"ïV�9���4��rB��2M?�$�MtQ���s ��Y� �Ԋ�]�A;��8~�=���IQn���d��h�W�9*�F�.vM���Q�4�l��ɦ��s�D�H�U�A�y�e�dsU��uf�l��qƿ���¡Qf�-����sC:�|9Hb+b��-�>��6��p����>d��i�2v��@q�fǈt7L=�w-$��g��<�-���,~E4I��;�����"
�0���D9Ӗ:Fޢ����ꩮ9�P�4���㭏�&�s���O:7vHYŞ#�X争�XiYwaǡ�M��Q���x0O\��x��x͔��y��jq���uk����;5���a{#�O�����FrG�"6�<J�aI�e�!�3Y��&ЗԮB��Zoáj��O��4���f
C�Ih���񁓵��_f���h�CQ/{�qTa��[A�K�-	�^`�r��R�D ��W�L���B&g��j�2��"pM��8F���G��#��o�*��t3}'�fg����Cy���cW�,'��@ͼ�� �cI+�/�|�ng�/�+J��i�6f62)y�A���*}(C�DR��[�.,��_�K�|�\/6��_��"��)���F�c�S��IZ�U5�Z����F�"�O�p�"���w�������|DuZ��L����%p����[6��FH(}C�_!�mGr>��+i�Ok����K�݌Š��z��[���*��n�3	2���	�
$M�z-�����jbn�|16�1f;͠:�uG��؃�j.G�lN��b�B�X��Nt4�v�Oa�]%���d�҇�ţ�A��3��@��o�mF���?�I�9��o|^U���a�~੥n~���d旌)���;�V,����e��w�7Xz�ޡǹ(k.U�j�9wl8qT��p&� �9P�&������u;�&#<8��*^ye��P�Y�%`��L'@xڂ`�XYjoľ61A�JE_Q�e�����ʉU)�Hb7,�n���3� �ܬ�D�����+u�ԇPHy|��"p"c�WYs���mQ�I���G��,���=B����M�������l�([���ܑ��׬�F�N��E(a�z݅�OM�G��=�F�7àW���;�*&�!όk�t��2�U�!�m>z)vp/O�Q6�!�8L][������,y,�8i�L�����XN�pb�-hS�9|����C;I�_�R�U����Q��D����� �o��x�{�۟+�;h ��b����8t�����*�Nr�4$S��M'y|��Bn��|��.�]M�; =�h��\�>���~]�B��?��D##��~���@�j�:�H��x�0m�!/Xb'�2p�.���Q[�%WX�:�gwv��V�h#jv�����Oذ�Z+�
�hۍ2fFUsl:q>z=O����mZ��/J�7��h�K1����hM���e9�y"R|~���Y�;S�����8P������u�H��;%UU���%�\�~w��	���1�u!IƐZ��v{J['�ߟ��c����־dXhB`0WB�z��1^rT�|9�'Y�P���m,~aۦ�2�{������3��"�����Ke����w�h��� �~�85��2��0�7}�M�[|���̸�(����F��l�5��=���ɖ{�B�xɿHީ�������3 _�ϝ��@+}yU�F�6%d̥9:�f~��ˬ�M�08���S��Z�]nz`�8G6|�{Ci��Au�	���S�y|��pHLΠ��n
���d��8q����;�P`x��"��2�H��pN�:��Ix��I;!�7����4���ᗱ�Ul��_�.��4����鱢Y�F����ǥ�Ah�r[4JsE�G�,}_�BO`\�J�`� h���`���m2b&5����j�oW���Sl'�y�h:R�u���h'��(o�����m���������|[���t���x���2��*RIFxĄ����ta:�DOxU����
�KS�N�eH�h�(EV�0d�ֳ�C�L��3