��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|��I�ɖ���˽�+]�Jf��N����2��@����甘������A5�N���n�nD����n���p�+^�T�������'��������c(�Lb|?�0����gb��o�YtJ��%-��8��7�A���**�Ǡ��2;),�,���G�� N�����k�V$}zt�� s$�@��Q^�L���n��A!�~��(��2���tz��J&S�NK�s�p7l�2H6�-;%+����{$�	2�s%����}b����ɽ@ߚ������F���A�~w�������GBĐ&���O�w�K���U�3cZ&w� E�Ȱ�Cx���eV��Ҩ`�n@�d�V"q�Hf��#v=o����nX�t��� ����Z��d ��o�!��9s���T�&q��7@{��N��r�U��N�{bXa�m��U��45���^�y#$�^��SBՄ?�!��u�b�`�F�n��I!��C)̓-W Y�h�^ �xR��?X{~`�S��\,P��Ƙ�u���6Љ"��)�KʼS��/�J]�e���A{<�~��U��c�[���������5v9!��ُ�_�)�[˖�����_4���A1Vkw��D|jj���RؑE��� l����3E2�+����GR.ሥK}P˅_Ə:fma�����A�Z�7�	7�Re
Vɿ�<�+�\	EL\{tH�j��8ޠ���͜�(,<���7>�Rɲ�����bʲ �ɜFξ��QB����j��vSK��a���:����*��R�1̱���g��?�,�ܨUo��-uw��L�1�n�?p�N��T���K�=�1�A�0��d��Jl�����i�+���8�W4��������EPk#��#M���@�� \���l>�+͔��� � ~^��E���p�,��	Ĺ��aQ��>qC�����
fi�0�N�.��1Z��E�|��©��^�'9�j��� C"�C��m�0v��������]�?uHB8{B��6!�a�^��gk�#�����y�;�bM�~AʀŬ�8���1ձW��!y"�+�v��WA.��/A��;UEI�7 �A�9T���zN��O�"��~�9:V1���^Q#��[Po��UrNE����f����#���by�9�� �Uȕja�H ]�Q������%?� ���Y��՗h��B2���th�#��oΖ�d'6����Nk�5��g0(M�Î.C]!4AH��|�(x�\�-���[w���]�u��ٍ33iZ��_[o^��n�7�Õ�<��).'#)��^*kX�Z����d��(��ӆ��Ǭf^���9PEb��J�4t�M�]gJ��yL�$K�i��"`p� �a'e�m���4)�*!��)ˎ�cs����_z���׳�X�֢oHMW�l
�sBF��b$����M\��J�Ũ0Ω �튳�_�:x4�v���s"P�1��Vt��V�Nl��@�q�0��ys�G�J�;0{N��w�θ�:��3��xY���j��t�"��d��g���������G�E���'�^�O���s��^Z��Y� �vpD=Ӏ�=s��!�`�qXM�H�c�|�A�ì��2<���`1&� ���t��@C�G�3����ϊc�u�����5��c�Յ͙Z���P=�$g�Ib���z�x�?�o{������
T\��)��p���D)p7�d�`�̖���w:�R/rU�F��V����pz�xKOx<��{�q��c��Ә���`�<��搧�m�cm�����șQF1�����_�,�@,��J<Cԇ���tCO����~�xn߷��$"��A�IWO[�Uǡm�^?
+a�	�w��⛮��+�^!oUsLS�\�0���ńf;�����y\Ug�[��+t�>5�T�����z��6	�+����t�:��Ľ~�:\��������*{�~4�N�^�"d�|�ǯ�i��>�]�	����_��d�\������S��Pb�'X+-�Φ5�����M�y@�tf@)ƙ�1���R�B�F�es�M������<�Yme��}�K� ��vT�>i_*oT�&YG{~��S�K��n�[��m�:v4���%�_6c�|@���{�|��PQD����`s^+	���;A�b�~��F~�̓��P���zE�z�3IӎQ���1x��n�9�P��pё�*l��^mN4;���t-�4iЉ2)��Gn	�E!�az�.��������s��c��_
��Bv�K=l�bO>���Hh��q�W�b<(
�j�Z��^ƃ9��XMf:�Z�
�^w����ŭ4�N����U�8��r�6m����|��t�Z��]��X�'`�KΔ�.�t/����m�Ȁ�r�WuK��\8W���h���x��J���L.&�d]�4N�b��h �1Z1jw���9>�A�SE(��C���3?[���yb�)��?.e�-��B��%�np9����P-J,��Q����}�$q0W3�6M�Ȁ�\M���[� ��P��Ȗ,�"�X�ç�C��n�w �_<�߸!;2���b/���-�~�֍=�0�M�0�l�������\g#����R#� @S&�{�;�V�]�)�K��!���W���'�9�̘
� WR���R1	�J�ӿ ���JPC���鑱��a(v.�`-��?�1V���0�ff���}�����G"w��d��t�����ϗv~K�6iv�""��|�< $ ���;���I�ͫ�|���n���CU�,VdN�`���k��V韀�h`��;P��Kp��k��I�]D���ޯ#�(j��L����,F!+x`�� D�}��G���m��^a��twRj�ɔ�82���è�o�t
�Р������\���g	,`��AaO�0b��*�����ֶ m(z��߃�R@)	70RԼs^Q�������؃���~�w���R�4�ځpER��変�!5�N�ZB}��×0�)��;�Mr��`��x��1�9Mlu��is,�cw5h��)�z�p�'��	��u��k�m�Dm��xx��6w�6��16���6O�5 J4.��u��m�I7�@v�
�]xY�7�D��$4���A��nT��xM#����H�w��%�:WD�l�c)�N��zP�>��t=�s����Wp�ϝ'�yXm0ft�wA��s�YY��R6���&�=YXDW��߽�v�i�@�����cN�j�FO�:�4;!�kr.�s�|o�G����(>�r��,�3�0]>{��g�T���F�0�b����{�q��@��<����%�F�.�w�<�C	a�������5�'q%8� w����_��ʐƲ{�H�D)�3�N�btea�8�������N94����0��n)��B,Φ?�"U�7�ĤA�� >էX����*����oˈh��B}��v��������E��S�������X�;i��l����y�ΟX���n{XD�H�1�G<��N�Uvq�l�<�(.��k�V���,����� ��ۢPZ����d�ۂi�� +����W�J�S ��J�f�x���ȈR��= �K�����a.�(��*�o(?Y] 6���K���[>�k�	{6JW�׎a��)cAOdI�C'�&'�,Q1�@ir���`=���ݽ5!���F�uE{�<v�' ��$t<�rH#��9b��Z��Z]�v�H�8��-�'�)�,��j�