��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|>�qT��>�z��
�����|�L愫�H��ɺ�a��w��$�YF���bںM_���,�0>��z���H���P�0��C���[�;vJ׭Rj.�
�1�?��a�IX��U�ܰꨮ�\��;(�Ee�-V���%��S�I)?i�^�r0H������S¹�=��OF�=H<P�}�4�����%"�fv�׍E�體|+�����Ǝ(���Y�����:5' -���\��
:�NdP- �LtC�ܑ�5�8C���&�+�����4�����*��K�!�P���RW6��b�#��}��cb�N��2����Vs�X���[�iX�K�Z�1�K,�*<�~8s����w�|G0�����~l	^��C d=h�~�������?�C'�W��(�qTKB=���������$�`� ��J�XX��Fp�/D��m����Év|�Mڶ��@��L��M��]�?�egUM��9�@���c���D�Ն4�͎F�_���u!d.��88��Dp��N��l�{�7CKA���yc�b� �<���uvaݦ���@>ry}���^;
�[����^I���˘b���>���<qW{]	�����x��f+�=����!�GOD 6�Kݝ������R���]�3~�}]�@��)=!U�AL��Bwh&�4,��K�����w���]x�4�DM�*�c�790k�������T;���{�{���LM�B�b�� �����B�O��)L"�<j�e )��R��D��Ƹ:�k��h]Y�z���B�d+<�G+4���A�# �J�لɞ�Kj������nU���N�� w7���G�E5��D�$��4�"R(Ŝj�chU��a,�.~4� �_������[�rfᓊq�Qܯ��e�
ڐ�J���ό�6]�pd��p�!�[�k�J!
����,d�f�Ʉ"��3��Ac Alџ���<�݃�q3L����s��"@<�E���P`M�
��h�q=�11�1��J�c{�!����Y9���^SV��2�sv��馞�Cvz_d�Gབྷ{���FHk"+<��f��5p���*%~�A�`�6uXT89��h���"�����������u=�V��S"aqc3��_�����m_��x]�
Wu�mv��f��p}f��M=�!�xv@��@���F�Q��p̌�mx5������C�)&�V�y�E�ٙ��������m?t<)]�R̲I��k��þ�F���3_-l�U��؅C���5V�"ݜZi�Vm{�j���%�`�jt��|Ko+���[�߄_T+Dy 1��6�/�һ���P�f�Pl�����莈��ԗ���ޓ~4`wyBȬeP���{p�v�bX�-\Ka�ɑ���GSD�o����΂�e��?�yۖH8$�c�Ƀ��7ϊ�E�f�J��<tw��#e��請�Е�rx�9���lW^�z��8�wM���Y@�LVǉ�T�bC��[�����E穒{���n�t��^D�*%�H�c��=��ؠ�; ��.�D0���ȿ	����D=X��oz]{���s��{l����&ORՇ#���<��ΌR�j��Rfs]Ө:�F
���Օu!���|OG�����K�m��!Z|���ga��lA}�/��
��Q���)��f.ZL�.B)c8�G�dݽ�p7$��&���"�G~;�ev�Ѥ�w�8�gvڻr��`��/T"��g/\��t�LQR�Qc�+��x��}���)��K�(8��	U�n��ʣ[�=}�;�t�U�砙��v�f�;'��7�^�b�b�$������e�9[��ce�%?sŭQ�FţG�^
]e�����B����.��'z#N��W]�[� Dːt@���1Qn|};Rx~�L�W7�v�[��Q���9���[�B�s�m䚀���O�(T���$��b���EK��|G��כe�L}��� 4�ə�ӵM�T:|w;0����\cL�z,	���j���`-����6��AZ�x����@�ѿtx�>1���F���� �r~��#::�J*��}�	�|�H�ت���T��,G��>��f�_�/.H��8D
2��q��7�J<#��[��X�x��z{kX�4d�`��]�+� �^9��u}�sc����R\n�4����]�8���:bLn�����UV����Q��i9�7R�<�#�_eT����� ��r����]W�������3c3 h�5�.ˊ"R<}e���c+��>��;�����AW��EX�0?t�^b�&[Lg ���>a�2h��`+�V}%g$�)�jt�};��VoR��:�
�6z˅�#�QA�&�@/�92M`�$f"��6�/&�S��M�'�A��ꠧ`����U	���$Fk�T*a�RjPxf����Z����{�r3
��\������G+� �p����|_�ߎf��3g�,�J�SU��'��Y�'�)W�s�49����`������|"�	�7�i�|~l��6� ��sf�ѝj��l�ȧ�%$a��KH�^+S!��g�N	O���fM6QL�zZdT�3�/?$+���bu�4�s�y!ݗ������I��dOɒ{���d����V��ykz���4��1C�[�$�6�Ǒ��N^��޺G�o�2��9-� ��-|w�>O�<z�W�V4����4�W�`�r�R���BM���Q< ��C��+�bh���1xz�`]���q�\���9�@͚q�{�#�ߟ��� Cn��1lJ1>(8�Ȯ�ԭW�y�	>�mر��D�	 �<嘦pP\03�	�P�Trn��$��+��Md``o]��+3*��/�Cv8������s�wd3-��	�|ME�ќے�5��-�M�Dzq6C_U+�1Oм2���%�\$��`�X>�R�[�����^�qE�+�ѡ"H~J�VRPߨ�C�G���$`m�PUs,�0��3��~�R�aC�e�F�3�J�B�VL2�)!d�1#�{Cb��t�.�YPĉ�)C�&'�^�z����K��h�@g�b����1�n�7苑̗k�Sԫ�����Љ���[�rH�i�}��%Y�B���=�$�!�yD�A�ژ���\���b��Ww.��_h<m��7�V^fi=�Kǡ"ҡ�7BG*B�X ��Y~��ؠ�+���Y{�P����eL��̤�2��}����A�����x����vY��O�|��t���"�@mC�7'ӂ����/��"���{�gqF�s�3�
�df���a"fא��Q?0Tj��6bC<P�+���&�{*�F����I��X�Bq�r@������>U���uJ_�%^~M5? c��d�8,d���9�G��#����C�֌�� %�r����P�^ƨc��H���vF��������6��-Z��c��A]��v,��q�� C������otm� �f����T�*)�Y��l'R���#�'~q�Д�}XƱ	�&d����(@INά�9�4r	d	�0�4O��?�G��_*�:ý,�������3�Z����"�ob�O(d�܃'9i�{>Uw{��l�6b
�y�4�@��z�b��l���69���%��V�ST�X�>���*z�zZ���Ko�d�9Z�F��U~{����^����u(�g@ \��QR��/B�a�WFm�%�}� ��&r��6B�)�h�+�q�NȻ�Xg͏W-��a
������m�d��g9�]`��W]��5G��s�_��|�QЄ���4�3	H#