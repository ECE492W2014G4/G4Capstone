��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P��v�"<ߞ��&'��k%P碶�R�ӣ�sĞ������FY&K�KFPT:�=�����"|h��ඣ ;��M��ͳ!\���yڮP�$
y�dIGR�TBY�dz��ԧ` «�'Hр���<<�̂�( 7���y�f�IT�߁�!�F
�w�����/+~S�,��J�3l�}� F`d� ��w!����j�%���pY���(Q
z�|�^"aq����m��f(��e����` &�U����qN�!������-�Y�1h���rhOTϮ�%�a�;�O�7Ρ/�;�a j�cyV�j)'m����������>��O�]�����i�yG��-��#I��_�.�:�n�Z/�4��g,٬ ��[��F:犫�;KF(��Ĉ6g����2��H�,¾��'������3&��$��Kœ�aC�HMr-3[�d��ا�}��K1c'	���a����_2<{.��s���hY�0K�e�N���]L�C�a*w��.<]v$�^8CRG!hi)�Nb��n[�*!�3�G,��?G�~��9���FU�Y��W�ӗ��.��y�_�-=�h�Ը��};�}�f!���kYT��=_�Z�OXZ� �y\���U��c�����������^Wm��a������El�#r��%�{e}Y��瘂��a����Q�f�VzVa�l�Ac��� ��e%�G���c��������O{XR�!�A�kQ��A�,��+��2W�#�eI���ʁ6hb:�n�'�kA�f�{�~2;	��@��%��x�?�>��=�K\��B�b�읩�A=H˜�CSW�oYϊ�8�s��Um�#��Щq��E������n'o��E�(M��'ֵ�
=F4�[�Nȏx��V�"�+�*�9�;+���G\4d�������d�<��t�v�F�^9�P�HVD*�����)��[�u*��ȇ�~��G�d~*��V�~��4�NERA�t��v
�;�(r![��y������|=�=�f!tO��6�T;?f��7W�q� �t��Q��mi��A�����5m�F�\����-�&�*�~i(`��%Ջ�16a�6HE�ݬ^��y|78��Tr�1��)��d��%Nz�i|��
��R���y����`|�i��}��4�R�!��w�9�I��O���RnG��r���l3���G=-9ּl$�>�E)>��Ȣ�L/Lz�x,�� +��s?��R�y�6W���ԛ��@_�
G@�6�´݊�"����cj�f���P�H8�c�AD �Е���5Jm�Ph�B��P�R)�j������h�'��=h�QC��)�oubiw�x��[&�֓?(�F1��W��1��Nn�q��ϧ�_)rq�>��	�!a�����C�y2�8��f.�Z�E����؟���i�;�EB!T�UHU�Q��q�e��"-�車��������}F��r�¨NA3UY��4%ƤĺQ����j���x�Z����b�2�i��p՗��̩Ȝ0b#ť�]�|H�l�@zkc���I�,����OŋG��9�?���˸���}[i�#}���y	����*[n͟v��G�����K���CL*���<?R���GC4{ ������y�|%�$#�$60�`n�,��OD����������u	tC(��`J�:�A�M��-ߡ8y�.��T�	L�F֛Z����[r.QLG|V_����+� =fb,fL����N�[l%S~/V��cO���[�7ӌ:+��G�G�5ɴ��Y;���Vl�=>�s��N�Wg�Y�ȗdF2ɿ�ҋ�6�n��r�oF��fL>:��Z�}�˯Iu�/��F�H��`����r>�3NGM�Tv��y�6{�>���)����������Ұ\!�|�e�1�)r.|��%�@�Ս��DuZ�G����V4�)�v�\F�Y��8�qԗ�oy<ep[D������SKA���w*�����ƞt�m�o���mzz�mV���Ns�am��V;K���t���ԛ�?3r����P6�V�ڜ��-I��;�C)�	��a4��q�����QKJ���kwA�_���U�\S���q���o�m�﫥��w*:������],��/W�tM={�I�1�,-L/���-��]&iR<�fq�O��7�E��C����M+S������{My+Wd�Zt��xS����쉌@���r��o8�)���8�Lu�sE1X� X,���X���d�(n@K�9ݞ;�{ZO�X|�6pc����x%/霄�Qě�Nܟ�)T���))"1�t�מ�䢝��"������T�M���ż4*h%{q*x�A�3$X8R%Xڕ��:�����I�h�?�l��l����̱c�,s��9p<p��#4B;*p�5I����/wU�ob�"�I�O��P�����K��O-�ԷD���bS�
N���[D.ɱ`vh��^mq�{��iWe�,� ����ES�ZT��GPU=��[�uK����Y����!�^g#���N���KnPOfh��㞋I�t�3`ޢ	1�W�a�^U���~B���`��Uʴpޚ���,��>����ᯪ�؎��8iԁ�ng6�d�Ő����h��'Ǫ����uF�!t�n�1����L��x�b�D�=C�� ���r4���a߾ �9� �Yx��(��P�F�L^Ѻ����O�[R�lRK��iA�^f�#��Ǝ�� ��߿����H��᠕k����)at��؆�	��[�E��'��cs�I�8���U�E5�Цc���cp�����I�2�������X���x�9���⸍,+�����0X䂹��F�>�d��Xձ�R���l��aR��T��H�������4�??t�"��a�)����)'�{�]|�'E�	~�S�VK��q �v����B/z��]�Ֆ85�W�\�`_��kl��p(���|)�B�m,��;�搟A��[U2�W�
h��������h�졷ZbG�邆WzD�*_(,V"���O���K��n��'�����f�������P��5���w�P��5o+'�&�3��9+��w�2 ��'؈��O��)�W_w�95T�U�sA74��?�L�~��ʧ�Ǿ�_R��}Ƶ	7E��ܢ"i��#E�׿�i�H�'�)!��7�@eol��nu�b$[!P�M�D���l?�F;�`uZ�^$�#�q��!����r���j@P6,p�h5��$wץ�"*�,�y��ȤB���y^��c/�q���S�������FG��f��Id�h��y�q�d9�X���[x>���4��S��pGb�T�ii��x=�P*��[��Qh�_$0�#����_�Y�]���(��&/p�����>R���(<����bFS�Өe��^7}8�6Ͻ.����w��d����U"h�>���8�1VKƦSn7W--��p��D-n�B�D���Ю�L�,vk�ŎπE�@�2~��ɍ�t~��kp�%r���+���(�=�y�ƖHB��{OS䀅�W(��2�~����|m;5 ���l�J047��;_ �z�7	�-��@�PtI�{I�ψ-��sO<�������� `�H�X�[�	������x�9�!r�n�UҼ�l*����[b`&FKJ� ���$��{�]�j_�(H&�0�,X�P�$���O6FV�j{���a�~%/P,��ܴ��IPAEe��70z
��v���ƵN�Z�l2�.���{�'�	��қ��#�<g3
����}���w��86ۑ?��Lӟ�|g�!�\�����6A��n;ۓ�Xl�c`��h��6U�a�^F]"~چHByX�K֩��������s��(� ��4f���c��Ps�R)���/��g�t1�	,����{l���Rbe/�c�>rx����S�q70�M�'W��w'���� �*ɗ6�����:�X��V�>!��c���U���A��棠|W=�83�Ô���Ҵ�f/1:-�c�Iޑ�l�{��l�W�J�kk�	��e���}�b׌o����̶��kL,گe��Cjd�p+�n;�٩��=��+ueP �ʦڥR3::�?\�23�8B���V��|J���t��ugzyj�:�3�1�-T�f�}XCWJ���97�D�U�!5�zE���z��)���M(����Թ�qv��[�lO=&����g�kB�O��([?�c����ψ�M1y^�c062R�$��p�M���PZ3�v@߼w�nv�l}"x���o��A��z�-Tׅ�][�1��ە����#�"�q�ܠ���XJ ��n�������p�����[����H�w6$���qh���fkX���~��k�`��<�0�ٹ�����@QJh�K����?�w�~�/��h�M9*�p��Ĳ���М~vE�~����秬<%0�-N��*�T�Y����"�-YM*��
�#�ٵ�{��l�3��,`h�=��tM�W�uж�U\cQ�!{u����ȳh����(�%EJ~&�|7�׀�=iv��;��+�5�;����ƒo/Bd�x��g���DZ4���f� ~�TU�¬�ټ�h�z���A��s� ���ǧ�'��Q���4����cJ��L�b�_9B��K&�\!�p�~1
N���J8�n�|-@Y	�E��&�X��o������*F�����2ꓛ��M܆�Y��ݽ��;t�����4��,�&��b:>�����l<*_UĐ��,��o�1Ŭ�tx�6��ʬ	'����{�+�d�?�u4�&�O�?���T�y�	n�
��򝵌�N3�	��8!����~2�-Fafi�rX�HE@Ud�D-�G�{�ϧ�uk	wZ_�xB��n3�o�¶,[�h���CI|�bw�,�`D˶
&��t�3�,1�O��h}`q�"���~*G�R�esg5��ׂ��w�s�R�RF��f���Rb<.HG��;.9`Yo�M�S�����j�E*��T&<�!k��³�a�ވ~�T�2�����ed
Ԫ)�pi��V�s���8Q����R���^��!�»�s��n��1JP~�#�azX*t������} �& IP�y�n��4����4��R;vRf��4�5�����S��y0!J@�,�ۏ��-R��W��ׅ���<d���s�1�+=�Ų�b9_���!�R�1^���)�ʤl�L��G�7�;\|���K�fA���&����\l��.ݘ�W 9�$�Vc���O�B
�]�
�y1O������X�A@��wMS�^H��Ė���~*��1?���ZpC��I���[�[ޓ��xQ��ws�n��S�^t�����Co�]E�-�T���`�E���5�m¼��
��v�?~�[�L�ZQ���/FS�-Ftb��ה �� M@�	O.O���PZ�ڧϜ�o��#���~W����@�-p�a�)���noS��<�j����z�ŵ���.�-��"����֦`3X1�*�'b�Ƀ��<��~|mAC���L�C?���_A�Lx3!�����ɀ��A�Tw�KҴ�����Ͱ�uѝ�hB�:i2/W��Z㴼'�Xi����`��7�DԻ��;z P�Jp���ӪF�� 0�1�,�jCr��K�U��_��l/���=NG�g#
��ݒ��M��{�wуw|�9����4�<kcA6�F���g7����r��C��H�����(h�k����+�Z˦����"}��� ��Қ0:;&>dש��� oG�<O�-����jI=�3��*j��r΅�̿������"*��1��<N���Ku`d�������=�i\�DqFR��H�_�Η-�#iO3j���TР:K@b��&�}�T��X,��1�5�}��[����+��:}:���;��-_�����-=,��H���g�u庐�W:�f �W��m�8p�䇅�6B~�]�4�a��Bhjx���qx�t�!D^y�@"D�/�����r�!F�Ή�h9[M�Rn߶�D�H�&��U��e��.�jUK#m���}�<�>�� �����"���t���c��Q�[�*���{q��^��ԬUr�Y�J�k>�t�f#����V�)��xo���ܮ^����<��3�
�mim�h�,��	P���"��M��Q��i�`��j�Hi��!�4xX�]�\J��>e�wŖ�&�3Mi�4N���;ib�����WN��$���M� ��.�m���� v�9�S=z���ޖ�̱��_����|V�8�k�<+N�&/��r���*X�i�~~�>D����?�l]�HY�>���F&	�#�KxK�Sh73���d�J����^���M+���^�W��I�w6~t*�*�{���d�\lݞ��,x���?�2^fKP���R܄b�ul���FŲe��cJ��"[b\��5U�Q�(�󡬴��+�	<�~���F�L�<q���M1���ι���N(�N�~�ks܅�`�J���'�܃�+��W|�<�q�7�}O,`�$��r�J�l*��+��~���8�,$Ѹ��֚ls��Q���s>�w�N�����(���)閟��^<��Ҳ���oE�*L����p��쀕�*�S�3_�c���E"l��l�H0��߇O�a��s�<��$�"柋����L�Z��wh'/���z����d��J��?�W٢,Y�T�i����2�L��)��V�b��Nv�������R�.a����8�.���^�F�M$�Õ��¸�O��t�2����RR=Q��W`0J�n��>�v�;��v꼢	y�Ѩ2dL=�y�d/� 	PS�_�+��<r�YHW���:P��>�K��#�7Q��d����ZI��Xc�j�{wC �-Z�IU\5z��j�lܪ�]�}!R�Mjf熤��sV}��4�^�p�Qݞ�W���j';!�W�c��bcm���DT���l���t�*�/[�%z�l�H�C-�+�S�]�5:n�y��v���N*�s5�p,߄�[b�C>N����̣��'Hj�Yr�u���F�l =l>��H�`.�R\Ҏ��C�A��(���as�������<C�����R5:�K�Hi�=%5���RK���4Yuif*al�d��[�Ҿ\O�b��~��6�;�BEM���]��{<`�]9,G('o{���tT�\�ٛ;�vI��4
߭��-��}^d��1_�똘w����j/M��?�
G���i(���qS���ʺ�����f��XKv�ޘƊP��m����
�ز�*:~6UOtA�P%���,��KE�
o{Ϟm�)��oc��b�b�2�
������Fݛ���|��aNͭF����Z�t�:�;aqaE�ȘK}o��(5SG�x�!�G@����2S�ga!�&�?p�� �N���>/�):K��0��*�:Xd
�9
;}02��Z�M�EJ3�.��eT�_�vM�pi|�p�.��'kUAIO�ZR�|�p@�*�;�-���ҹ���]ŪQ�%)��U���{j&��z�0���*�v�y������ER]��D��>��"B闗��$[���[q���Ư%����O���-�˻uK��a+��ju�9l� ���o$]p!�\�rc����Fv�b��ejs3�>V<
��A�7��v�CY����|7��aȌ��fK�mH��D-qc������R�6T5���`�e�_�અ� ��"���E�Z��	��i~��7�L%�>�7X�}ʨ(��ɀ�"f����*���@�EM�Y�+�	��_�l�]��R�ħA�/

��w&�<T��81��#�Ƌ�|x�'�FM�&��|rЫ͋&C��f�(���]�\���Vh"tw��}��H�D������oH�K��Ϩ$-�C�d��9WYD�N'EW~�O@j̲y�7��g|�#��Jb���~ȗh�������w������� f�U��u�*��n�U���E�8���+�&�Y^��<׳O�4�^Y���h�LG�A�S�N�w��ʋ�"�{Z�q��8T��Z���yK^(�^d;
�×4#u�K����_�"�uO�������^�I�x0� �+��������9�d&f�HR�k>ed�9���˝��-�m�P����f��)�q����m��x�.�4�6)&��u�"��3�3�Ｇ0E��c��(� �<,+��/(������o?�����N	�6(>��v��ag�{��ޕ]?�`e'�鬗T��?8�dAv�)g���-+W�~�I�ֆ�喖܌N��vQhz�p�^f�^ks	������9�h��i{���)P�
�xOT��T���;cذ, @��y�s_��ڐƵj�56�n�K����	n��=ܨf CL���=!�7;-m=i��;�vc��9�����J�)܍��*~"��2��4�I`�������v�u��[�)f�wW�'��e�9�=�U�@�Hl�rx�u�Ĝ �a$v�5��,��Oنb�e�moO��ez{��uX�{���(V������{Ք��~5���h?6��m�l]�g�B�\Y|��!����[�oAC�g�٣�����	ǇkҠi�*y�ys�^��?��)D;�+� �.�e�U��l�c��s0�V�B��L��m��K���F�P^�U~|ۙ1��'�Ė��8JV��ů�/v2��tc�����=���E!�����|�Kd��p�h��S��p|�OZ�d��s��<y	_E��MV�\͠��m���?�����۳�&_�JM����[	VDOr�"���M���fc2Ɉ)�����^g�~���ַ�U���&����]lFD�y��T\�D�R��j�_O��2�^��xǗY��5@x�d< h��N�)4/:X�6N��+��I��g��N�j�㽢�g���o�,�D:�Y�z"B=0�92fS dxX��mlV/�h|�ev~p؏T�u4�WdM��طvYO���Q�L���T��~$�|����Y/l4{g�FhFX�GL��!�RfD��Te����#�{�$[��N���\�$6XG0��<���b�0AF;R���]N�0�JN"�p��cT43�7@DY��|Q]���G�\�":�M�y����N3�	�p�m]#,k�4��J�O��XB������~�W;~,�UԀR�Z�f�R�\���Ă��P�\UG�(<NJAY�BGb^Δ���C[i,i9DF���j�K1�h޺K��O�D��r�v�+�f���*��O�4T)�PC��{��iFu����r��|��/ �&��0�� {+tݞ�*��H�������a���9�R��֧M��i�k�	.F�K�J�oY�/]��I�z�7���1��0
sٹ��]G�$J��}�]	Gk�Ī��0�,YrH^�`!�}c�>4���g:֒}J��-n��Ζ�))c�k[^qS��S .FZ�T~P���g�
�1�cVҬ�b�rE���M�Y�����f~�.��v?�":�V�h=c��42P�ݳ�{c����Dj[���}����jrV��P���@����j�������ސ�ȷ<2hS��,�6��X����;gU�8�(�}9���};��!�s^`�M5��Q�*�w��~��j�TgM���0z1�����"�$ww�Kҽ V�?<DEl6^��N�Ǽ��)�+"�	]cV �#��.������u	��%�m9dL�U�F�/�!�^�&�8+F\�c���Z3|�e�9��k���s�����%�kwNw�vY��0����7p|������ty�}�o��^sXRdOه�~�@���BN�]�@a�E����N���-���^�:��i�s��ۇ������]E�!-���}1脾�}��f���q��t��o�!�[�c�N���d�z5®6ws.��]p��l=���u���� ��RJ�)z�Ziu9���ޢ]x}���3B@. �S�V���\�p:��8���0'!�;qI�V�P ^$!��ȼ'f%%�M����'��%0�]�������몼n)|�-�y��r{q<����$�z�A�y��&��o<i����u��~O��;�-�^���Q^�	�݅,L����p�����H�G�{h0��Q-��&J�?eQ%�Hd�XG�F���Z:CCQL['ښ.��6#��a7ː���1V>,W+v� {�0�� �o]�B�䏜0=�1&}UU�-�:�����x~�H݌�z~�iN���D���R�ݎ\�nLn����r���DO��Τ��� �D��a[��\<x���ʠ��&�@��g�}0���g�	IID�ե���H���ܡ���cj���D��D��)v�2	
;���� ����M�,���D��K�U���K�'�/te����o���J����b���>�~q������|������eźG�O�S��E[�]7��l�]������S�6�4o=1nP ���lB�Uc�ЮV���hN�?�r�!�^��1�L�훽�Ӵ�<AXU�o�zV��aV�v]��I�4�_�T�+7$�]��s�������u���T��RN��/\#�c� ��?��yb٭�iA32P�����=�a�E��������m͟�hMC�����h��<o%�C�z�2|^O�:�u
^C��l�7����~6v�Q��y��)����2�*>ŽW���IPP������Gb����]@�~>�#��
��WB�z,�#%Ok���a��P�d�r��8t��ڟX��\3���G]�?,HO�%P������3��a6/��k�m��m0�VN�yŐw1��jO���C)��@Ӛ>�&�fxL�������Ɋ�Ty�@�D7t�Js|�Cf[��D�v)��ˆ���-�![�Ϟ�,�,���rc�u�F�|)<����$y��;���!f*Ep �c����<��.y3c�<�u�9��O��Qʸ�xf!���u v��֦�%G��}j�`���tt*3J�HBqnr4�6|�����7ՃT�+��SF�������	�@�x�m��	�T�0	l�|�Y�q���/B��������Tr�J3N���D�U�MFl�X9&�X�&������6-+�iz�����������y��ǱXU�f���~���I�ds��/;��ۡƝc_sUX��gˤ�T�e�_���#k��C}�^i<i��th��2�l�Fp�;�1e7�4����e�5�ec3�� ���*e�9��둦^�L���w�/����`�wf<��s؍}7Y\6,�M�Y�x�Z���-�5���3�f[ �'���"��fVW��n���}�!������@
m?mC��j�%��}�@ԝ����!��
M%���Gv��H���n\90�#��k�����w�����
�}�TB�((�X�Ug>�;(�Nf���\�Q�$�QfzY�[����:3O��6��BvV�E�V�>W���М�������L�
x���K�c'�/�H�O��JX@x?���x�5\��y�S����Je�i�`|PYA<kI��a��3��/t�R�i���C3Ǝ�����V&��Ps�+6���������E��h��W`�M���7ݙ��L%��7J+�8��7oc؅�m���X7�JH"ts�-��i�ނC��Z,���4�~`&���㩍M&MYD�:�!��rj7}�H�O��W�z��bG��H��������y�\��)��w��r4ֺ��)��=�A��"q|j�Kt;�do����Ӏ��zȣ5uerSH���W�>Fv�e���vf"�����,%�,֜�SI�P��O��T�8g�����Y��ʹ�C��64�}-?���^:�[�!-��q��WM3�T�(y���+�y�J�(�H�.l��h�!3,�R͠|x&�&���O e�r�W���2S�l�NC��I�rS�p�S�p\t��?N�پ8C]�hLA�����-B�O�eQb��Im�B�����:��Y�u�V'^��Vk��=>{��L�'������R@�FBM�M��y��bV�˪ �WAE��<A�A�4�D���[j�A��"�#@-Q���k~�e4���z&]7W�	�7�9�xV_�m���I�6ޔ����A_�����Z���]F�ŻB���ƁGb9��HpG����;YzCv�?Q������*�t�	�z��O1�=}�<ao���(`�rhù�-�
eʙ��#,�t���O�c�ޙF�M�'�
h�Ù����	=g��O�����7�a�۹D蓼m��d��;'�x]�☕Z�&ׁ�lc�\Sp.{e���aN�uͭ{���D�ʰ�bݐv�J�I�.r�DaNX@Nb���~����[�؏���<�>��-BF���h)<E.2�B���^o�emzq��(�K}Z�be'��3��F���)h��xP|D$����_,�%@6O�A�o��ܼr��t5/�b3*�9�aŏ�P�2���ii	����Q�������ꁓ8�X���Zֆ�d1<J;F�Nł5Į_��sJ�0f�D�,r��SO&���6��OZ�U���b����,�V�R�{I�$�I�796���(8�����0+�P{8pׯԊw\��&�+�'%#�/r��y���W����Gg�p7�%���NM������8�K�u��8�D�_�E�h�#E��X]N�cd��B�E��A�O��D/6P\�d�\B	�g�����Z���t(�HN5�X|@2�QE�o�$���(���M�[_�|W��<8�e_*.����'"sn:0~�K��?����/P�討?q����l[3q���q`���� !7D�`:�-,�!�����*�!����,}�3š����_gl����Z?���w�̂� O����בscdI+�UC����;w�� Q�\��d�(��٫A-QCJ�ϝ�`��C�(��(4���eU#�G;�j'�b(�Tϰ�w�Ѵ�I���=��H�Cђ�	��O�\\�N�	�+�Y_����[*]Q��W����u����&8�eœ���R��ʤ��V�� �J�\Kq���E+���~�:`���B[�m��.��uf�M_��E�G�����ӊ�)KƠ�<��6����c�#]`�����v!��̈́.�(�AO�I|�����ܵC���uw�?h b�o�V����l8��c��7%��?e>�S$KNA���K:���x5�E��A�>b��v��br�ر?蚍9���)5r"�+o.nn|��Ɏg�.zJ."��=1�*m�y��l�o&(^Ou:c��^o�Dk$Y�����1g!I�}�}Xs�hՌ�"�BN ��p}ms�R�8�A��G�8��/y(<@]|�V&.Z���~
D&(��
����N'����#y�1��,wm�M�㾲��Vm�;��d�M��}}�O��φ�W�^rN-U�/�z�8���k��e���A�I�~R.
��:U�.택!0D�B���*N��w��ÉU2��" �IU�@J<�(��&ʻ�G&��� !�n(Z8+8�-h��F�ܘd¦���0�-��;Ćr"��7ԯ��5�|�[��,���O4�K��<�F��x��r}ft_z@� �FH��ԉ$e��57l���ֻˈ�D�݌	��� �3���D_�;7V��~�BE�V4DF�~���X��b��H���yv��vB�FqZ��S�Mb7�r-�3�K��Z� Q���r��;rP���[�HR�m�1#}iU��O�F,�z����hܐ���ܗ�h������?��&�����j�7����z����B��g��R%�	����T�e�=��"F_���H�7��L09����Aذ+d��]�F�
7nip����M�t��j%�[�-���% +Е-'X���)*�*����'��幺v�:8���)|ӵ�Zʠ��!���;�!�����.ɽ��m��+�nӬ���~7r��W̷�����J�����^�:�WN|j��A0ƛZ���
H���H�}�8�'qH#��w�AwbL� c�wtXT��=�#
�4��B��n$��%kS
ߠ���O�ȗy������]��l��{k�)c)����l3x�g`,{��l�9e.k����L�<�� =(	�5�y��G �p�f͹�K���#8���,�R�����7�����}�?��a���R��4+`�v
	:.����݃N
�NIF횝��Z�\f�b��q�:�����'���B���!t${iTf#���w2�N��q%��-r��;d0��o+T~yRy�����,��1�؟��&����h���o�]���5˗���ҎYO(m<6�#�G��"��z������ҝ-e`��w/7ĈZş�Zr�1|�"��/KjWOs��e�T�*���t�{hU��)���GZk�U%"9?�AE��"�l�{ז�O�-t��#�t&|��H#p��P��y�I)��d���bSkw��j�X	�h,�aҋ�cPmK���?�Kn���(���X��+! �;ѳ%q��T�2G$w��)r\� �B3"f�>�Bp���Ջ7@E�:YS�[xs����H����F�;�X�KL�d>��XE���\;���,Ҳ4_��������*c� /�
���#�9��$ˇ-�OsJU����S^V�V��0��ҞQv��$ N��В�\�ɥg�6���`��5]_��XW�h���GU�����9�\�MF�i*]�DM�D�B�_�����R�����Kh���^Q����V�����T�r����u�r�L��7:�X��,��E���s�a�b������t�iI�^��R.��餏U�r!�z8��Q�R5�R/�E�"hz�څ��z�_��T��o�8�G�I��CVz���	��c���by�nH߼�����#�,�yʝ�H�H���s1�Ǜ���zm������(��B
�c"�w>�r���j;���*=G���o�&�~e��!�m�q�:�?,ƥ���M)�Y��z!kp�1b�=K�.��#� �9vo^��̱(G�K)�J8��8�M�20�]:j9�����m1���M���%�W��*��"���Ȇ�ʐe���+�ql
5�Ck'
3}��zb����aw����ߵ�����`���n���$�/��L���v�����Y�d��τ���n��/3d�1�`�͝��[fg̝��������b���i��G�����%�{��]���:�����a�>�y⎳z�l�ɺ�չ`����bv�
Dmo������,5��Q��E*�@�cĳBsG30a��)��l׿n��Z� 6�t�3:��R捔�����|%׀�7�jO�`G��0B��>O�s{?e(̙��#�r��F��ZW��D��$�}U�ؕ��L"���w�8��o��*�s.�����YAI+��:�F��F�8�s�kA��/i/������Mm&����+��5�=�x��N��xl�"��:o1>|���b�x�
*��"/��ԣ߳`���}�S��##�Kb��ʻF�����]Ȣ{�}�+B���� 9!�����o�zÓ�q��@��\o%9DV~K{����T!Vx.�j��~�u
�?W�jH��k��qĉͺI����{�1}1��W$�02P�7�v��p$y�+qv��"Rp��?�q�R��l ^���0oR��eK���d ���gS{�׽�MG�����QS��������`;�8{���	��D)��ȭ\����}2i��(�ܯ����P7�ee��tɟ�kA����'�5ڐh';�Mci�����g_�Tݬ�{�Q�x��4 \"E�Ǟ`xb�l�U�s$sU��.�w~�
r��!l���F��Y��6��F�F���{��=��̔GGe�Yy�S3Y�H&ҳ�9N��1- ��~Y��Ⱥ):e�(�u'�w6E߰jqKo�k� X-.��\��#:���"�׷5��L���[�"��b�st�l�����N 6Dr��G��z���,}s4��
��M��8���	�����F�]�����<a#��HĐ�a���[XT�q����Pw�iv����xr�W��@��	��d@� �1�&� ���!_�z#���z�p3Ԧ��4���E}]zqN��,���FI-3 ���NL^���A��+=��XS�����Xw��"�]�.��p��H!O����)�#����>���b�(��Re��_ː�ئ,L�ZP�U�)�h��c}���[%��۾�b�L�]�K�81���-�|cJZ��$�`���;��ժ�Jk�#���:���,�R~<��n��d�5�s���G��%0��Y@�E�u�k#���G	F4r�����\�����w�D]�\c ���(�[��Ig_�*�E��L�L^W�P�h_1�@�+bС�����>h��l�c~�#�(<�\a����^��X�N��"ajc��-{k��;`�7e��p�~G����˰"twpT�.=7g��}�C�䮈P�5�t�9�y����=�0�]��l¸�X* �E���F�U��fO�qg�=L!�Ӂ���t�2��B
O|�b���q��rG;PJ�tR,�#�sm&3X����`�F���
��:�ew�:�6���r�>��U�>'��=MBBZ���z�e�$���|Dg�󛑆�
܌�8KqI����kgI��r89L 	�_Kw�_C> KN�ٍY���֗�,{�yG�G0�J��v�5$���La�ֆK�47WWa���"�52[0�D�IXJ�&_q,�`_Ͻ�C���S�XЄ�2���V�C��u�B��\�N�E�إX#�E��&sG�e�s�hͣLt㑚W�H���S���e�Vd~�!�i�:G���Yʺ9y�9� ���AAc!��7Z�5��WM�­��fJKfSS��0~�'f����&���L�G�dľC3:j%$O�|���WSh.`:(�D@%��Mk���*F�����{1{C(�nS;n��60x��=F��+p�Q���z�ž|�a�&�E�u�>S�%B�/���ğþW��O(CT:��Z�+g��Af��m˘=͏́�8�C�8_��W�e�!\v���ǒT��6��ƴ�_y=G<�C�����υ}�E��a��S�:O�o�x����\[�#��9Y{gf8Ta4����%��7p˸���<���qS�'���\����`�ۻC�U��\��oE�Aѭv�'"�0�m�w/��d[��
�@�S]�7�+'�?�x0��p��D�Jjz�YtKx��o��ȷ����������q,P��j2l<p|gHPMn�����KXuʘ���~��M��f��J\���T��1��YǒwK[�X�M�f��ח�9 V#��$�s��N�G�i.>����8��~���z���Ho��؎1H�X�,��f!.�Zn�`�7���!�������
%�g����j5�YzSʁJ�̳΍w)F��HviL#f��ܵB�M9���n@��?����'I��r~�_Yn�UB�D�г�MD�@@@N�,ع���Ҫ*���?rR���:Y\�߷��r��^ַW�[d��=s7w��G�g��˚���O�p�ۭF% ��f�����CуE���f�{�'5,2�k��:O���R�'���$�Z�&�����Azu�Vr�q��f�>d�|�u�z�m
<�Mq֒�S"��:�� LK6Pu_f���%Bh����86��ln�3(�ԕBn1p�gIy�5�)�>��b�;ќ>�d�������2{N��޺�G-��#6GE󳴷#?�=Ӛ����cj��?`��e0aL�����Z�z�@���6,��%�9@��~�J�*.�f�f�����2�s�(t�D�\NA�3rK��tR.��tFa����Kw{WU��&��0��"��f�O4=+}x�NZ?��CG��y±��G���WX I�'�E�4��4"��!�q0����uW�'Κ��F��Ѡ��T�}�bzd��O�����Ͱ2��V�|0_�rl|�J=�L���ǕI�e{?]p�&��#���&0��r~��g��f��t�+ ��S ��7�
b����CSy�u�X����l�&�d1�x#Mcr��̅�^�_$��[)�#� ����\�<�`,_�{J�����B��@��7��v�*w�7��R���u�B�P�5��:3Q�wM�Ў��\	/��t���)0DҜm<x��I7a3R �l����p�m��qFH����l��?���R8��Nβ��������3^���{4�v#E�;�ϙ}�Ӧ@6��F��X�M[���I�ŗQcg�A�Z�U��堷
�td�α�ʃ8�w��1�A�We�~�U��+@ �\�~���ί1'ͼ<rB,�4v���	b��y��Ƣ[i} ���z�b>�Zؑc� �/�wKTʽ6r��cT�1�Թ��a�r��g�^�}�j��4�PP5?�:�"j��Dl����G�Z"���	P_W|-Кp��|����F�B��Fn�=6 O}ag]���,�;5�*��,"�#���YZ֭D�0�gB�(���'���A��je �+��9Ay�A��b0����2�1�8�-�ߔy,�PEM������j����®�3,&��m���Y�,ͣ�9Ŝɲ�����5F�m����ΓEHg1�;՘��tG���yI�-Ņ~I6oU��7V�h���ie"�*�xg��i�;�<_v�NH=��aR�T5������]W^�L�������:?߆*+{�sU7KY��T����W��!2FS���Mۙ�ƝN�1MK>Nk��.R���%u}_�C�M�g��E�6��[J=��`������acWQu1|$&>��GBg �R��v�^�Q�L�{9ul�24��C�t	�Ư^�mv4C�����2�+��,)Ce|�Tb�a`��2�^}8���Z��srI ����
10��r��8�A�͔(*uH�Ƿ)GLN��se� F�1D����⶗8]���u�U�E�m��)���2�#,���]<,x-�3����g��,G'�_�5�3����+~0��M{D�}��h��D|/M������U������+�0BB�6�k��kj.Z�����1��%�@6��=�n��R��I_�oLZk�R1'�>ZC*�/w��y�fXn�)��N���&D�ln�%%"���|�ZO�0�u�y�?Y���ĸ���ͦi��D����؏�O��1���I���!�:�{�*�3UCl��_Ԉd7������/�N���x� Wn�Kap��k���-�TԡEֲ�����21�z!뜆����t�M7��nc�ޘ7�x&ք���lq�c	����K}e� ����0���S�3?ejn�P��=�WZ͢��i�����a��4�k����	�8m���x5��j�b�g�JA;�����nW'��=J
�)�G�ɟ~���H�6x�F�jY���s��T�i����D)8mhH�\F��7WiGi��6o�Ь�b(H����x�Y֙�1���܍\�=6��Ak(�>�����,\�P��B�	�8~8��d8	������ݚ ���7�-�@zFP�O�զ�)�b�}��6�K�ʪ�2En|�r��~EQ,Ĩ�,�}��KE[6���&�n1́/ e��y�۪���^�U^�-��ă~)�N��Eg�4	=LTT3�]��^�~CAV��HYQӘo & K^j҃�U�*�KHb��q�,ε&Z��a@���D��Wn�*�[��4��������,X.��/F"9ȹl������T�/tT�"�������x�Q��R��P����V�'q9�j��I���_��������ٕ�4	�[��)"��qs/t7��yJ`����B����]�b�L���Dz�fȬ�e,�[�Na��'�iU�I�t�ȏ�/���eE����^��D%��Y1��N��o��~"#t}�Y�� O�Yp�����m�6}��%R���L0i�bq�L�J���D_`Ko��W3�n��K���CEr�\pn������f�Q��dս�|�r�昦��RF��X9TX���W��ƥ��-!����<�]���8�O���l��h�Z/f�������kB��V0Iֳ1g7�0�g����H2Ee���`N��ZЈH��c�&�Ҟz���F�W<g�c�V�ZSl�z����	���ih�I\>k�(��%�8�#>j��ze-�����2��m��JC�u�A{톶⿨z�Rb�Vۇ%�j�
e�n���1D��!.L�XM4Ƨ�2C���u�G�X��CXk4B� Wˈ`q�t+<����!	��N\�ת��=z�F��UK�=�-�{m��GtN�xn���+Nq�7���RӰW�C���E���|��f��E=�@(6��zN��9vh�H�zg.\�>�c��>Կ?����r�0�'�t�����Z�ɛC��v6-�ٮ�@�{0h��֔Y�ה��E��dV��#����uN� m�+]��P'}��οm N�,�30�t��F��������91FO.`PC�h��]��aV������������~�P��K ����-�K�/�ÖE���*�Z���wO�@1�e�,5@(�_���E���$GVi"=��zY.M��Mؼ^9�1,� ���'���Ti�YBS܁im�����DB�qh5�4������'�pB�Y�؜�Y+S+�����i�K"ŹC���[���}�S�u��'H�fW�$��Q�Ž�J���B9چ�6F��]�f�t��v�1��<F���T�!���e�jq�O�:���W��,�f�Y}���>Y�>]���3~�6���TWtT���9bi�,5R�M�Oic�%7٢�yk8��JgŇ^'f�[���P:��7�-T/i����)�0%b��r^�do�, &�%ڗ��ʯx�$��༺;˵�:�P����b���o{�[�f����ʲ��d�~��k�(e�x����Ҧ�����PhƋ�7s������!﹞��!�=�`���iQ_���*�	E���4B�BQOov��a* �TrD�l��+�wؗo-����X��N�ηʅ�@�����e���n��<��ր������t#q����u��t�w|��G�[�[enE8�EaV��Ͽ�%�G��H'�F���r��/�>��M��1�S/ԖZ�в~jI�i�N}~e�?��g��O{a��Kv� ���75f�D@R@�^�ۢ9ۦ�ue5�������N�o$��aQ�b�O�By�mг̸	$�@�@ЅO�B��(�J���w�.&g�%=��{!�CxTs��}�6��8�ZG�)��@�;�ł��U�'�-�7�g�~�����U��/���Ya dXj��m���[��ґس�hٓ��?+$��6�[\}���:Lx�*C�N�ܗ�w���hiE�;��2�>۔<�O.y��H1�F�f��z��Ս}OE#���a�lpp��k�V��
�d4Yw�f�"{����)vr(H�y���b�{$j'_�m���z����������Qh�qIhWN�D���w`��VUf��nW:����5��[=��j	�\�;D7�w�W}�8��p�x�L/�P��%�&�S��`�m=n�&<�f���3�[~����E��Ȧ}o$vY]��Q8)��=��-B�*��|ȡ��ԃ0\��g�� �wT�0MeI��P@�5�]ÿӉ��|S��z���	{vK�1����z.(Qj��<*���b3�z��7��G��;��x$R��u΃{z��.N!&���gz��ʻ���)Y�3����d��?d���n�R	�LӁ�?Ow���ޠ��,�Ȅ��,.�l�"q{���s�>_YjD#T}+?�|U�G�$�X+[����Mz�R�-�6�����CkG�L�w涯a������G�iB�A��"�E�:,�MM�(�1wIt0V�[_�>���Fa�vwAo��J?Ծ��=U�Z�Q``d�L��Ԃ_ �R϶�A�Ke&���@�"�z�:뼳@[����@��h_�\�e6Z�-��ղ$�뿟Je<~��M�����ſŎܽB�oW?sf��e$~}���2h*m�І�ъ[�����QT�E?�1��49{���u���:�r^ےbn�S�5�%;aj��T�qi�5�0�.�}^��	ހ�l�u��%&*�2�#�3�rW�ɊH��k����c�n����aV`����CS�
M�ђbuF������mǬ�J����� і���^QZ�L��'(A�$�8��*.���ikwF��j���l0�t�$�8�L�V=Y��lWJ<'����LD��uT��F=��S�丸�����SA����}x43i�O����-ua����_\�",����h���Oc�g��!��&(ò%ŉ>�GW�5A����I%o����v�+p�S`�L^.0V_G��'�F�$�}�S^������ǋ�~��n΄��smv5�敀!yx�G�$��Tz֖�ʿX�*�u`�!��! W��z�K�?x�1+�(�lXS? �����m\U����)U$��\Ϧ�k�@[(���r�K��/�
S]!�L.]]���4���;�@7����*�܇p��!��F���7�#0����)K7%�%�;�P��Dp���( r�3��֧;|�~���K.���C�1�#a�g���Rѭt�Gi�VD�9ۗ��o2��?�n�*+�$<�P�Y��Y�����4�se�����.��8A��l�,��I0�/��ECM�`y�]���X2֪n�4�w mѾ��i��^*���1Ee�,萯�]Xߙ��">���yt0�癍=��lҽ�=I@����q�@M[����#QpLu�f�+*��C���'c�����m���>[���&�9��l�q3T�M�U&�u�*6-�`�,�5
����^Ky=+��޶Oj���q�|a.����琾���$>�Wr��c���sllȱ*���~��:�2�M�nI����i����}��R?k��Z���,��'H�u+h��5N�l�`1s�u$�8��%R��5.L���������� �Qi�2bȄC.)Uzծ�������E�ŝ
yY�.;��6�&tzz�`Z��0c!J!�uv������g����}W��kc@����xan6/�D�C/���>���)u@ϾӸ�BA��.�U!K���	۔X��0�;��+��yt�Вm�4����gw*���Z=�|̡f�hj����#"�V� ,���E���2�D/ ��sƉ˼��&?����T���Z����ݐ��r���L>V́��>���5�w�W�f4E�j�V�?ѧ��?Ė��)t��R��Y�����N�M �\�N5��-��s��J�1�i��F�V������XC=�#;\^
�-��}c�U�(��7���h=&���כi�Od���1$�^p���HN�y��12s���AR� tD�~�f�_\����=�  J��6+�+;<<���MC4�����g;[[�HnW6�<H�[�����a>M@ ��K҉X���������]��7Q���!���1��~��{a�2Z�^}������տf@����k�SW��@�-l�i��y+��)W)/<V�@UK���/�%Kԕ5�]}"��F�fj~}�4n�t��.��'9 �b7JG(��BHt�
N>��8�&W=�.�{��#���mlֱ�
��	S�L��������oN~^�y�<x���
�%��-�����·[H�3�Ǡ���p��I��A�~�*cMd�?$㉽�̹���|0�@C��=���ˌ�Lf#��>��s�T������U��T 6SJ?��t�������{:IEs��&�W]��8fp4jy��LC�~P�z�����($���Ɩ>�.��>�Xh�19�q�`#D�]ޱ3G��̭�p�)����T�/���Z���:dʫ�3�zM�4�\>��O���7�/ﲲ&���*d�u88
Fs�e�n�xL��7����Y?:��M�s�VQ� ی�F�Z7�<<B��������`�M���2l�`�G 1�~<�V�7�P�90y=R
��?��`���^l�>qN���o�.� !��'��Ö�Bj��n���i��t	�<�X��Y�I����f�Am�3]�=WZ��+���*��hyLɀ�eH���7�	 C���ȋ�×�7̪³�G���@���%� sOi�c��A�$�9�ʈ�����jvg��O
,���:�b�Ȉ�����9��,D��y��/,�5I_~�"4��Q�ǓE<�%<�.Q 9�ԶD`@6���9��Nz�-zo��G��t��2P��֭7��6<}�;:��ͅ؉REW���^m�Y>����������vA�FSן�rHf��zF��z���k�I�A�Ȁfɒ��j)�r,lʟ�~פ�`�1�yڥJ�6���`j�%Xc����`�7ly)-�ŕ�S�"��:2�0}�d$	Gz�>�d_���j�x�ُ����(��H����s�~�g��q#~y�?�?�)ҵN/&�
�/��������ӏ���f[�<�U~���=�}�,g�&��tP�o���;�{�um���nʃ�b~���Oɶ�8��_���a
�I��k�_��3]��yQg'�2ǌGOyQu0y���I��-=�r˺���m%���z��!P�����L�/h;����-�M'n��CO��Lw��ekk�X��m������YƌcM"���u�`�5ˮ�j����O4��5�=�(`U��|����h37�)�R��踨�4#��p䫜l~�FPw�6�y/i�8�.S�7�W�b)�RY� is�<���~��'�3`?>:;X�{Y7�HQ�!�Eg���݃�;ĕ�u�����(��A�2mMg�u�9^24��ijc��K�Ϫ���N�<��e:@1���e��"8pY��#ߙ2��'���S�ڗ��m����I�bȲcҩ���5�H���8������}:Q����"y�52�� ��di���j7��A��z/
��k���og��� $��2�[k�K(d^B9��A՟���7��:���~���?��\��a}��Ee�hj^*�{jY�UL=AC�W��d�̲M�"�$�����_]q�/db 1��c�3
ؗ��nWX {��R�t;�j+W��ki��1CG�I���ʻ
7�L�j�qtg��������B�"��j.�^iFuF� t��Ch�k�ZW�sK�9�[�g��;Wȴ�)h[�|)�� ��d@�?���"ܻ��/6֙ҋԭ��aZ!��0_��IJ��dޮ��y����]��-���d�������r�v��y�~�]+��L�n�Ci�l�M�=�X� ɕb�rƾ)�[�Z+>�ƇK�K
�ݺ�����fi��v%a\�Ag�&�ES�gG�EK�@:��w����r0�jy�TЅ�C[sa�ӷ+�������5��P��6�%��"����u��X�%db�)G?�m�kP*3�V@��U�=�^na���m�@�nĳ����@���h F�%�:SKb���Q�������g��m|,�����X2ܧ'�wK�@�WZ�(S|����t�����`㪑��%�n�`����:}�Yƈ�@E<��c��!˞�T��wo|'	yN
u�(�A�;iU��}����¼o��Z;�n4�u�Td��4W��aI����Z�� �F��O��"b�dt
�=�m�t	����`ܤ"TC�WM�����8��}��F�}��k�o�n�zL��ܖ��6�X��n\��k�����S�;��D���y5��}�Ի��fX�>��8�	;��^Sσ�IBT &n�c�>)���&z!��JF\�:�Hr�!�dc�Y��QK4�#
�Z��s�Ϯ,7�шw����)*�;|�^K�z�v(�J��K�AB��3҇y��G�R��l��ѥ �m��p%�
G0�Q:����)EH>���9�W-<wzdotNR����}�����nebS�����R.#ի���`����[*�H��Q�k��FF��О��\�{4V(�eY�xL�2A��?>��j�@q�R��}9��g�����0l 	�I��G(l�{~'�Y-��1�C�?�[>�sAth���}W�^.͵T��0��U��HDmH���&�Wp�Y�WU#��+yZ]�hƼt�4\����Muz�ݪ���~�(Sg��G�Hz����9�<���h!ҍw�ػ[�����Q)�% v���1Q~清��jEq�a�\9�b��vwu}4Bs���P�R'�y�o�mC�	�W�#��1�X�y5Xۨ�٧8���~=,<�,��_�
y�@�D	_��Ƕ���� �BpP�2q��p:,���R��e�!�G���7�X�2΁E����[��N��pKkTT: k7ݑ�Μ���!h{�rg�F���H��8k����R����f�>�� )�.�FzO!2��3�X<�������%#5$��)4{�$��2+��$*&�t>���U��ɞb�j\ED�ӑ�
%���~�R"3�d�i��՟��NqcN���Թ��"��ݮޜ�1�N���+�3~wB5]y������?Y�q��f��Ӂ�k����}p�JcK�m�0�N\l%w[�%R�1��|9]�e�0��ϕ�*U���N̖dy��B�d�;u��/\�����Q��J���o�+r�W��}���,R��g1o����p��I�9%,I�`�/�*28F)��z j��4�'����c�2:����S���.b�7W;n&�,f7��Z�>�{��q3�c��x,KƂK�#M������7<}��-Y���n�����i�1��h��K�9������sz�+�C��;�@��Zm�c$�&��K�d)x�Uv��}8"�}H�t�?߶��Iv��.r����G'�:�q.�`qf�,Z���_䜨�H�!��{}j����]��;$����:ؼ�3?��9�z:t	��{�;�ZM�i>�#���V;U�5qDy�SaW�s�}�7�a��(	x-�l$����C�`e$v�+�b j\_��|���׍	lI�*�ɫ�����p�;T�tʏ����t]�� +܍/K<�b�y����/���M��.T�V�i��B�ڔ�ãO��#���в�_�����MQZ�i�Gʞ�e�k�*�y, Z"��]VN��)j�
c��3���JӠ/�:���K@\$���gCϞ&I�7�#t�