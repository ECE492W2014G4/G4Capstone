��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�"��F9s�`&���a�oq���F�g�O�]�<ݲ����eCL��D���{�5��8̝DFI��Zp\m|Q��
�}�6C���UnF:<�jΈ�2�����<����sf�k��,jڙ�����2��X��Ss�HL��	�������+g?���N�Ż�����|�v7�{M��VNB
��Rs�゙�Ld\��X�'��R :�J���^�����kMkx�Q���3!P}�e���Z�Y?.�U{�RP	�)��lI{tI(S
7ZF�I��!X3�f#d��l�%����ڱR��v.:������S/��3ob����H�?�Jb�<
��%�Н��:b`�,}� Ҁ�j���1�����Qa�F��hL
��VLd��a��>|�x�[��A9���loN�}c%�o���8[,ѯ�*>�L������������3�g~@�-<�#�鱓�j�7rl��*R$0���z^�X>��˧�K`ï�6O<q[n�!sz`Ømi`��x��4L����*�Q��_���$���
��Ő����2bhr�C5�ArXr��.)�]ź����tqV_b0
l�۟;������$�b�d�<���7��-��I5�����i����@d�� �)a��in �"��]]��q�=���x�w-��@~�+ޓ�Ly	M��>�n��JȺ֫�n�����>�8B+ws ��L��5�_��ԝ�f.h�g��+eޫ"�,K���a%�F��9� ��ɫ�
�_��i�)���<�
E�c�eU�j�=�b#���Y��ȶ:[  ��w�s��ގޑb��c����Eg����M�HU@ �v�v��E6�:|W;J��Oh������X�s����+�7C7�2��"i%IB�IAR�<�u��_gܻl��D/tr`����e��dY�l�+���'��4�0jd����M���T֔伓�~�~6��ީ5�Gb��^���V���O�"fTpU���e��n��P�Ұ�(�ɨR��*@\ɣJέ<�9��� �Џ��®2z��55)l�e-"���3u&�F����/ڧ����5g�
���n\�:��6y8̓��$���A�Q�Jr:���{s�CHa�t��[�e���h�tzȰv�[�]W��)�YC-����b���M�;�2�ȷP���_���p�\H�i�h���+��I�+�_���O�	@��8	[��3��;�gH6u��r�����DR�$��<�O̽��4ϓ�pC��Uv�:)�G���=t���$���C�Ά2���/�W4ʨ9&4�~���e0{Z�/�
�WX���8�G�N�'�sd���:�ċH�zö*-��v!�R[BH0�R[�:��
Q��D���r2�	�@����uL`���7<�E�4��:l���dƳaB��CB�D�nu�]#V;��|�-,pß�{�'Z�^�����q,K n��� �y#�|B�-=�ݟ8�`$uh&FF�)�l�՗5޴d�\+&
��.1��d��X����� �T�9�{ܠ��7l�/噞�x�U�n˔�Q�� ڕ0D�xu7��CK��������G��q5��A��y��S�Ʈ����%�q,l~�(�l���.9�3���#}ac��3J�����2n�j��*�I���#�q4>w	�:��k�lЅ|mw5�吸� ڑc�J07\��Ho�Ǭl��ѣ0�u�\K~����!�X_O�z��K>�NT�]3+����ʎ�:�m��,=�)U����Ც�./��s��DC[�63�}&���O����O�تG�S,�c%�>6��o_���x6-R�[��^���¢ǜA���TW�^ꉌ-��!~��Z����LT:�)B�	f���lz���C�����tmK];|�m@_|��2��k�Ӻ⤅�5-D&I����G�֌`���ަjп/,q����r'�F �<ئ�479ksև��o�yD�)�.�Z)�u��V�.*gf �Ppw��}�/��6�J��7���,��'�@]\O^�S�9�A���ʉ�t֫ʟi`u�\��1�!�tB&�9s,�<3Y���ϛTp`+�)rP�y�D���[Fե �\�3.�[����:#�ƻ%P�t�s�$z��-%��ρ���l�������,�<6�8󇰶�����/�.�iW����K=�L��5���y e��|��������"W���u����A��/�J���A�λ}��s���I��9D4��}���"9���{�m���zN�{`b�kk/�t��9�
<��"�	~��o�;�"�I}�Z-M��?�����s���6Ŀ��F� ����L�ö�A�m���xJ�{�sRM�	;|
[�Q{͵D�����@HX1Q��T�����cvq����Y��U9f4����c��Ɋ1�]s(Q�6%�<�$�ܲ0Z��*���A�w�C2z"���ǳ�=��&.�Y6��ݢ�]BH��H�@ϡ6�nLH��N�������ҲI&�8��V3�#�~��2D���:h5�,��ӧ��"��iRy���KZ����,�&Ш,3*r�bz�3O�o�185��B9�Ϩ���ݠ%�fa�]���mυ�d{yo7ϼv1P4L����t��U��.��=D?�����~k������D�����ۥ�v:Sy�XE�����J76*�2�A����}�w3�G���%T�!���z�E�ѴA��@���&l�	���W�+[E_x��4lb�Z*�AL�E��t�	]�.Y����f�zZ���]�I!��/o�2pp�w���� [��R߶B�bf��2^'��qe{�)� �e��Q�V��/#!�R��%n�������4��0&N�W��F��� �ߚ�6Y*d�p���Lr�>��|g+�r�Ik�:�N��*�J{^5�����H!6��svq�]��D^�������ڦ<$;$��\r#O+�^���ۦI��X�.y_�@��ʲ�������}q��H���ENk�7/n��	
�b�!IsLQ��l�[U���&�
��������<,4�gJ�h3>DGO��=�Y�y��u�Fb���S�
H�I�VY�<]�odγi�Ȝ:��B&�~Fa��(-�N���x�5sB>i��29��uw�HM58g��Q�Dt�FE\���ʈ��))BX�7Y�����3h|(���3�c�:C�q|*��mZ����0ju�k�*�z0�$��KB���'c�1@1A#��fY�B�X
��L�}v��ez´꿒��ڄ�:��hʒr[� ʪ*˲J���p�P��/�B(�lLTvr�S8Zi��D5�;���u��j�reB@wH80��[3�Z��L����>�|a�F����W�DD8���3q
�������f}�/��ܗ<�40s��%f��j�rT �W��|������;$ R���xA�����8���E7���J�Җ���;�&%]���"!"���4�bMVm��k�ʬ�Y���H<No�͌h������~��L]�U�Ĉ�+�?8Ȇ���4lG9�J��5�Ϫ�c!p�%oV"������������ծ����Q'0�``ߟ��������jP�G�����:�����g-d��3	ڸz	�߱(��8�V�7�:
�	K��c���#J�{3��ke��Ci��������{^��ɾg��dZx��G����"�F�jy5k��{���
�Z�9jR�J�{��)���.?�"��Ӊ�I�
�	j�8�x�o�n�%�|��ό���:!�̭�a��X�Hza>��_��M�iC7�j�����w5=�)&a�լrba��v&��W���W�7�>�;#ݲ��M���n.8!@�#ȉ#�Z��L��ܐy�oս9��޳ ���I�2�f�|��Y�O����1�>�wAmPop]�F�����~&�( --����hqE��F��u�x��sֶ��$sR*�!������.�s7��Jo)�
��K����4�����2/��-Ag��j�E�%��A��z���P�	���0�0[ɭ񔿉���O['�0�������&0xP1;�?�cs�*���MN5��j�}��>��1�h�sR�L$��c`Dʧ+'��e�!@��0�uA��H[8�	^���3k^��g�s��Ԑ�b?����qv���6k���[o����xGy�%;������W��N6�T�+��=A/�#J����X"X��Y�Z��!L���υ�SO�?�Y�*�T]�7�X�q�6[|u��&�� �E����RQ��h�j3w5!�*�s@A���'U���י����쮴�b�|G�(�Q�9�a���죞�b�Z��؄d�7!��<��Y�=�z�7�tW���!f�}q�Gd�{���"I=���/r+�no�\*���/�).wK�tʬb7�?��-;�/��n�8@V�wg t��I��G�7&�>�����7 �)�$K��ۋ��Q>-o�@���P&0�q����e��˵����hn���5�k��</�F����]���ru�B�3�*���렯K�����V�z���=�>��B�҈�_�z�,����.i�ֈ1��O>������BAKSԐZi�p
{q/���5@�9Jq<@q����]7*����~�8�O&�_&�l�s\*$��	�/H#t�b��u��0�����s�zQ��<e���
�*�#OsV�EE;�@&��
�^
b�b��{�o:���y��Sx�W��MXP��X��"yN�Dn��BS�|�VQB�w�l�|S���[��fi�w�/V3�͚*s��qXО�wGGs�0q��1����;p��F3}*�/%E�͇0�w��������� � ZS�~Ǫ�W3@��Ϭ�,a*5�n.gX=ݏ���$���n��f�V������!Ҋ^��Û�>�s���cL�����t��L�]�B�f<���x��l�$��OM<�)���-P~�9��z;�4a�����,p�gz�cǶ���߼�N�4D�����6���9zI��ԥ��qS�P��h���7S\[�C�oM0
t��[EwBluA�3Ja�|[Z�B�@7�qC
����a���BU���c����*k��(B��W픐\"Ja�,��Y9�>�X�.ˎ�M���Ne^���:��s�������J���?<��j�G �T��U�˚���ʊ���E�+�\۝:2ml{Μ�Ů����D-��3��!��¤TV�`���@��xB�.Z�>A�5*g�7���q�D��L��%���P �������A�<R�4����|�5��&J-2�B��r�b�L�@W>γ��`�D,�s�SE���3��J­�����g[��ubk�\�BR�}�z\T.I`�4��a-]=�Ҹi��[rKYL�\�ɞ,%����E&"�*	����\��8R�����M��J�ti5�7�z=�H��j���a�w��C@瑏E<��~b�3��B���?��@Y�u�Q����h���X����l&��9Y��i�c����D)�"
���?�J�!���Gxr�����������O �[�K�7�)�V���О2�E�10���Q�!�Q�W����tm���L`�j�#�j�zj'�z�q����{!��}R�?ر�|���������tռ�4��|�i?�*���(�gq��E��!�2�(`�v�%�Qa��V���y���aw=.��C����|>�,w'_ar��X3����/�=���l��G��̩��m=�����\=f!���H��o���X<.Y��I�q�Y��w��ʍ�J�y�J�&3B ��җ?מ��gX9�Wl�sZ�&o�Lf������ić��a���Ք2��<]�7�~���4��Ր�p-7&�q�%��\z�Us�]ch��;HQ�[s��1�ܡ�uy�L��P�&�75�o�~���]�2�ܷE�j/���](;��<@�_s�.q�Զ��H��H�4a�X����10��5:F�S�e�&���gJ��)��5��<�$�=��7ObsY��߾(�2�#m��}�Ȍ��q'd��S��U��.ի�����θov襏���F֮����	&��Rq�4Qf?ˎ:�{�hf�3���"�������B��/�'+��;�rMn#P�Q�u���� ���X>J����~�(h�Y>�պ�?�2�k{����jp��k��͟]�je���JI���#�9�W��A�q^�K�˩	U\	�<^T���	��9�X
��C������pmC��=�|d܆Qm��ث�0����ҁd�����4�Ұ��`�ӂ��2?�ܴ�����pbA+��d�n	D�C?au9�����	=P~�E�K���Sڍk���2��[I@q�_�r��M[c�ᓫ���T.w�fK��Pp���$��Y�O����c�ɽ���d�����2����/����A��Uw�*�T�ވ�<1��^��?�5xk����q��i���MA��t7&�x���n��H�V���dW��-ނd�jC+�����}�R�����M@�g��~����B��h���:�^��Wᾋh6:���ZV����	AI>�"�+���v�GY�TE+j湗q�յ�&��良��%~�B���������X�?h��5��T���FE�%�l��s>&$d�Q�����
�:��WEW3n�1����7��9I�Є����I�ӑ��.q)A%_�Z����EO�=�ǫ�O=�N�F
!��aV��7�OJ�<uaR�NA����9�0�K"u5Zo��x;m��	Y�͏��O�����[��Z��)��R¸y��w��e><t��]߳*�r�?_�@cjٰC$ 
�;����G��'T���-�/��#�=�u���8VJ�[M���^%���:b��$���U/�U�I�%+4�:�{���û��'�hd�w���CTæ�������y���@��Fq��&�U2Jg�(�s�N���
�3.}��OY"�'���c`s�3'9:�E��?<H��L2/�fT= -�ƽzl���y	pO�S�.T6�1������'r��&�~�����#�hGEy�4I �!����0��p��
���;	B=�j��i��ͅ�|���X�� �� H��U��"�)Q�Zw�{"� )��x)
d��\�r�M��!�u�|��N�n�0L��{x�<tsT���>(a=r^	�N"J�i���Hu��� i��(!i[paG���&�j��`u��V� ��`�f�D��Ħ���m� /<h��i脎 c�׳	���8�*Q��)��ň݅f<��8�!�����i�c@�ϔx~$wA��Ţ����``�Pq���J������U44�I�K{Q�й�hL7�lj���s��od��L���ؚ}Z�xw�va������G�k���'w�r�:x���EHJ8w;gzW���zc*�Բ�E8E(2��`9g[��?�K�
g[�/F�����g��LDv�����8��^#��\|��GW�hD�J-�������X���R�=�W#6Rc"0F�����y�� �1�9��tj;X�Ѧ��F�� V2-�S�tP�Z����]�7��?�>l�}����/n�zN#�?�5y��1 ;��C�%#TH����J�/�|��Ip4�M�/��n�> ��1��F�ܯ��k[��X٪���T���������>�(���ɹ���W�[�Bp6av����N��,?�z�Z��1G+���{T��Tc����:�q��y�N@�.�.���Y���@9%xM�A��b�����F%dș'G��a��y3+�����P��~7�w}�jt����)u�ɋ�Ӓ�-dj]��C�N���A'3ޱhcx��HO.(�a�:>pJ�(���	&���b{��喪����c�j�EQ��9����ц��'ﾆbu� b	*�W�5
(�4OU�c�I����y�{�wHk�a���$
�ki�-��	�V����SΘ@�B8��~z��\!�j��W�NIe���9H&��v��.+GgUT�G
�Q�o�%(+�om�yj�t+,���
�S�6Q���4��,*�g�#����2V?��EJx�zo����S�C<s��~����r"�̭��$*$��q����7�M��'�*�"4������@fWD���}k���s5F�i4gN��zpT��7�oa�ܩ���5/�w��V�xjr'�ƀÌ	W%WY3�	�f�|�!�����Q'9	��uogs �nhb�v<�NJ�tm�����Gu����
��	��Pj���?(U*{}�L��T.P��x����!k���>�o�cRF/��uE3���|{yD������D�Jp�![�(�h��)W��>x�r/���76pࠇ�+���c�`h�ď%z�������Z�>I��R�-�����B>�q
p��.c�J6���o��;
@m@mҲK�˦iUt���D�Y�v^�0|�fZ�^�d�blM�M��\����뷚�\�WI,��6S�\yq���> ��j��|���L#N*�(�ԛ[�z���d�9�HG�+��7Z#��ZۦO4�9AUkw��>>��n��(�0�zh�c��Y6'���<�GV=�I�~T�ƽ��>�Wg1�_ƍ��O��0�H}��&������i����7�F��v�ר�[���a��1&���K�n����$k<�6���c=�͋b"yQ�&�Q	��e �*Z��S�^�������iUA5�+Ku��̷��ļlGA���Z�y+zC��{�_u_(���b1XNzKb��mKng"D���sv� �"M*�i�rPֳ��g�pG�ɉ���`��o�Do�;��-y�J�~�F4U`}�<f�HX|�Ő��[�f`V}���(+\P�cpN��o���0��@��=m$��da�֤͔�g�[)�_`/��Ze�����������l�>Q�-�)vtv:C�+R��T&	��>|G	aǷbSr\���!��;g}������I�jI��B>Q}棁)��o���-Y�T�_�"�?�=��zm��(,�"�m�f�آ���%��}�Ue �����-�����"���3�/%�^;��;~p�21��I�y$M�m�`ݎ�F
ᷙ\y�0�������~T�kA�O� ���s�zю��j�4ML��� �~�g�8��W���/��a&:oU�3�L�k���T%��Y�ěxk���E���k�פV�7H^+t{�%�7�ȭ�P壩���"�1��֌�o,�;��� �G�����X����@O�2�;b�^~Qx=�7$c���7О*V�w�4��N�++J9���}���=��8Trb��q��j"���T���~���>p�7��Shl����zM��`��X/��f;��%x�ZO+j����f�Q]��3�+�1��p��KwJ(1�^%i�s���k�ߑl��<D��4�}����7�!�b�� ��������xĉmO�����te�n�rؕ ��H#��Q�\�W$�A"B�ݬQ/�F�1�>DL����ݠ^Ic�y�?���'�����~2�E���o��(��f����J��4�p2��2<��,� ӎ#s��٫F ���E����a����;��Vnh��I�Is�w	�����:���"�� ���t���FK3��&kG(��A�q�����Ղz?+�B�;U���Z|0�5.�m|�H���0q�dD F0���3x-��ix����(��DY�9Q�	s��$���n$�^����d�6��Lt�)iM!>�>�p��^k��_�HCK����4�x�Œ��B�-%��8�ǖ�MI�o����wa�XJ�~$�v�6��X����hW���Bl���KΊ,�Q9��z�6��N	4�h�!Ƴ�U� 3�a>�N��t������Q�_W��`8OXc-��A`��ՋG�.���D�bm���_i��~����;OϠ�V��5q1�)�ݞ�T��ƶ�����A�(��C�"tc�,)떏�#%b}�2~О��7�Y���=T\E��8�}�Nqm�ԩ>�|��U;D ���9kR3�����ըゥ.�+�/�|���,�f7Xӆ����<���.>�[�+����Zh_��گ*�6{K�4e@e�W�s����y%�.e��������t��<�fmY�kZ: ��I�����4 ��]f�fӀ��"��
C���2e��7�ު��I\3�� ����n_ Ղ�⿌%�*���6�z��Ӏ���@��Y1�$�߁��!��ozamh\�p�@�,��m�v!���d�(		�E'v�Zeηl<�LJ&~��J��flA�g�����O��}��+*
%��}�~�kr;�s�Zem���]���ˈF5��+kJ���2Zz�w�mf�;��� Hl=䲆'"�&���Y���8b�!?vv�t��KX�*mx������L�㺞hc���',*�ʹ)O�O��v �p�R���
T4�{t�믙���Yh%:��DN^%�8Ӕt���3�5g�a�;�L�;G��-����^�|��r0�RiUuY�]��{�=M�^5J޵>>���\��M�vPN$���I'�4��.�q�m�9�b���7�bF��̩���j$	- �G�Ĺ<\�}�j�ߪl�$�~4n�n�U!6�}��x�?hD�.�9C=��A0�L t�
]���(&m9�33���T�6X�����n���[��M�q�?��T�g��\U�w[X��0�!�Q\��hP�aG��z���FQżVdMr�!NBR��6C��a.�7��b7c��k3��yŔ�n1�]���O��y8�HˠKѩ����b+%>;�!+���,i{I����>�TB�=�<:�����<_�d��w��`:��Q�<���I����˷�pR4�|�������5O�Ο��jxM�r����FF��}o~���	:�8���=�z��2#���O�h�����I0��H�h����)@-���Y�繘ii����`6���6���^C�6��&�+o�C`��P���0І�I���,� �ݦ�T����g�˟Y����r��2�r�˥�@�t#�~��y�,uO�|$2�M�&������[��I��R�1F���� �#q�]��&Y��頧��~������g��_���X&��}�l��x���S������Uʊ��mH�W��2z��R��M���:�w=k�xÉ�6lO�]x-2lHqиfэ�o�� ���&�R��G�[?�]�0�G�h�LۏZk�ǣ����� �{S__G�mV�R-H���B�-� ��[0h�7���'��	I���'����$u�"��@�s�H�a>P��*E��\}S���o赗�����r�ڀv�����rD�p?H�9��`��C,���S+���J�����u����B~A;�K�0�7`�B��ð��ʇ/�r�Sƀ�ǇY����b>*'-J÷��D����o2oͦ!�@c�{!m�K3j�U=H�V�u	�����,�~ۍqݯh@J�f�K���7j%{.0�Vr�	"�C�E���Q��[i1 ~M&P+>b��E��ݚZ�&]�Ӈ�p5
�[J��#+��ˌ������W�����%1����
Ս��O��&����*�U�� q�T�ō���`�Tp�L~���~+��+P8�AI��kt�J#���< �&�T�����/ʡ���$�K|S��Ut��0����h$�#��)��⽔��ʔ�:�=�IwF|2�玡R���w<��vC�����D�TM.��s��|��Z����'�FM�Y��ΔD����Y|d�Z���|����
�l�ϰC�b�kM�9�\�����L���K9B��}=�~���Qc#5H(ccL��5��Yp�؂�
dri�B9U���5�G,#�k�w�$f�yTneiS=dך[Lo�n���'�N��9�8b��uF��a���|Fp�`>u��l<�p�`NuʻTv�ی�&��F���$������￬xlRR�O&����MƱc;������,�*��3���z�Ҋ��m�����+�}�\�F)DBE���3㕧�}�d�&t�=[tf1�d��A��0Ǖ�� <�����jx�@�X�R�w��W��ns��t�r�H>����`	�pW-2;���P���jg���9@�,6l3�9���>���R\��+��*qV��|U[�G8D$>��JU�_�~�ĂHN�%^��2(m�)�Ytb���^M��s�������'ϛ��W�U��r�6ĸ�~�g{���� ?o�aK���r�+"���5��d{���y�<��uml`H
��j5g���4�P��9�������*��n��ݴ!}7d��X�����M0�LQ��у nz�.p�������;�"�ķ
јS��,|k�@�T�����+;��>l�է��#6����O�Ub1�I%�K�6-[��`y�ֿ�R~�ļ#�og�SC���p8��8w��U��s^-��{r��:�X{m���5����pS�9���;�/��Xq��� ��3w�lTx�F'�>g��,�]`4�)|~�u�DP|�mB8tG����jJ�u�(���"J���
Z�Ўy�t����ߕC�d��h*P?�b4��6��d�y ��:<��&!�G���P�6�0�~��E�T��ݢ�b�o-'��+V�����[�+IA��pH��YklFНr��%��-��F�@1h�֎.bb��PԊ�֎o���nn��o�q����ϧ*�b����vm��6��9�	���?��!���
^��,�����E�瑿F��<F;�ʣ��g/�yYe4MxߦG�s�^3/
z̹�X���L���|�o��b����cb���)�)E�f,r�;T����n:�}K��еo�c·�@y�ʒ��ȉ�ڱѸ1聵��/�b!`������g"���ba�i��ΚW{LXўį�i�s}3��%݇��<yX��#�I-J��D��s��fË���r�z�MЅ�;��XC<��	��Ȳo5��H���^N�R Eݪ��d�~͏��R�~��V��鎱��p]�K	 UF����wփ��͆�5r�<$}NRKQ$�]�FL�uވU'��u]nd,��~K`�?伍jj���N2��x'�*�b����u;���O$�pc?���j���|�Wˍ�T��+�iQ�a�����(;�O��K����I�����u���6��<�t36��z��"g��uL�l2��b�D��Ǳ�ꙷM�l����6�1�l��QF1��y08�ه�@*� �dYpd�L�� ��7=z]��D%a*�<Y픍�(j�_�M�����(�6���a�-�9"{&�	�/�� S7�!���/(w�-9ʔ���	���r�H��P:�"�Dq`�� k����tB���rm�pw=��Co>r�+u���G�SϬG\����<<�\�s<ZɄ�Դ��z���Bd�.񥸡�7�r�k�߀{ғ���
��t�,�>�v���vc�Lw�+=�/0��c\sOiT�_w�ꅯ��Vf�nZ��Ѕ)`���.���n��G��[�.�s���Qh�al��(^LfN�e�?_��7���"߾�����O�Y��sƒ�$����"�A]��o)z!@��ҫЉz����ioе'�y�G��lm�\c��6������X�����h���&�6S�3����������|d���*`p�E"r�F*�h������Ijר�ŕ�+�Zfo���A��r�P�L�Ќ�!���!��;�O/�����2/��Hߖ�����⚮:U��/T��$8�e�6b!��h��v��\�e�J�?�E�$��˞=�Ұ	�%Y��u����@���v`y*;<^\3��IC?:��5���Z2BEQ�s��A�,!2�i$f�HJ���-$�	$�[����j�,Y��x�*�~���f�x���1C|�;��}��@ �h�V�z�PM�j/���0�}�Ȃ��~�I�8���\4���2�,�J���o�tp�9?���CFJ��ɠ�n�*Z��E	{�l���7��������rwdO���!E9��X�8&�୫�3�-�Lt����Qn�V�y�xȗ�eJ ��K�|�r�b�xD-"��)2�em4�_8|�^�H?���O��?]Ւ��ya47�BȢ�v; 8R	����P3I��H�z�_즗��\c>A��V�	�w��@3�:DZ�\��U�	G��+��8ȋ#QP�jc��*��cB�๤<in\���*TM��pb��>�4)�YkƬ�wޢ�B��Ƣ��p�!׹�~�G�'1����۱-%�G���i�r���7筁|���1���t7��)�~������_uT���<�:@xG'ɯ����h���{n�D��6�
!KC��Hal�4n�A.A��?#x���:�Lh4xWpR���0F�:���X$>������.U��xV��\CܳZ/�@�6�z���'F�-�����v��sF�{y_s�EAe�R��S��`���|�0�j�|f�:���j)2��˵����>��s��>I�\��HdN}깣ʨ��<�B��D~7��ɚ#��1���C��46��_��ǺF� ����S�P?�}�ψ��C8B&M1����t�6p�e��o��Z!t[���=�gWt�bHs>�	ӓ�ԧ�Z�"�z��ǐm�!~5������M`�f��xb����� �F[_'��=c�"	$�h8�~M=gy��1�dvt뿲d��%�\U�+J�E�'��攜�����[x����LpFe�r��W�G�ޛ9;����6ꋩk����-J1���?ڊ������*�u�ք"��K�|���.P֎&Oz)ܵeѶ� ���ɟ�r��;%o��K���M���-pw�;*�ya����+�����<�39�:se���������[�pQ<���b�����@֋|��s��t��?EZ�ș�'��T�U���%�~O�˥nN�R��A�_7�9B�z��2���{}�4�`ipf�|w�z�L�"�6���:�uL�u��wsdW%�����7z���B��\I�5�~�g�G�<������FT�їʙ@B�����8��Z�
�]`-�+�@A�2c'=Y�`��u�;���� �B7B��D.�Y*h�On�	cC~���8"-e�|�4�~���㬟�F{D��I�ݿ��=��RgWN �(��l��ݞ��O�q�-Y� s��]S���(���D���`��_=QY.��mQ{)o�� �D�?���'u�2LG$סo��w?����Q��r�w��w覀���w�I�I�m/�HbY]U��̇RC9��@�(������o� �@�e�ǌ7��ڊ����KZU|.��b�ne��A��@:��ʔ�xY?�k��bc��)E� `}�b�����"�p�i<9Rܓ�B�q�ub�Yf�o�?~�z#aHM��H~����?n"�ӭp�Hg8����`�	<�->u=��-0��(b�J{(�
��{��ᢿ�3�S�,�gO/G�|xD1�&\��v��d_�$�=v��I�v�6��ň�a�:��Cf�vɔ��(w�4��z�V�a��Ù�w��lh=��kv��`��!��J�UbR~�e*��Ș*"�M:��O� ��v����̬B�"�\jL�fFSt|��a�&�wk7lp7��}g��2��*Y�	� �e��)�B���h�7@�ѱ`g[�)���J$g���	n[҉5)w*D��(hR "2Bu�>~nX��G(�������$2~�2�N�'vg�P͌�ANE�pry�@VP�C���~���Ϟ�[Y�R�/����^�C�-�������͊Bʝt]V��y`)q5m=0k��y�l��d�¿����/�~�"i=Y�aC�kl�s�e5v�m��;��?ʉº��O�!S�mM�C8l��n��CO�O�����\}���%@uk'�v�`�7��mn�u ��N(��RPBr��<����b��!$���IsT_˾��Ԉ����RKHz�ۏ�Y	L�g!U��:�l�޲B:q5u�������'��l����8�쎣eR#��#�hK�N�6���uK]�s�?�Xڱ/W���pAZW���v�r�o���=Ӱփ>�:���P��f�����'
S��%1D�s�	#2u pr5Xk��7~��|hxEA��h5F0*q�Xi��,`���ji�:}�	�v.L�%h6Q�~MB��~��C�Dine�7�\�P
w����L�Mj~}>%7�<�N�Pm��w���J�u�� o�麒��I���&�U�K婑���z.%��Y6�K�{���x5-�u낉�0vX���n�q�����<�=��5"u�_l&�)�^l��	CU��9��9�3^.���
��L�C�8=~$!����\A��]�_����*�Gx����Κj�A�T�T��`�/V�uo��r��Y�3��R�?��jm4�̊���q���t������+�aP�T�&����.�遊b
@1Ю��qJqJ�X��,ژ�n�u�PN�=���ӄ��9�-4d?�j^'ҪXm�A�h<�c�l�$	���Z�e3�`|��b����|V<�O�ESA~����_�'K#��B�4Ś���ݺ�J�g��i��r;zZ;X�ӿ�hR{�o 6o<��M���}���`�i��M>JP�y�a(�@f<8��TQeta��޷�@���Y��y���M��aE
2�H�̀�.�"�.9�c�ؚ�fg.��#z��)hy}L�P��թV�B�������Ý����)�It6߻�����`�d��:1��\G:���,������������&�����wx%>(����uX���_1���i-5y��']�A�rI������
E��E�(
�m��1*H5À��O�m�!]v*�c�3Q�5�����r� Pev�>��0�)q����L�~&�c�Ip{N�,\ �f#[a�-9^�<��-���1�_�hM��f���Muc�w�b �NΞ@)�"����@�`��8i�������A��#�BÝ��"
V�h�C�������:��?�o�G�`�k(��tA% <p�ȡ��>@
��˶��Uy1gYo��!��g,����T�|S):GL��|��|\���$e����gʑ>>�4S���y���a��	�s6q��^T ��xsԲyv���4S�ё�]��$b42�(�5�b �̑j���}w�k�mA�J�zǸ��ā�6
��b�Q�t���޿5-�"&��B@�m�|�:����&�V�BQ�v�,>�p_B����u�+��3�ӫ��w�il�[q��[:�5$i�����a�&nO��.�:����[�����Ҍ��a#��_��+�"5���>}T�9���l���.�"+0�Ò�����0J��ZY��"��.8E�B�"��g;�G{���x���{�����1�����@��]t+��I�X�o��;55P���l-m�k�Х�su� �.�_.;|y��1�O7K�s-�*��˪�m�'�A�x�Z�i%SG�ʘ���54
�B�G��]y�籈mHk��UOכ�XI��n:�J�c��ۺ��;q �s��?��R����c��fC�u���Ad��z�@��q��#ZK+���Qv�V��`R����p�,�n[�:t���t����{����]u�Ȋ�8�/�$p�v��lT�`���LɫqOFJ[Q�5"�e[�Y��t�6#�!.���]�=�!���Ia�t��JQ���E,�v�a�>��0X0�Y�w��B�Kf�υ�RHd�4�P�~4�ڇS�S�͒'Lr+5W��-��9�E��s���o��ׄN�a�{��O�Z�#��+IIR'�7�B���?�~�B�T�`�π|Pw�����H��[х*��(���X�-���X��m�U`�=yǚ�pJ��Z��%�y�R��ψ�Ҝ�ؚ��/�6���X8�,�Dij�{?�Ȳ��ۂ�D��V�C�C��D1y�U(�:�aI=�G���&���}ꓢmB⁥�UL�{$�s�s�p��b�cQ�S�;��^�'�I�_u��>�_w�ō�r�	���$ɶ�0u���5�Ȧ�5�Y�a�z<!'�9:��
k�:y����^��x�&��4�N$ê-���\�WCn�}!�BaC[�Q���Á��c��ENED�c����;,\k�Pe��Q���f��Ge�n���a��g���@Q���=)�NNL�l&U31_F��ė-<�׊���ƫ����c3��m��$�ѯ3xX���f-���ր�-����Q��!�ub�0�8J��hZF̋���I8w��@d{FR������@!�1ٸ1��K��.�U��fN�@k)�c��ѹ���b��u�����9Ru]�3@�!ϱ	{����,���R���ÿr}�g-��E�Ƃ1� M�	�O��|��>��3b�i�5A,�b�p"�~�����6qz�ݻHǈ0�뷊9m���БZ�וI>��E�V��攆�G|�|RYp���X�����p4j4wߋ{<G�x�Is�+�C@�䤓4����	���˘�b�j��� ��XU���>Z�op�R�ӯW��>�ۂji�ڙ���|O�$bqX�n�pn��� �!�/��d�,�Nş2q�bC#�,�����i:�����O����R�7ƭ��M�xW)�	��q�� ��9���x<���y�5��#87Џ)4�	%X�W��҉~�T�.��M�'��=�2Ёl��~�����X�3n���a�ltW�	���������