��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|��We����kɄ�Dߒ����{����}w:/�$|�c|/^h�c�4A�|���<�r��}_�����SY���ʹUZK��;_��+��0�$0"�E�D%r6��2C+/S�o6�P�25�z+R���.��I<�%
W�,����\^���Fw���S�#�(>�m�u~�Uvwq�U=w�i"�H�W<�nޕ߃�#ǿY�����^jx���8��E���rFn퐵��b�9�ˑ��4�^p�n�e
0�_���F ��������R���NQcI�~:Nj���QY\g�k�G@�}��p��] �9�jLE�܈��%��^31D�!���,=�ðuǪ�2-ߘ���)�2��=��SQ�h��;��8�L&�"�]c�շ��,�]0��J=�H�b� �� ���)5�]u�R��ěI�̰F��:K�����a��@W�f��VD(5x����t��|�8 �+@���{1����:�-bfw�1OD$�Q����u��s�w��?�q����9�+�j2O�"p�Fw׌�����ji�ޮ#���Z:%q:���"W�U�>��fa�`���F���B�j��'�y��a���T^�Jh�T2-�O�i�6�B�_������5�a�a�)��Es�u�f�?t\���gl`��v���>��g��p�K_��"K[Z`}��j��W���O�6���V�J���[��?�
bQ�l�Fc�UJ��i�����\naIkj|U0����H�F�J��v?�v��(x�j���OH ܵ���U���;�.���62��$Y��',���[(���#��G�ym�bK����e����m+M��d/�=�a��7%uR�l
8�'�
�&Y.G8�8yH������ktV�LKĂ� ��ۘ��LԄ�����i���T���	����D��ρ�'������ҍ�bu�+ �t8Bb��ď��gpǨI�� w�Z}ё�\��I�����34��#�����Mì�g�v)�i���b�S��QE�5i�&.��� (�d�h�󇴨Lp�h�*�٪�m�,�$e�g�^�f�ڊ��2��A���ݘ�;fM��s�'c4T��Vm �7}�٨ӸA�^�I��G{~"�\7h��qų��yџ�=^|\��H�@C;v�sE����iN��ʪ��ţĩT�eu<adYW s�)��g��ʃ�6��+� ��tl���D�ʽ���|4�Y�>���IJz�
R�SE+b�^���_<��ܽ��k��Ч����_�p3:|�)-�R_���o-���+�(� ��0]�����m�s	�/&��R[9l���&�6�6R�l��#1\�����8�[��O�c�'�x7��Ts���%������;-Ȓ�tsyt��A����J���t�:L-�hp2��Eԛ^���8�)�{��1c>?h�ȖHPb�؈j~t˲b��7����o�V��_ʕ7����6�C������g3�%��`#���ڐ�N+vg!�_�*X�5]��4�8��9&�H�`�	���g6i�վ����m���o9���t>>}�^v���>1�����ŝ���1��2<��]����X{�m�H��h�0�w��c��nN�3�m0g����">�@���ʳ�l��?�|lcr�գ`���!�5ݤ6q�������#^�y��(*��2(�q�UQ�N�@����'�?@QxJ����'��L82�n]UXC�ܟ��nDQ�>����>\f�>�ON�ј	���_�YX���B��휃*JQ��s�����{��R�'���� ��#�jF�j��F��[Z �hrK��w��M�l��)��ܓ j�#]�.�9_�З#1K�QA�b0��T�q���K������}/'�m�w�4���v�+��0��$LL��E���23��ռ��=+�'��R��q�`�;]ڌ0��i?Rh����T�Ԛg���P��Z-�}�W!�)��j��D�e1��.G	���dVoޭ��V9ԑ�dZ�2�/!�F5���)�N��*6O����en�3��ۼ�9���3��J��z����T���y-s$̮�V٥� �9��C�H[��s�1�կ�5l���S7C�%J6�ԓ0��Ļ�bjb�0���z_@��9�s���g�ˮ�8�O����l9سӪW֓�8����������f���?g(F�P(HL��������m��ڙ[���A�E��?:�t�T�j�Km�ӂf�����c������Fc"�mЄC;�o�k�1��0�y���t���<�v2)��r��@~�z�W^�5רC�|Sd<��	j�5��{<1���,8}D�~糧��&N�s7�j�������_2��7ޤ��Țq��`�F���s�+՗;�l��ޙ��gɭ��D'|
蹕�{ml.�U�I8�u!;���dWj5Ӊ.����ˆ�p�q���a�����9	�jJ2�=��?"�]T;}ޜm]�;dٓёo�
09e+��d��Mn�J���k�/���V��E�{V�Y��>NMm�+V`-AL�=�B��T�aQ`~�ƞ��O���C4#)�a������	"����� 0�pj�[�D�c\>v�D��ن�Y_5(�Q�Yڜm졶8n�dL�W��}�.���d_&v��b�+1,=P}��\���^u��0[��7��k�L����E� �0�9Q�:(ևKYN�������&��y�U�|�7 ��.w1x����7�f=�4F�Uy�9�+gܲ��FD�F:iY�G�B�׺����r.C7UA������T��<�a�����HO��f�s�7�;_��j+
�q���G���^��oN�����
�G}~�"�H�l��:��hNRY��7��9;��#��J��,)����;
��'?�Z���X�L8�
��f�߼s�
15���v���
5kTn�bxlif9h\��Ɯ,Bh.�f���6���zl�����Y+����0̮�8�|	�V��U��/�@�&�,ۓr�]��x���������w����b�%H[��S��uZ�"�.���.�x�0����}���w/��x[2Z���&����p<-�e��k6��V���N���B<�����h�t)�*�J��d��G;�b��KD,���'�S�iK����$��7[�u��)�>�Զ$|�>�ǥ(���Xf�ݫ��_���6�����oy�$oS���.����%���6
���"���2u�J�^ب�
�և��c� ��<��n����sR2%$p ����c���߳	:�L���k# �����[�� �EH+{r��N�����%�R����|	'�}9�Z?���w������ox�+U�|���L�s�ړ��ǡ�J�bM���PC/�B�\��R �5n�k��l�S7e�c���;��G!�~^q1�M_<�_=XA�c�6,�?��e��0��FIC�Ҟ������5��A�A)q��O�M�:7���F	d�`���B��:C���Y���Vk��t�71G-O_�^M���m�[ ��o���$�+ b����$�nA�s�г�&y�ܶ�=�����5M�6�#rYtO7l]����[zK)ڕ�bGx�G-c������߸��4���w>�8CIx�sDE�:���<��,����GȎ;���Q��2QU�����\pS�O�d�v�A���s�'�~��e�7���Am/��c�i8��}o�Q��`���G�:
͟�JRQ��� e�F�9�1��,�KI(��([����х�,�%�p�X&p�:c.ϋ�*�0N�b�.��	_�kC�����S�m�f��k@G�h�m�l�,]]K���M�X;��T���t���@٪��6��y��}|QaƠU �� �'`)���C�8=��>`�ey*�w�'�K@>s��8o��@i��X(���_Asy���\o��؜ӫ���Pk�f��ro��|���
����1���.�g�<碟7Q�H�ڗ%���!^`�u �'��Owa��ш��&u��z+�rO���L�d�(���9�7��z/�;�>\������-�#S�uc!;����90�.��|��JC3�G%�����,��d��xȫ�A9���~�B���<�����S}#	)h�;�?L�s�5�y�)�2�.�kח�̈s��eX�6�q�~��?пd���逈�?�������a��oH?��)�S����6��T�����VJ���6����L��y]^F �5?�3��`��%hYn��i�'��!�����^�L�P{IDʿ�nx�n~��q��OO�.��/�	���511�{��ճ]�6����k������f�33U������Xd������l����"@t$rǽ��!x�GL}ɘ�ީ��{X�ӌc�Z�-��sw���a.Ɨ=�����刘��T�DDjZ}����>ﺦ��<�QA��\V0�|�I c	!�4ȐN{m���� ��?�[2�U4�dv�hY�m���j>�4KB3��<��;� &ub1C�vw�̰��S���7aѰ~�θ��09; �����״�p�d�&�ۡ�����F9�y��\�_���̺�ϝ���D��fw���k�5�&fot^�ȟ�=�)����689�IM�0��a�խ�:��ZV�cd2�9�;q��,:��WX֗�0��e�,���o��(N�*�S�N[^��������Q"1����>��f
y��~��Q�gySku�}(�����OK� ����*Pgª�?݄�#����	�q�}��[$��mƒ��H�u-k`��ق%@v�n�j.o�|�I)�hU�e(zO���)m'M���ڒE�J_�I�]jm$�S���hZs�f�x�A[��9Fʠ��n�O�]Ʀ<T����EB�-��`?��;T��]A �CR�t������@����!k�ȑ�
���/���ez��)�HSdV�8o�կ��H�.O�cE������-�`�F?Qޚܔ1 D��Pn)�LT���8��d)f��J8\2a��C�{�����p@�1�ɿ���k���6O��.�Ʉ�t�(G�<� qs�uػ���k��9��]Vr�&m� �u0=��:k�?Sr%�|~�<$C�x�}����_�d���B���j��A��@�~��HI�ɧ�a��y�k��|��?�����rՏi!Ӟ��8/��ѷ���ٓ�S��3rs-c�"��0}E�&��SΒB�Y��A%ۘ�&�.��9^6��T�>4�~��m 빇F�V�onB��p-�Q���.NWƹ��B~��׻� .-k�Zsf�O?}j�?��D#�����~s^�^M39Ҹg�$ �hЦ["�e�Y�6�����9��"�Y�د��j�v:��r�-���LL��󓒕c.��J�ؾ���ޚ��ɺB����juaG�Ze�J��l�qZ�.L\3�V�Wɿ��0���;1P�t�Ҕ����g�V��I�gR��bnyIAt4�5�~����칶���ET�����5h�����]��˸��u�_.��'�{ǪQ ?�x8՗��;�¢����	����]bi������F%�V|�5Y�jz%���,D#��A�������q�o��-Ƣ*�?���?f�1�%������$�L�=7<\�>�mV����p�l�w�%s���R��%t-�5o(��0�|�.��L�@�!� ��żM\�0���'(�.�y����&'*0��C���һ:ófΟ�#
T�-�L 0���i��i<�=�n�H)�b�a��=lpY�2�������.����.Q���6�8g���C��C������VlD�(��a*�<��<w�rL�ɒ�K7��a.��AYO��[��|0|��(�l�q��m�E��-�������l��+y+=Ĉ,
�%�%WX+7�P�T�Л�NC����}Wbw��"Ȫ�$��f�9rp����G�O�@
4)j9;m�)y:�����6���N�Z�/�$$�;�_�	-#��ㄩ(Y���i	��3n�6�9ͼ 7�5����A�r�2N�x�ITb�n�W:��I����ǚ��9���_���(,���sc��aU@�x�
�T�K9�}8�j�7Y\�դ`]��jQ��KJ�)��I�и��D� ��$���>������,��=$H�%J��_�:/�Q�q~Py�����R��4oH�KW�׺��z�zٓ� s��:
�h�0��`�@�)t����R��$���4%�?�-� �FB[�֔�(H�ʋ��莢q�l�HӜ12���D�϶��e1���WK��اZ��#����k��R��!t�!ʦ@q���ߓ�K�q)�#�gB¸����� �6�ӄ��ky��`�,������|#�+=����]�����)���]5Hp /����L�������G����2C���4�=;F�&wS�v�W<p#/�k��H����^�*½�7�f]�������M������˷�tcy֛Ot�|U�,?}�C��y��g�D�EQ��@H�M�=R=(�s�+�\��I�¬�C�y�5*�*�c��o8�"�3�[�`'�hI/�� Ő��J�&fݍh�d�+��7K>@�������~��:g�ȳ!]�]�+i�ٍ���&e�_�Cj��^\����-F?�I\ibm�/��'�C���g3%�Ӹ��@���P�s歨ͭp�v�U����v�04X��r��=���;Z	�R�C�&l��I&bڽ.�����>�����m���/�p�� 0p�'�=�D�1��E�I��%�e������U=�x2;H�>k��\���f�=�WAQ��D��Y>\���7���J��爕�e��#��jg��jw>����R��GQ��E�)�%����h�|�4���j���>�`���K�>2blu��j �Y�I4�~��%���Fq�&�G�lB��C�:fF���uq�W��j�:�"��8�<F~���I?.�'�Ytf����X���5*�W�ae@�\|ߕ�/�,,5<gW%���1�{�z^�5��Pŵ�6�����;�Y�52gL�(��ú����|I�����NY�\���8"8���*��߃KZ2B�m�	#X���yzD����%#Jb�T?�jG��q��?C?����c[;|-�NM�1B&��!��P��7�����Q���2EE�.1l�$�?Uh@GV#(��p�S�T�v��W9���%r��c���!�s���i�/;�dh17�\sԡ_��hVM��	���d9T��Ȅ���)ߞ�gκ�]m�S���SJ5�%@���.�׆9����얠�"$��@��@����@���dN?u����08|�fC��
��zYF�Q���q�2ޔN�JsL�`��ґ$'8�[:ᜲ�7�h. �J�w�[�ѻ��uX�%9�ځh%�M��?/���u�m}ط}��N���æP��B�z�S����ȲA�0��h�;��N3��iZ�$z�e�]�<d�=�����p�+�X�]��2�+/_+JG&��/�ws��W%�����O�Mw����� ���}~�σ����*�!g�$�y�q��.�4A�M�ώ*Waz䢙.Q���s�
_��ڢR��X���~�z�X|�b�<������2�� [��`a�	L�sD�,�<�U-C��TrOY����j��q�Q:N���-7Zp�x�0Z�2Z֊�&�41ɞ>^-oz����/ :M��W���(���Yk11&"ol��EX3��~�� �E�������_a����5(D}�0�ҁ�&���7g��x̲�a��%���_/�JgPG_�]�x)�Vr��C��*�-� �G��SH[H!f��m0/������I���?�^Z��_���_n��\�r��<�m����6��m� /`L��E�r���V7^�������"n�q��*M��5!���ܭ�o�E���Z���wCs�U$yUI�y����L�FH;Z��M�a�#��c;�+�jO:=�>߰�_��J�O��a߲�"!%��d�lI���f�V�����7������c4����*�A�SKCX����\�j�KL8���q�����]:�Oe�ϼ ���*�kN\�CN#ѫh��qa~���*�� �-�&5��nq��w�mL��C�$]��h���t�Q���k�I����b)/�g���C�#�}���֔cJ�wr迳H�aO*|���<���,�?p�GI�u�9m<�^�1�a˓���SbF}E�$rd8I�d6�oġ\�*�(}��W�J��bN��u��۶�pu\���N��oO�����ڰ�����jz��Z�p���j��ًoy��I�V0���:��s;f��$���=ȹ�=T�΄���W��˱�v��%�zl�։0��8��Kk�i���=�Xwgt�Y���[���VIhT�4������K���o���Dg9���K�_q����&�
��7�s��=OJ�@��X%���_V�����{Mo���J�Kp�h��K�&&#����:)Z�H�x�Pֻ���	� 	����S��2O��S���h�p���nQ�� ���|]�	�#a�g�ό���AͪX�s�=�u�����M���OM_w��H����S�9ۍ������=�>��{�K�ß*Ud���ͫ���0q��Q�\�sGV�����k��o�~j�	K�87�{2~M�
Ĺ�O�	K�f��q�y׮ǧ�~�!�=�l�i��B8�U���e�?P�����# +�f]H��͚������c��=�?P��`�<��B�����z���љ��Q�+bCl��X���_��>�����9���-B�%Z�R�� �F�9�fG��i�؃�ʿ~� ��hkՂ�9z�&=�������x�A$M���A�ă�Eg�Үc�^��-��L^v7�]��E����BX0�!�	|C`��L�2��nλ(�t��TU�F#.jEvqb��D:>O�y��#�%!R���S&��b�Kθ��S�!�"O5��p����y,V;J��:;_�[sWᕮ�~ubms���ِ�d���?�s2T�w��Og#/f��¯k��gQ��5G�mD`��Av�1���%�G���]N�ӶROAf?�2 ��Y���{�9^E���4D�(؉93�.��Qa�]������yD��EA�=�bc9�7Z�Ӆ�H8ɚQ��G ,)��=�ɰ:�;�"�ت��S�IJ�7qd\��6��Z��=y��u�㨽���m3p(f@6��+�<t������Ch�>�xT�M-oǿ�0=Uy�W���㕀Fɣ��	�5b�CC���~���,n��ʻQlW�k���qb���XC+ �Mf�K�D�`��}���8lS=W{!��r������7�L�8��&K�s�_�@��q��@m�6�:b�y'�AA��<s��tQ$c[?\�/���8O�@ʅ�
֦HS{,�K��A�y+-��L콽6� y�?�XR���I'���V�Ԉ�8��Ax �-����9��0�9t�������������+�"!�x���*��9���7`�������B��i+���=�}H�-�P��UliJm1AX�X��Ôe��I��!����Kb���ޞ-�����R�^,>A�ܩq��p����&8�Xg<�k�U�5p����
&��֖Lގ(�5��ı��߼8�o���Paڰ�̞W0p
B�S{�0�1˘�����@�>oE����.���z}��.�����u� �;p[�p����7Go��cBN$��mULݍ�x�I��/���q"�TT��p�z��v�`�(|�MW>�(�K���:g��=�=0��.b�x6��gj�>���os�|@2�Ur�V�4�Mz�؞9�"�"İ��ឧ�*�@J�y�.��zSS�ݲ�"XJ!3f85\���qJ�i�L0S���G�"�v�}T�
#�rHq��c_~��o>��qߍ\�(���~V�����0|��| ��a��F�o,^�4�Z~P��5�z�5�m;����0m.��I��KW����A�Ӫ��Y��#T��\�����)*�ɩi�6�Bo�{��n�@a��Y֣�2}�_�ݝ�&J���H���j�d�T��荌��Bb!�����oT��T������b�;�_8��z���%K]�up�H��͝˹@�S���z���#�
?�L����� ��ol���Q|�A� :����KU:����V�u�GZ=�I?�6���uڿ=���g�;�U�5����8 ����0��ɝ���M��;W7*�$ҧ�EkwR��1f�$��_o������<rZ����n�Ʀ,/�2�ge�y��
 �F�M�"�5i�8��r�]�L{o��?l�hp���Yq���4� k�QG��ǰ��3�DYS�7��(����Cˌ�e}������^|?J���]-����p����b��3 O�"��e�HE�ȘZiQ��>ܞ�RpIrt��<?>ɱ3�=խ�����ۅ�n���+8�Q�]��򦌴L֕y�U~�L��6P��/lk��KNb7�u���ݧ�kc�H6a+Ɖ�hF�����R��V�+�!�	���rU'^llX��:Z+r!
�/{dh�'�O�G�p\�̹s�/\τ��Χ�����Ԍ}	���j��˚���(;��h1����L�Ԫ�p��0W�n�O��A���<Q=&�3OVᔐ��J��nR ����)�� �QHꔇ���eB�h���
ҙ9c���eY�S�M�'u),R��@��4�'	����ŘCR�FOŁ�0��9S��T|�P�����,xpȏJ�- x��?`f��pG't)�ܴ�P��3��Nm9��tG\#n7[�4L�[g��(�[����H�G{y�_:�ؑ~<�jrP_ܳƃg��{�9b��=��Щ�bpW�i+G(�� M���6��{)�<����H������)�3��q~���/njh����.������r1IN9�ع^��S��9�5KF�n�y\�d�2*k��Y)zj��v&�d�U�O��