��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+���]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�O'�yz,�_ ���)ZN�6��dQr�p�x�y�C'�m��H.@'�!ѽ��Ќ����M�����9p��s���v���	a���y�A��n�M�1%�P��Jl���� �k�
:�q(T�F��l�F�j��;*Sc�e�op'Ho��$��'�*>��e���y������@�%X�9��o@����&RY/�~f�C��31�qĄ�J� ���2��:<��-��q*J�����>+e�!1��]4q§ �]m�ԫZ����v�����F�q�S��8�00�F�ړ� f
���O�Q�h� 1[o���zp[ �c�p �2q�:�W�9)�t�(�����1�B�ps�n�ri�s�R�ng~r�t.��:���\�d�@������P�R�;^��42��i�i�h���71���e�9��9��X���z�]-��a�g�g���w�4��i	�p��� g���؎m/�/�1��~�8V�;�$�5��V�xo%Di�%J��� rA��/h�}�	&�+��;��+�����hs.��,��ӌ�*�:6 9N'{������+�q���a��6�hszx�ݒ}�����_��9���*C��x���P��r�*�C���¶"�[fJ�c�.M� �3�ls	^�I�i~_G�X,쳳�V�U>h������.`e+/�|i��U��=��dF+n�I{V�Y�����azڬ���_�r��7�}P;�}{��+��,��AN��'avVhO����V}����[�����.�*���Q4�VB��q߻$�	��
V���y��35>~~��9Ƹmn"��)yA׵X���~�TO*�ad�m^�J��
O��f�o���sM��?��@��] (9έ���.�Fr���	6D/���e�L��Z���t�k�'�`xK4���ܛ3�/�d-Ny����Z#ŧ��:%�Z"�R���U���^4r?��4��Z
s�	Ȼ�#��x�O��F�-�⋀��a��\�S�����*���̨������j$��ʨ�)��i
Uݳ
k�i�?]'+��I��hk��� b��=�qy�Ok)���&>W�Q��ˇ�͑�/��es~�;%֫S� �f_�n~f?���Ӏ&\��bU~���Nܳ֏�N"+OS�,�Q���g�\���K��5��~����h���aT�l.�n4W�D����M�@��/-��kt�����lhFTp�dO0Jo�Бl���+#>0Ts'h�V���|e��H�Y	r* ���\QD<7�74�ǔ�ՏD���ֳ�=�-�zh{eg��$�S{v��|8�w3X��`&1,��Р]�&��+�y7]�E����X?E�"aQ�@d��X���FhAJ��j�I���fg��dAsQN�!ej�c��)&Y#j�&������v���@f��f�J�w�2��6�6t��'�g�n�����Kn���i�T��Jf��V��AW:�8��P?�djȐ���&��8��e�dY���/C��m��J���Ϡo^K��Va�U��(ⓖ�������ȉv��� �`�C��׬X8;�>��9#<xV��w
��O�k3�����7�+����Ax�s	á�ŏ�WJI�j�o�zQ/ت�u�3`i!���+>��>?H~�K�\/v* �^K��};0�U{��|�v�q�ږ��'0H�p�����[��d�� 鿢���R����3.1a�+�P���9S���~��T�-3i_x/{̾[�<
w�~����DNo�;��zU��S^L���g:���C+{�^��3u�94a@��)��C�^�<��K�]8�7Q��i�M�	p�2�N�6��U�[R�@�^p0��&!0��&�l~dZ�G�w-�G����]|Ѯ�؄����1Dc^A>d4s�#.M0f�8��c��;4��޺�V���� 6�G�S�+9ww7�xG#�E����`�yg�J��Sf����Lؚ՞��7�Fdp����N�4i�e�,�/]27�1�"Fq��p���K����C+�{����-��IR��9�O wu�x�^��/1�hTNIlkq�4⼁�Z����m�k�Ã�!�����������yDPz������x�*0-�H�ܑ��	�8J�9e�x.�А�ë���5�^� �9.�Y�����Z�΀�큇p�A����tG\�3�}�D���ȦrgJ{��	Z��mꈪ�� �ڏ�2��;z���v�_m����Xɤ��׈pc;�?m���D��]Q)�?�;p�yo��A�::�b`�ʍj@og���ݙ)�%�?��\�*@8��톬����d.$=,(��8�������ټ���������#���_DQ���7�>|X����ဨ&�?��W��ԧ�D�IU�p������-Ԇ<����ۨ�L\R٭/������#�� ��n��pq�o�3 1���_��Z��S�Q ����B���q��B���;q:������-v�#�i#����0:J���N�<;�S;h6d���Q8����Ӟ����ݘu��d˪��qy=�0i�Ň�D�Nhs<�=�j.?\��Cq�`��9����r# ^�G��>���a�׌��N��{F��+8�x�YB���JZ�7��|W�&��K>�丫S28t�Zd����ϭf��V��{�H;u�1�/sS���cT:��і��s*N�p���T�B�M#~��Bt�����ZJA�Y�n����|,1Tz4���4�z�uD��r�\wJ����Io\�(��)ێ��Ҙc�ҔR�g���i��.��b2�_�z���ְ���f�g����(֖4��߹�W�_���IZ�����V ���dc8 i����K<��W�ￓ-�������d�J�.h��q]�:��������Dɡ���������<�zF��m����F�؄b�t&��3 ��.À�+%���y(�&5������U���4���K����}�S�&mgdl
��=5O�UT#�|~�Ac8�gu�%�NOK����*� 0�1�T����j�*>;�����Y�Y���51p�([��ώ����i������2[�=Xi�K�w���̆��}$�=E`�_�O'��dt��+��(�4��;Vif��i�<Xk�7Ri�+�8��\�o����#�k^c�ٚ��̫�n����Ď�Kk�f�����Ԟ/���,��UN��ݻy��Ǹ��g�Er ����u�ڿ�}t����w^p��Q���-��;�9��J�Q�V��z�F��_
���|'4W�b�o^� {���ٚ#������ �?S�-�qp�R���\,�'�މ��L��As�s��YO��U�wܗ�Fa|H�=�`>l�5O��ҳ2�=�R��VI�/Ua��~���vx}|/�W(�dY{ ����{>
��b����*��y7�b�H�G_���a��J,�s7�:��O8\����� ������/Z���`�|��������4R,n������񕘄��`fU�Yk�	,й����h��:lm,p*�<�Hp�#��J�`�X ��]z^ ��JG5D������GMm��hn"1kcB���N1��ޟ��� �e]8��C�)@	����В���/
 X"���
z����tMZ㥫,�sMh��,T�[�*�G���Q!�`�T�
>�^

]Jf�쁜����/�c3W�k�M{�ZMSC~AQ������U�v�NԻ�V����̪���`n�Bֽ
q9�ueY�\��!KH,�<w��#�_����E���ɩ���j�'�l���֖���ރ�*�Y���¿l$���:ӊ��n��J��T� W�km���ç��W;�Ѱ��kHq�V�3}V_Nu�WF�5a_w&�M������T��Q��\�_p�s�����AX�u+xb4�H�aY<�h^-9�SS44�;=��l��(��HI<	�/v�Ps�\�����.#w��"r�L��~�U�k�L���	��;�6横"���t�����������������K�.�,1�2�������t���r�RP���D|��4��P#��7i[�+cb�V��?Ɉ=�>�,�%X�{�����>�/2�ma���o�c���(	��/��C%N;�#}�ߊ!�fl�Nށ3��I~|UT8�!��+�T����L�41������T����Η��#*X�7�*WEv�����U焻��q��4�m0���f�'��O�\�A��r�5&�D8}�L� }��
�RO~n@~W�W��O��R4����J���B��
����}�P�JIE�r٤]m��m�h.��H,��즥�z���;�6����]6�ѳ;WO��+#	6U�E��'4K��ϊ4���s唷��']�N�k7)^;	yk�=�R\�Lb}>ck.���y�l9��>� �o�/�1�Pa��nI\��i���� {�m\R�j����K�6c�7��r��O�g�V928�|�=8QԩK�c�׫��a�ғ;�6�B��ԪؔOl���gvmH���PO.��"R&��:P�
�k�	(~+�������}*�:��3Y�E��T�<�Zr#-dT�4?��(���֏���չܺB�+�1�n3��ط#/L����!��������`��88���[�5s�	%�|���HWm�Au-&{�ޑܶ����ػ�%U�o�;�$JEK=NHb7<��}�Y)��%o4uQR�̧u�(��<�J����Z�w%:=Y�
�Jq�1ө�}� �r�Ժ�&d�z�S<�� Jg`0���vXP�qٮ<�y$?F��#�fr<4TL���]�r�z%҆�ϩ�$Y�l<J��|�N��S+;-��'�o�z�)�t4>�D��p(�x��G���p4�\{V��"�����;4�2 �皩,����e
ѩ�8H��3��}�I�oZ�������1�;hOt�������E ����PO$[�i�J����xN��4!��V�ص���h��۸L�z/�N��]1��R�:�V}S3g3�x�y���헆�D��|���G>���b��*p��7S�g��p48Oj"��w�C��M(���hoab�h|]�ߏ^�� և��2IR�tS#���f����Ư2�D��g<���P�j*��2�����EJO|k���C���Aiɴ������ ��$�w��p��0��JetG���k$�H��Wwr�͑j�Y���	5f�+�pI%��_	�ZS��� ��Wr�p��[1r���mm6�r��'C���m�:�p������J�B�F��
h9= ȐDW���Z����N�Pd�py<)�W/���s�[d0[� �f^4 J�w��ye��w�Z�����D�1��0�8e2�ε撰��21���{��׶�P"���OAj�Vѵ��r�'���&?]����r���+T@�>��䙧�[x!��.���ފ��P؎�=k�H2<��'��"K�.���s�^����ƚ���?��k�G���1�L��X��>,J��N����ջz�;�gx)�ڳ�1݆K�s2^�|Կ&�64�����U?�9S�Ǩ�-{C�9 O��jd��>�m��2�p~z^����T���>�A|Q0�.��W�l��������7/�^a�6䳂D?~ImY��_�K�ɪ��o�cz�Ą���J����B`�Y��\g�Z��;?|Bq�: �����{r-o8�6/#���Z�K���G~y�����X���>�
Q�������w���K�"Lp����N'N^�5}o���:+4,�w����$%�^bڑO������-aUD!��\�u}����+f.�N2���.�-!�����A\�-�En[)^w���N��f��I�ì/j�yW/z6g�xU[P�b)�Nݷ1re�6v�1��S�2��dq
��L��D��	T�/*`�4L�gXNEt��?7K�1���8@0�Pe �x���D�['���4�*-9OF���WR�N�fIGI����h��2EX���H�j6=m�DB�zu��5HE"R�I>V�"�,�O���4��x�@̱w�ղʺ ���M�
���Vq=��D)*�ܬ���+G��L��X����3�;�_,��nF�(Uvp*[�%��|! $gP�`{�̈́�8��Iu�N�,5���?��n���T=[\[)%*� �ۧ.������ݾH �L�Mg��-�j�G��Y0Ů��w�!J �ح��|jC�zb�D���.�{x����6��s����܁<�l������������)љ�o���1O�����zB�%`��L'7P�,���d�8y=Bj��x4N�6�X?�iߧ�H3s:���"ȅ�T���D�����VO-]6����O1�Ɓ3��_j��
m�'���˓�7s��K��`O߱�K�l��է:ö)�~�L��_��&�@�@�he�%�s`B�����Nql�\���Q������dq>��Űm�Ci!�͉��eZ@�3�y_�Oį�~;r��5��wZ�z��� ����6P ����ͻ�_{�9=\$���gcb`0ʴQ�Yg<�/���N��Y"߭#p�R�,-�����,�����+����0��Bz��ɋ�������4N*���U�-�j���{:���C��nb���mpF'�~x�Y�8VŶ�=&�:]�����]o�fHp���u�#҉��\�R�?�ꦖlQ�wM���z�Q��t;���W,[���Nb�5�ҏ�Z��Q���gW�A�%�	17�&Q3_d��M������̏�������ܣ)�?�-�EXv��<���Ƌ�	H�M:VR�)^-\��	���r37.��B����-~Z��EG��ޝ�/s��_�^�?�ٮbgmD28Vz��E'g���E{E����bE��:[��Wd�G�Rbd(��+�T:^/[+�!P0�2rj	��`�7L˳�A�Rpq����=�Tc�P�(�ֆ�t����WA�~�eg+U��E!�$��}�nE��<�l��>x`^��C�F{��*��?������XLt���k�?�a��_�qґ��M�
�����N�o���c�;���2<J�8�L�'�Q#����0J���Mh�%���7�9�oM�*�xH'�s������S����.O���ۡgdjF�_ظ���G9��t"0�	�4��IR&�'c��x��N2��Ń�8�ML 	���B\i�u�b�U=K��ue�n�*5�	��5��a[<y��S�nL�K@�Nk��f��&�|`����g+r7�15O�f���j N��^I�)	1��E��R+1���n��w�%�?`I�'H�unQ�ƥ�B^$aY'�Q�nAW��C�O�d��oP��,+؅�P�E�n�U�pT�6�Xz�덧�p�� 5�/65�t\��Ƽ�09�u��)��=�dp�*LՆ�Z� �^}<B;�Ҋ<F���4��Fs6[߾Е��f�����?�M1"�ic]��z��)��X�����[Z4��[Λm����cwzE��e�@�A�кh3��$���|=������b���g�)_����3zzIn������W�t�q?ؤqY'�X��8G�o��=�����Ag4#nW���M�ͧ�ҍ��������}GW�i���B�����+"�����*��+�ĸ�*1�U�}�
�5�?����)�v�,��Q�!�o����t�Jۏ��K/Q~���e�E~ح�1����Ȏ�	�H�Z���L(��y�������ԇ��[R��2��������LUZ`5�0���Ҋ����B����L��ӑH�n�x������k]݆�zQ��S\H^#A��wS�) ��y;&�.����n�$S�|�4q�q�k�':6��H��`��N��"���Q#���bZe߳�t8��=�KeU?��τ�}�����mߛ���9�������KW�
q!L�K�F�?A�O`�0m=-�0�Ĩ@�#;�ΧF=n.~�=�
�!���gp�6�T�=p�R�����]����b��]� 9��x.�¼��*	�'�!����w�ks�Ӕ!��yCvY!Q@"䳰�[�+W�ss5a��HE�cC�5B��>��c�OP����w�,����R;\�<���ن��<% e!�b�,l1x� �Ҁ+�ly9����F(��"T�|"D�q��s���:-�F�;Z|�+��;��Х��Q�����x2j�d�=�LBB�.l��ҳ�B�x#��i���	���i����z#��'h��@�|Ě�|�
����;�|գ�}h�Z��q�a�n>�!~h�s])����ģ��ꖦ�"#���C�l ��?�j[?>�B�0�r i�=��ҭ�s�˃##>�rPT��8RF .Dnͣ�<"�^�Զ9�0�&#ez�N�[�eϋ����)���O���ב����?F�LO�����)s��ĵ���UL;\�����	,�Ҵ��o�嬫���Føq逋����b�HbIS5�R�6O�6"FOAΒ�T�^�>�����ŭ��D����{g�@�!B>��Y�\�ߠn�~Hjs�m��L���ڂ��+"�1y�t��"�r䕪5,���7�l�O��t��%bs~^��w0��'��]�4	�����T�$��&����L&K�d�2Gw�@[l2��7������"��E��(m�?�� �]�U7q�m��b����a��4�XT�r��R<%;�v�d5�;�!��� �,��{�	�9�bO�c�P�[����^2�p#���GߵC�J���x8���{4<?��i!Q]9��f��&�x���7���|�G� !�y>����oh�7	J�X�������kzǍ�3��~+��� l�!G���#��=c�p7u
�����d�:�;�bz3����e���<�B@�� E��;�l���뵞|C��%/E&b�	�:u��779{�_�Z��n}�l69��N���3>ܕ,vW�_1D�e-����TGNM����(�[��q埖�9MfL|�g�ϳ��[�"k�}[�?�kqfo�>�Ca���:X�������}ex��.��}2Edy�\����J��Ϳ��&��8��6S�N��kD�#>PMz��$� Gm�o(��phI-|����^ַ���D�wd���i\u��@�+��G���<nJ�ƚ2��3��BCj� *nc���&���6�F6���n���߁n���tnQ�IM��$=oT}����JxO�Ka�5�p�+��X;DˮW���T�P>�-���΍�rlb+�i��av��'���Pݔ=ФK�I+�N�a"� xe=�ћu���ڡ��;;1����~�,���W�Q}�٧1WMn�ǲ��t
�u���ȋX�E�^��-	 1Rc{����)@<��b�~GRŚ|�c]��IHɈ:Ȝ�h�E�Rt�G>ԓm��cp�:�h��<@R^���t�.pǕ�Zlu�D��v*:h2�F�n	Xj�N�TQ�b�����ܜ0�D��G��D��P�f0�q�V;�$K�%��u�@���O���e\�Ψ�5�%�Z�gC���
i�T��$����{�&��Q�ӎۖ]�[U��1�3<�nT�^&��ft�_8c����H�n�-;��	3P�e�*lV��n�t#�*�μ��F��Bp?(kw
.}dd�Ԡ��e���6���'���s���$��*���U��[X=yr��,/]���ZU��π� �@?��@�V����l��1��}pS�u��/(X�*�wAӿ�^{��i�:K� �� ��C�q�*�CM�q�����#��WdZI�ig�UEֈ} }8i~7e*��jr<����+�Ʀ�H�$_���^�X���%�i}ePmz8�v|ZHCˉ}�!_m�S���/�Or��^��7� �9�T�����o��t?t>��t��S��bn�mQ)�� �������M��m��8zY�wg�����{���4��D�~�gĎ�����(��п��N�_�l<�;F���/��Rꀆ��S��bp��{՟�"�"�V��a���݁�<_��EQ�u��Q�i�b՟:ڿ�BҪ3�6�A��D�T?���	���]�Y��:�j��%�"�C�u%�_�6�䟜K�ӆ���2)�����@t�z�)��l<;K�Z͘ox�+�eKCm�@�]�=\��������<��P��}c_ȟ�J�@�/H��ө���מƃΟ��� �H�S �@�H%e�Q�n%p(g��0	̟���>�ҁ	q�%��\����d�u��t\Ghs�a�~OV�L�%��g��~Z�Z�+�9e�3~�7 Z�o;����Pj�/"��&��s�%`� �Iz��W/<�n]�"��N+�7����E����,�oCJ`Q��F���I�Kxs�b��3K����fs�Z��:�;4B�k��7i�GdK��m�4݉���9&@�ɞ l؅26�5R���q�ch��l���_�*b$ݗ��u��b���|y�v�a����h�v�%mK��M�6:_>3F}`�to�!�l𨍼�"�wwF��V��f'8�yU�Ό��fB�iؖ�p(����v��+�H&;����Y��do(���i;3%���×8,����bLk���S4T�'�C�#!��hXx����J�E
�k���=�٤_�g�\���6wK%�w���r{�eRh�-��N<�Q�A��p��a�a0[��[Շ��0��Wn���b'	W���ZzZ��$u#�[��,�j��B�`�(.�nxX_y�o]3:���ާ3��,��%��~�&��L�~��^�����)�`hu(��JA�ɘb-k��Ȃ.]�4ص�#���{��W�t�0��32f�s��g��+�'dNM����V����e\�"�w���d����Vx/$�)��|�X�����х(�+jE+�@z�{"C��(&P�U�Ҥ{������ L\���C���FzK�`�(��X�p� ,ÎLg\3ǲ����V��Z��u�j��'fk�r���i�c0@\s)��ox�r�=��UX�5�=�JslN�c����#�)A���T�4J����D�rhN�$Iw[�I�,�*H�d�]d�0δ�>g��n�7g����0QO���Ձ����uy�9��:�+ ��2�m��bw�e���A��!��ƣ;7�*dQW�J w�݃��7xr��ۏ�	J���g�}o�x�p�z:o��,����{<����d\�����C���v�4���a��§�)�I�� ��4��e)�u{�q�o�dPˤ�bZn~���c�#ϰ���7�R�^�j��٩����g�U����o��6;�<�U�F<(�Z/!ɕ��Ū���TG����(�)d�P_�=�k,�|�N����%A|��)+�g-uFt�Ͱ�L��2��"�\�ǈ<�,��{��{�_嫐��c�3�@*�:c|A�)�(���������%7���3Cÿ��U������5O-Y�(_�`�
 t*#�4�O��(���u���A!�Z��l�Eೌ�S$Y򒥂%���ӏ�SR�֒��d����	��8G���ū���f��cSn��,���u"�x�&��w�g�ͮ Wǲ�m�St
�P��J��h���|tB;ˤ�8�;�����B�dz�xZ,U�p4���>w?bߢp�l ڌ�
[���Vx{Њ\W4�_���Kc�k�"��#�� ��6[���/�c�`�qᏫ���J�gf귇�o*Q=�g���s��Q+9Y�٬��0��X�)��>[I|���&D����`̾���[~�ݞ���#FC3�(�%�y�{׵�5gMBm!f�d���'L�e뷜b�SD��>��ff6�~�4Y�������Εpܔ��v֦�ڟ�ĺ�~|��l��c�g+b�k��[�Kl�XՖTea�����C ����w|T;����a1�wW;�:_C*�@#��0��ޮ�fצ��WܚcM���,�5'V�z�/si�K��Ԭ�K�W�r�1c�-��&�"c��[�-T{��ń�IEk7��0V�Y���2�Ct��j�.�!�X�l	w@��ه
�	�]�紶h=���u�5���R������C��,��MY�F0_��:2���Iؗ�r*��|X)0}�"g����Y ��%Ì�V�����RJ��0����O}�eb�C5M���M8�B�p�ķ�.ka�L�<9��$��c.@�Sr�4�,�B�}�,�N�Vߔ7�{"�2T�ke�6@�O����TY��J��E� ⫬J^�D2-�{��;�qa��o(�����h�㹨m��2�{^��c�e�����xz�!Xpj��K�*�u��(�tS�ނB�uY�J��D�Z:�ӿW�mý��[�&vI������\�Ry�U�(��Ge�������;|����9�����֩��v�G?Z�
�}r���:j�3K)����6Ĉ���k��Y�@I"]�g�t��H8���E���F���8O�+p�Č��g�K�DبȢ��*�*x��/	r����,�u���Y����Y=$� >K�1\V>���o���w����h:m����%Hii"��%��Ȩ��+��I��X�~Th�Ez��B��r.����,c"�s���©t�i1�Hȕ�$v�|�lNӛA�ӓ�A>�Σ��Ț�M�^��k�����'W�ե���K������wԜ�W�v�eo�Bf7z��cJ�R�������܅KȳЌ�Bۅ�fe�}+,�����֍�q=�;%�>���#kK�P�C;P��/kP�X	%G��
%�B7@�鸷��͍��+܂�q�y�]�;M�5���s����M��Ώ��P�c�'�Wje:��$g�H]t��uR��o����2RȤ;E����Z�l���g٬��U����O���;��k��MV8�K �Q� �1�lm�'�?5��=�h�e_���o�W��L�����*e`D����)�a{@��D`�M${`Bم���D���գ�G �),����w���X��m;Qr�FM���V&f�6�C�:b�k�����^	-R�V�þ(��J|{+s6����l�fʡ�W�3J�%��/��P���.ԑ;�7�Eː�5y��E�rM���g��V�Ug*�+9���ޏ����X��v�B�g+I�}K2^��Fa�J�c�.L���Q�F�"D���Ѣ8�g�3��/��i�@�y?p��HWI<N�y�;���U̦7W�+�"��P��}��Na䳡!V��t��>#�&�9��,��aj�O±���?c2u_6fQ���/#�L�5����(D7��Ep����� u�l�]Ys���(e�H�������X�H�0hu�H�߽�ʴjk56�����,G�J�/��󯰢��c��̬��*fJ���vU�Qi{x^�+�D}�=p�]-�9�dw�z��xa2n�%�p�'��U�u��Vm�8�&���pDa�Ix�5���?p��I#��N����p�hM!���l�R�q���y�)=Id<��j&�+��7���	h�Mt�L�͝8,�B�%�(mo��p*�ʙQ�eł��=ISfP����C�0�5�����w��_�{�R(�K�;�+*H/�Qq�����I�S�E��N��T&Et� i��b{#'�����N�mA��v�N'�k
�=�������0,\�� ��ƪ��LV���L���2�N&1��l��I����M���n @�`�Xﳫ�ϻ���Qj�����jH��z�`�n7������������=���l��:��}��*���=�i��,�v�Ŭ�8<��J��H�`���� ��v�?���;��t�RB<����/(	C����Ӹ"��rl��$�b زoS P�p�(ą���q�򮽩(����=���>Mp!��X��*�[i����qP� HVd����>*r�lf#�?/����f���}����=.Lܶ�A!T��o�(�����N��(�x���\a(~1ъ(�a�����2�n-ܓ෵�S���Q�������t�zķ��6�m�6B��0׮��
/=�*!:�0~8d2K����#��#E߾\\�<W���b�o.^��Y��3�?����p�	�K��6j��}�n#V��(���8�~��/�ݛ[AW/����j���u~�z��?��ّ��x������Ȧro�$��Wx�G �z1=\u��V&o|z�<�ˈwט���O�~{��PB�����bz#�k)S����o]F��{a$c)P "�`��Ph%1�TJ_Op��G$b�#�ۅhQjL��톗ev����v�,(��օ����a}mp�;P[���H�z>�����G��������=54���F�BD-(������DE�TG�<Ih"�ѣo����C_�ev#�˩&H��*c~ɞx �����]㱮�f7u���]5���u�w�ϗ�C�+�c���:�h\Y��T�=U��y\C�#�Q1����	�L�o��V��Q����?��'|D��Ê��o2�!��_��'�0��O{�$�Y��*�r!��1j��+�c&m�ö_�{�y����݄5�����;C�?�	�/�����n=���#ihTEOJh�fv����m�ɞ��_�р���潗a�u���=�ip��ްS|��v�8
�f֐O�f5�b�.��ow�^xMS�� .��Kff����2Fؑ�j���]�p-f����B<��}I�*K��?v�CY�3�H9�^7V�b�`U����~ />i�����W�z�3F@�,�8ɣm���Q��;�r��k�'���-Ih#ø�o��ƙ�+�'"��wU�_n�gb�ꪎ���� Hp���u��tuӹkץ�b9�:`��"��qm�V����©	�w��D���o�?
rsn�!m�b5�-���1v��f��yM �<�������x�ށ][~�l���-�n>��U��_��#����J&%!1�YFj��}�y �Fd��!ߺ,��O��8�����d�=%4o*7Y�S��߄��oB�D-�J�Ψ����w��DҒV� 6�����}����.��rPI���MNvԫ�C��/���Z[�:f2\Z�wP�^E�T���}C;C\���Y��I#���E6\$����x������-髥�i.��)���л���-	�]cF�&﷬4�rݖT�Yy[i���bgFy������2�hߊ�K�
k�� ��b���� �E.�#���O�a�;Ю$���J��3b���w+g68�)���Z��}�uYW�fGQ�� m-0����b�x⻱d��{�;cʹ��e�н���8���Sji�.��t�/|���khGO��R��]�^_z��0�~��2��\t�\�ǳ���ݔ�e��mJ�Bi��=7����r5628eG�n�̔�S�l� J�W�z	M_�^�8ǀ����۟��ՠ�|N\��� �#mJ��N u+^����Ϋn*��$�X��،��?Vx���vMo��)����_���,�0��L����~�JPEب)���!�(�=�X��˶Y��7<�#V����s����<�`[;Wu�P����Hn���g�aq�C����yd���z:��-� ��6�����r,��@�s�P�j">���֜[Y�����ڷ�T�����jꅉ��4u]ǽ� d/śY0�{�������+�5Nq�w{��2{����"}t�q꿕	Px�?��U-�Z4��w��`���m�HLr
� c��(���l� �Wy���@��p��Ȁ�IMcr�#�{,�e2�R��=�k���ڵ�_W8W�ی�v��Dm\8*]�;L7YЦ�%n�d��RC *�@D��j(ץ�_��xf8ݸ�"y+4�9���p��/$��h����;��'���*n��,�v��#��=�� ;9�B��S���3�M���D���^��j	j;�t�Fo ��o��M��sb�7R�Ira�D;��h=�O[�Z���'� ���@)��:y/��{����
[ɲ�s�.��)Â�f)ӽ����m��Rqc���c8��`�>��i������*�b��d�{�qCG�F2)=�u's�$���#��4�1������Ո�9񇌁fl�oti:���K7Ab��G� ����Ǟ����4�h�|����	���=�������B�G�6��)�Hv{���/�DC<����U��T�J�<�}�ww��d��ד���]y����RY��4[�u<0uM����pu�D��Fp�W�vY/�����������*ǵ�5|d���L�������A�?��9�3�!��J���t�����oz_}�u��zI�i�0j��t�G�tH�����MdK?��c�Ӣ��w(`�7���|�4Cu��&�C/%b/4dI���JxB%�Cl
����u-Do4�e�������`^,K!hGF��eӧ�/��@
��*U�R���z���6@y�`u�^���޷ �Mƃð�*�da@D�v1"\�t<��"+*�C�%������r�0���Ɂ�)a��>DZ�o�S)����8��r��v��`.2,.*3�i�M�1�Ř�T[g�V����������;��M�V��	�� K7��jc��äaF�)V�5ͺ�$lsq�C���`w���o<")my��5E�#�&�_��w�����;�_�%l���q�g5%�1�D��\�[-�Lv&���'e�?倻���c�+<��+�NO��ZR.m��酯ڲ�����ݎϼ����`O5��Q*���;`V�L�ϑ��ƿ`e�����JK�IK�cj�. w.\�����@J(L��4�"%� /zV5 ]�5!1(ސ�=�R����QYHDV1]\�^M��}�!��q�	m�{D���_��8�q﹑���X��?P#Z3���s�n�-(i2��1�͏��@��c�Lxl�I3���&��w��	6{֔�w�e��J���1'���S��4�_�Q���͞��EL�p�0yg�Y;-f������!~Ob6R~7 �?֏�����1u���D�NI��8����E��.9�	jfշUmc۬�C�Pv�(�L0�DPð���v9BT)�`v�Ց��nv�'�7�I|��w��{��2���XZx�O� �ր��1��d����v�|o�.���4���34�7枼��˨/b6��"�5Y67��W�.Ed��zq.JE?p-�Z_3��+��z�@BU�r��~��bo����V.~�OI�<v^�,�
(��Aa���晡���;H� C��y\.𶹡��t�"_���^Gv~81s=���
��� ]�T�|n���L�)D�ۋ�-3i����,��}>��h���gwo�%�����'��R�]A='MQ�Ū\ꘊ��|i�Ft�&B��q������T�Z1mZ�QP�O:hHhS���d�p�c��#�#�$K~�> !��Yc�џ�[����c]#��'���J���W>�P���6)��O���犏M�M�G���3<�;?%�/�P,Ya�>3��:�G���O�ZŦ��_C�e�I��蟾�X�|�5<�̳���3'��UZ�Wdv�l�ڻL*y��>���JB�4 ������;4˿���!e�h=����<����`0�C�����YZd�?U���ר�����l	�O\ժ���JU�5T�)��^W�ʇڍ�փ���ip&"HT�؏��Q#�K�[�u��6~�1�'�{�$F0����bo(�Oe�1�f�I����Os,Bo��B����2���y!/ϵ��j{�j/"��
x.w0u���_}ղ�p��K*�ة�q)��+���j�mn�/�M����dW�ՠ8��A���s���~�@�Dwe��"TMo+�
������g,�x�L�`н�7^��,`�YZ���Z;���������6sNdƒUҴ���i	MF��\�����C��	M�R��{��mBj*���f���eo�5���
U��rM��$����O�]RgM
x��%h�Y��O�����H�0z_;I�+��å���
�^����4*����t��Z�����?�����/bu��$�cS=x��Q��;a�v�0eV}���Yx{	\[`���ԗ'x��7�+ecS(O��A�_sW��&q6⨻ѽ��b����8�	��+�-��lIk��YNU\�a|��v���U^��q	I���9�)���"��G��$�&|n���9���z��F	Ґ��,�R�'eg� �z$��6^{q��Ͳƒ�����T��>�H�w�|�r,p[��-3��S�2}V������6q��9�6s����B;�%w��E�y����p��"��ƻ�I̕=�(U��`%l�W�kЄ*�8׹{�T[Fy�k���O#c@�3	��������]E_i(�U\O�W+�^ �0n/1���/l��_���m������4�yǍI�ԀI<����&��_� �3�"&�~�h��	/~Xݺ��s��jɼv5ʓ�E
>�@w�#���˃7�6ǁkp�}�';d��ï��x�����к��](�7���G�;c�$���D)Z'cn�w�����_���OP��Q8����6m��P�O�!%�#�3iag%���(��!ߟ���8���Brh���x�r�
)���8#��[�;#@�*��'���6E�N�i�n�i7�"+c�Rwȭ�-"h�B�J_M�37��gͺ�� ��J.����c���@�{�P�R�QϏ�۫8:��wc����;�-�擳K!�Ҿᔘ������`x�i35^�M]ڼ��j+�
7r�g|&��w<o؄	7j� �ܙt�E�o@o���{�
��p�w�F�?z�]�Z�Aш��:{�F�y�]|�]#��OК޲�e��9H��Gs|*�� ����uo�ڟJ<�y�}�,1gwf
 ��g^��ҡ��`�}9���(���P��	�]s��_6D������t��r/�N�/�����j\ΉrE��c�
��&1X���:=�N���,3<��)��Fɯ�z�x��ef��nO�7wn��,�WC���4�u5��Bn��(<���� ��_n+���a�ު�1\樤��U�=Bǥ���.0�c�܄�4	�<wTb������cg�!���荃	D��}�˨5�����q~n؞�� ����ϟ��Y Z���%_�ys@�J�\t�����L���C{�$|3IO�Vd�K#c�����j1ڰ�'w1c���p3��`��tsQ=]�`)�4�oY�yP���G3C�1��̤���x{�)G��`iM,�Aw�?�� ��^���;���>�H(�E��^F�L�B���B�i���1u�8��0z[]�A2zZ�O���	��ܐ=�%��$Ǟ�� ���b����
ߡU�3�ۮ�mb�6�O���ʩ�5�64[یҒd�E�]͢��8PU�<�Z�v���k!�b@��,