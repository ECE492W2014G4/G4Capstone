��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P��v�"<ߞ��&'��k%P碶�R�ӣ�sĞ������FY& �c�]�f�L$zqi�زwk<OKc8VZ�6�Xș�;RQywSW���n��>c��\Z�~1��̀���E���`�"{�2�/���3�\��J��p��b��[�*��.@g[^�ߡ��v(]Q�����P֮�cq�
�㴋6�sR\,��@0=�l1wāA)�:L���~���c��/y�jmS`�8K'���䄽�K���z���9���X`+8hܿ���(��Z�ū6	�!g�\.Uÿ1Ԣ I>�u^�8=�u�ra����'q&7��t�|T�j�A�
�(�@���k$�;�*�\�7���k�c��i3'��Ōx�;�$���_��u6A���,��;x���h&-2 �`X�N`7~�A�9胩x'���>���"v��D*HD6Ib�����~c���)q�dn3�	�s�:�I�u
��;�k<���G��%����QE�7��ŀ`�եS���������]�ZGg:3��@�BJ��+�V��C���B�M�]���Ԁr�ب���bQ{⧇"}V�!��C�������g�oM&J���	_�am�wX�I/��j?�􌯮�id�="�-E�Ψ�����$Z�N���ny��� C��W�ζܡ��c[��U�����a��d�l�m�㘺���~���{�Sfl�{#v�oN2Pm,�4���E>�qe6�<{��b��G�Ż�P�S/�Pi��y�"yw�u����{\����y����M�#?���5QVi$r�r!EM���IW�,�.��!oDZ�J+��Mi�ƷJƯ��_j��D��qx@�dR�Y��G�2r�")����P
���Rw��P}��M�|���o�N����F)6��l�[���9:Z�G2��5��T�:$�0�//��܀}pU�ex�k�!��x������.��3P2�,�*�Pf�ӊ��iEü�7�(Woe���R�gT����6I�̋����ןv�&~��������3�/X��aj��o���rF�G�Q�6����D�њ-rQW�y��m̎T�2��{(Y1'��Fo�վ�㔘W!�(��hP�7(9����G�O�����Ƶ��E��ii֧�pi�/bf����JЀ����Xg�|��S_�����K��~^Fŉ�4����qeA1V�[?z�э��q��V�L[#|'_�hq��p��D���uˉ8p�󟥏o���5Tmg��*ڜW+�;�}�C5����6d��E��G��Y��kY%b��(5�
�:�u�D`pԩ�j�xƯdY�N�Ӭ#����8lѹ,s���d��`���.�|i8_eg�-0W$�\�i��?#[��!"JAY�R��o6��t&_����uE䉐_�n>�梐ڛ�P�H0�{�X���T��[�l�7q�H�0�H��t0��M�-�+��,q�8\X��<�V^$*>ڗ7�4dd�E,�r�����~c�(FI6�{}Ws�L�Cv��zH#�|[���F�f;��Ҕ	���F`Ð/��*K�q�7���(�p2e���}-�/�* ee"�X�vf����~�H�?g��ׂA!~V�����4�gE+rdDey�K�JA�R����o��	�GO��lP�7,�/N ��}���F��I�%�ͺ�����K/G5C�jF3���E�߱w�JF�!8�����\:��.��{r��0:j�qsv^��`�м�r�x��]����z�!�:�O�\q�Op9��r_@�G�#~��,Q�G�B�V���h:^���\|!�6/ү|�Ư��ؕ"�]�s�(k�>ڋc%�A�&#���}�| -%��_3���a�+�|�z\�Ų=[�)�\�l�{}x;	���?*4�7�����q�㖙
��d0a٤ت����ݣNB��rƹ�����w��X����O=����xY���D����1Y ���1{j�7��$���2ǭ���p����&�x��r??X�����
?�T�aߒ���J" O���pG$E��T�>�`-�t�ˉ����Е$���#n�'��l���"��K��؎�^M�n�Gе�k���lu�iu�w��2Z�w�r�Rz�c��?��E���Wܲ:���,�KB�;�߭�=}�9�3VTɤ�S�ȠY�B����i��&��*VUr/���!�ۂ�� �H��.Ia��
^&9�p`���*�I]\*r}��ԧi�eh�.#Ƌ��R~�/钯�­�ZRFMp�L�<ɿV�L�����>��d��KŪ�C�AU�QIfL��0�9ķK>�x� h���}�o����Q��΂�:Z���e]��Vh�/���U�����ݥ1�#g�`v�X��f0��r[��=���(v.4`�v����Yą,����h����7�-|26/L(OuRlCl����?��N`Ӷ�0	��;E�������1
��kdå���߻$d2��$$��kY J��\4��ݧ�?\�D"�GYs^��%/8׎aA�x@c�	�1�t����ڎ4�Gs���"��Sφ��}�$�
s�<����si�i�2rJ��3g��Q�IB ��"cL`v�OŰ������xz��� 6܈��E2�����;񝈀,Vz����²�^�4!f��>@���M������������Į�+�<���0��h �(�a��pU����?(s�q��D�'0�	�6�W��7a}�A����]��g�Y��黆n�*���;�{=����V��(�=N��R�]��КC$���_�N��A�P�_��J$�U��7a��3�A}�o�
�p��	�
�x��1ڕ�'�;6��䵆c�&ȅÜ׹�xƓz�"�qx��u��9��|��&����B���>�<�(�S8�<Ť����e��?�47�g2{%ܘ��l�V뜧�fÏ��3o�s�����O�� ��-�u��Ɵ�!�`�ĄK<�
ܵsΙ���; � +�~��z;�U�R�Ę�8v�.�a�O~QuE��h�b>x	���Րd�<_E�����<�X�b9�CX���L/���Ed%��27�L�jN?��>8Ɵ��q�vy띔��':`
i$�8'Gut������"ÝziePZ[��q�0���`I��=��զR`�QƔE���{@�>�Ҷ���;h�� �r�_Y�us�U�iߡz���7�:�4_N[��qJD���~�xHO�_o>��Q\?����/�3�G�"J�i6����+7�����h��+��ʛt��KΫj�gѫ���"�bY�)<�`TA���AI[.�ׂ(1��f:�J���gO3	�LQ�W��Grae��K�sx�SD��
#m�β�X�"<��\��v��&�23ic���	~�F|׋�3^�����򄱖�m��t��QFrU�&�`����_x�V�'���[p�hR��N��7B��7��.��;SNYlf����=�Ϗ�g��nx�&/��p�W~�ҞfN�X�zw,�BN�=�%�l3����/]����Ҙ+f�t�u�OJ(��?/�<HZ�����<L�j��2A@��ƅQWy�KA�keK���H��B$��ی:,m���/�-����oKz�8y}��2�Du�ˎ�����|a#���kX���^8���)��}T�c�����D�����!�b�KOO�Bh\����/ȏ9�q�g�a�4�-V��O)�7���gaa7%:
�����-���`��H�����0a ���+��7ee �aBoj��C[�'�$�� �Յ�|�t�S��1/�fo�,$�8]+	��wPuc����T�:\��.k�5��{�YE{L<���Q�rd�!�-��r���2(�.����~�|��}�5�~�tK�P� v5B�Bʎhg|�=i��m��;���I9ލZ�ǜ\<�R�m/��g�B��p?QqtM e��M���+Al�A��F2L���HM�����_���"n��>��y
1�����"�Iv�E�g� �W�Fl��z�Q8�`��g(����5�ɱ���Z;��d�b�2��|À���om�Ga|�ݾ�+���������cnx~K���:��w��	�x|�K��J�f���	��uJC�
ՈA��:v�m�9���-{z���#'}"���<R��h�4����"0/���,J/����*;ȧ������Nnq�Ht�t9�}��@eT�ZƘ71�:F8���U�;U�d��Bb�J���@7ǝ�����ZS����A�0O]I�� Yg�S,l��Z��]�X�=V�A��Y��b�F�Ӄ����5�G�zd!��y���,�m��[�V�F�Ye�'K�hڶ�J8�_��Nc=�/ϋ@\�]�
�-�������}�UP%�g����jo���(0Rw��0��ϰ��畤�L}������3p����v�
�F�yA�~'9��� ^�����a��wpO���Ͽ�:���BH���>Kf�l-��X���77/��d|_�����hz�ަBS���И�ť��ѫv�vH��:ؑ@�K�5��mQDj:�VJ��	�8$�$�vl2(���d��%�D � ��rV��Kw���a���a.\�w�^�A�;ůJ��۝���F�h�C0��v:	v���D�g���ĩ�)��N��Z��8@��F&�ф0PPY4xЯ�ߢ������/� x��u��]����"�y6��mU-�	����/[�o`�Ɣ�/�^�q��X2 �R��;��� �؉css��0�X麂D�ci��˼yI�]ߜ�!%���=\�<�� ��7����Pnz���2'��e����yWnI`��ͦ+Z2"�������� 3�N� c�8��o<\��6���8|�0���!/��5U�·���&��92ڮ#�s��D/uIlo��e�z���������l������.�9�Q�j�8Ve_��:�Nq��ﳁ�h��o�����l��cՏ�1��[�՝p�w��q��/Y7ĸ��P��np<k���YؘIw��5�$u����Б��x���(U������/tV`V��`d:�v��Wxq�T�����ƻ�)i7&�AM�S.�Ɩ��>���8ڒ��n����a���b��e�q
/I�vw���KR�@�\��V@�]�w��Л���%��}�@d�D(��q���<d�J?�b`����E��/��ݰ	$Q����\A�~�;͊(m��qE2y�3~>���N�`CЄb7$Y��Ը��f��Hs��KP���)�FAD��H��48c�S8��B����?�d� �b����OP@�l�b�:�X�CZ9h�2��� %A���H�%��9�ێ���LYi�6�V�Ƨ{��Z�D?q�>��~u��E��O�uK#\�Z��|]I���;0��վ��	�ϖ��8L��b�봅�5�-���Q����`^o9:ze��������"|q��+7��2�M5`~j-�X��R �����<�T���;���q��8L9�0R<ӰsP�S�+��yʃH�|U����^u�J�Ɂ�����Ga����<�;�h��.|-)�U H�K[T$�7����K��&��-�^�
]x��N�D��{���ď�劳{q%c��(�f��m^7S���<� 
2�Na52�%+?��րs`�O�
��UAȜ���|); �5��q����:��,曹q�)��|�J��1�S�����/�KQ-A౼pl�-�XO��D���=�\��B����r�Ģ�DrJ}v(G�%��-|v�ne���i��������f���͑R$��N$�t�\&��7{׍�10�j2��H���WT|����Ac_���\F�ى2s�g;��	(���R��0�R���LE���o�~�8C`F���8�t��GD.Ķ�M�ͽ��p�3O~,�p�$AC�M�Cy����
��s/���o�+��uJ���;J�����|�}��ą;k}g�4��X#	(� f,_N��D�S-�/s�N��T����l"g/`���ur��JQ7v�4n�v�'��.��n*�| �b��P�?k�rD�[Bf$�(�r+T����ԇ�ZG?s����{�ޥ���5��47���xk�:����i�.I3Dm�Խ�0s����T��8v����-"�����]P��$f$G�-]�)m�S{����C��W��w��#|�;rXoB���0�G
�BAN��=6�s�p80����$�d83np�N2�wIQ�+����G�|/&���~3����;�
n��@����\0����ZŔ��4�eݳ��Nߣ��B�U�#z3�k�TK�{vFF������ �~���L`��E�R��0�&����f�,�ݥ(4,I���}R|�m��P>��7�l��lLU"=K�k��[Mb���Ml~�ݺ��d�z�)ZI�#�z���&��~r�~�Ö�O�w��2��ͨ�jV��� 
�}�������g�~}��Y�����$(��ᰗ@ �⎂�=��$��!@P�������Ǡ�FY�? TO4C�Xv����C�3�d.����ԋ�'��s�r��V���D-vC|4�=7���j���w�'ߥR3�:��[���O�KꞸ�?��$)��2���'��Q�+�_�]u{Z3�Y���Ѧ��H�"�T�	N�G���͈��c��8}�(RAv�����"���3a��#f�sh�+�.�G���t�U��"�@gln����Woe��46A��>'ö!��+�٤�ަ� ��8��󴘠�k|��1��NZxX���F�=K��-̲��a�T�������� �u�Eθ�E?I���|����lV�*��/����.cp�{��8,bU&���oF������Iʮ}��{����%��_.�#���;mN����>��2��J_��Hγu&�k�� ���Jt���{��)�	N�\w��˅4�d��2�,��F"�YC���+�e�KU�L��F_��G����b1��;(8�=��� ��޶��kg�Lg�P2�üe���e�E��l6���ߊ�����6Qy&|W7r2��ʯAU��ޢR�.^�JȂ i(Í�����+��x*-DD�w��_��هx��}�:Z*��)^��N#8yE��A�`���Θ��&$�����������ߕ��q��F�^�l�/ ��g��}A�5{��#�Z�@�H�UBW!^��S�vA�⓪^^��߆�l���~pֳ���|iZ���	֫>�a*��t���)F��3��44Cx�_�Ԏ�ɉ*��(��;� v��$)������Y�E�P��z�ẋ<[|�4o�	/!�����i_0��UT��:l�@Dʘ{2�����a�<�)ex�+ ��J����.�u��I��=��S��ԑ�%k	�p��)@#��B���4xI����ů� ߏ�O����$����;��U[6�M����'�'s�%�~���N����^�|C�t�_�R#w�>�*B�|oh6)� �_��AԜ`��2T�_r�9f��bs���Nd�� =|ȝ�0�B �v�<�X��,l����bZ���{;�^��|�+�b�3N�o�!����U$&�@H$&\7d�%����}�褻�lpR�C�ۑ������Ji��y<~��&u�)ڵ&�p���G�Ş�1�/슆ܝǷi��!Ai���؂ $mKV��=���z#�]��\���+�݄R�8R��_��,c�)��I�F�d ������fPhĭ0��Z뚫�c'>��7�!{W��]��L]�*	uǌ[��
2�B�]���ʐ:aG�sԌ����(Ӣ/*D��(��D]z�SC�M.yA<' }�[�����
��zT8��s�*��Ol`N��Q�__dDf�iC)˘ۿ��� ����wB��dg��Ay3,)F(�gn�WrJ�w����`�����h�
��m$m��'l �����=�#�F�0#�h���&<�Bǉ���/K`L�����fi���+죱4����Qc߿R�^�b�I;��nѶr_�z)��7�8����#T�O6�N�|����ĉ�U���^�)�%�]W�R>�hl�7>ݽ3�6��x��Z-��q���^N���K������x��D�=�&X̆��Q���R�5(�c�'�􇊔LR�W�J)���G��Eq���P6�C�����(���O�Y�y'n*UK����R�P�~b�p��!�`e���������1,��J�Ę(���t���*��y���"��oru5��(5���ddg 4���o�c��
�Ǟ���C�����m$�I�c�������8��\��,�G��Wf��)Sy��8�Xc�%��}��σ'�b�*;C�6���I���_{~�����Ŧ�f�Q<<�����8����	/C^�E����n�ˢ|�g�������8������Y�T���2��\a���U1Z�9��FB��]	�y]��gh~����a���֨vw&]��aD����@=�<�[c������!@�_P��ފg���Z]6o~p iWˈ��3��K;�m�T� 	�_�9�.�Kε�~ �#yJ����ն��=�s��/�R��9��n�5�m����ˁR�4c��f����_o7��Z���&�Mc�ā����'Z��E����fH���i�<�2��v�T�������^��WM�[&
�_����Y(�G�i��;�SpCR�WR�p�0:��{|�9R�H$�����T�N dP�7��֚��e?-�\���h�]��5w�d^Qn��rB�"{�d
�q�������|F��t4i=ȳ��=�Ⰲ�\�J��(븳u\�+�(WQGXu�i%y�����&��Ĺ�k�9yʕP±8�EXl=y����d�.%�2#�-�RMX1��
�7 $2�Xs���X�����7��+o"�0�Ap�6¯�������6c�d}w�{��*="���6�ŏb�t�V����\�/�#O0#��+�{��|Ux�U�~���+N��1k?��_�D?p��m@H��I�cR�&|p�7\��:4�G�3�A��d��ڳ�G�v��$3�AF� j{�������ε�_�ZƲ8?f\#��Av�11^�<@`l��\��c�M�/��&�b�t����U1h�+C윸:�W�u���,q��(���K�oVyBeODG�^W(�֘4���j1�xB7b~'�E��u~(������H���?8��H"L�#��-�C+��ՎbdR;�4\��}�������J�6ԏ����j��bE�w����tv7��$�� :B� �WH��Cq3M9����6�)^f�S�^�VoY���!��y��ty�̣���
�|�6�&J��n8��lq�D�7&�.�Pe�T�eҰ�P�'_X�!�u�@� ���}��
붬(n�P����n[C��+��醣�5\�l�DB�|1KT�ܹ����Óݸ�Uq֮�X,�Hk�a�������QQ�ʕt*4iSW`[��!����N�_���w�I󢤰Jf���q�m
��mo��mb��G��?L�RB4�f(,�&J�u�C?vg��w�q�UJ�Y�7Yw$�r0$T�����a�>_�ȶΘj����;V<֊���r�[>����A���lV]W��c?e��k|��kzd��6�ɱ�G�R�����Ⱦ�f�[R�_ǽ"�����T�h �7��)q�x�+D��S���dzDwQ(A��
{�Wb�c]�)�ـ~�q8ȣ����B��(mX�`i���&zu�Pi��� qF�c���jȏFzo�n	�̄/�Ìaz�B�l �,�Y���������^/�8@TFط<U��*f�o�,d�S��=�AR�O��7;�윋�	/��3��ْj�j`BZ	ߑ58W�
w���"�Z��~�BG��+{�'_Ά��+� G��qx��k����K��ࣞ�i̛�+�:����D����כ�L�+�$F�/�N�1",�I�8?����)������.� ��?�!�z�;)�w�wہO#MX�����E�EwKnZ�P;?��8Zs��ܬ�Vx��hn�e����/���gbL`���~t�Lz��*q�}n�<?�k (oo�����q����u\P�2��M�^��u��[Z�����v�9���Zm_�)?�x������1%���7��^���ҮP_��3U��
JTϲ=��ݓř��gy�K���ޥ�e��OC��A'r��8�����%��;Y?���}�����.�te~?������gA^�FS����>[�ꉻ���)n}���).���f�2B[�D���9�g�Q���᪤w:{�~�Ԑ&QL����z�#��Ώ����*)�����/�3�5�(��dQ��F�����C�<��K�\��Qàɓ��5B��)�nt��2F�jX�`h&�v����if�LՀ�4X���RǨe%պ�vƩt��y�J<�����Jg��s�m��씘��������%S��5�����h�Yg���Ф]6��*��<�!�,�9����w�<�i�w�$�q� ���(J���c�o��N�焏BD������!̨�/8�;WS���ç���9Э�d�&����h�WU�LѢ��'U�1�Ŕ\�07���!/���qk7��R��Bܩ��iD���U����^3�uc��q��uH����*�a�bݤ��W��a3�R�l������!G墆/Z����������I�J��lT�k��g��^ZP1]�����C��IQ��mzG���v4Ԩ��S�bt�1r�:-�w>;���r�j,�y�)��Sc�T�