��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_����m�e"kxu�Uٲ"#oB2�-g�j��h�p� M T�(�P�+M��&�[���+�=�n9" �2)g�ݕ����r��J)�a��m$�ke�xT+�ol֘B���zUz��}�+F�v�yC�V�`�W�#ƚ����?��J%!�i+���5�����5!���o0ٳiBk�욃�ٕt=R��bZ�r�85�W�\n
�*�Guu9��>]X������˄��?��]������[����.m�5>	^�ٷ�����<����߼�PU��0?���! TC���ֹ�0#�t,?��uNE~�w�qH?��C�]��?��٦<'�<�����o.������lE�e{fQ$���(N��0E~�ԗ{q�9k��Q�G�&c1�掆]�p�@��=?�هq�#V��H�Fz��wP�WMe.V�.Hi�۔zw$2��d�'�U�zC��V&MI������$�=	YL��w6D�OX2YW������'8��=��n��>�6� ����v6��c�E:��h�a�ǃHT�<����;����Q�8�<�������4��S���A�t���+�A1|C�W��_�t�i|/(",������B2GV���P6�䎛י���Q�!©� 3��''�dz�Q}���"���^w��Dn(P�X��֕Phһ����m��l���f�Fb�T[���2����U���~�+|��+�&0�h���_)�~8msr��뒈��`�k.�Ϯ�V�<b��%�5�)*������f�HsZsx>D���~��;E]� ��/��<f�%r�׮���8J�6E-�Y���k�nl5�\Ec�N��ҩ���(�?L���b�b�d��=��zqE�>�B��Ƒ4Fs��P�bq΀��6��!����w��PG�^أ���"�U���R�N�?��J"�߮h���H�cFE= ���@�ylz����|�kޘ�8n�-��H�?zy��`�f̬���w��"nvF�H�"�uL��ud/�yc8�k��]Up�e#��o�`c商ς�������Ь�bR�r�z7b8B\�A�R�l�'��|�T��@�� ��,�SKC6I��j
q�l9���$� :��#�}�
�����k�3):]����Xi{�X�o�>�:�ޔbT��YwxG?�I�{�A�ԧ����r�!����xn�]AfQ���f��9��HK<��o܆�<���͔�:!5�Z�V5�~Sy�4GLk��a"����;��9��xeܾ9{�](����߱����u�t�F�O�XS�B�f}��	�@L8�Z�t���4Z�x6�Ὺ��P48�`�(:�O�̂��W4�%\�\�=�QfS+���^���ujEM;���h�n-��0��#])5x�	"�����z`�G^캂�Z�4�r��p�>#�#Jҿ�����������01�0�v�� �/eny�ө�ҏ�� ��)�R�u8i;��%��X�p�N���]\G��*�6���B	J���r�H���x��X��Sַ�<c�д-�g�N�=�x����/�U���m�N��\�q��T	'��:��	x��a)1b��t��c��,\�R���:��S��i[I(���a@�S�J�I��?�wߚ�	���V�U����aK!q��4�U@���u�a�7�ٻ.D|�6;3����*/Z����	@T$2�<zcl��B�t�D��U]ؤ����eFy~Јs�}�W�3е�CK��3C�~��]C�K4�>Uz��*}�/��ށ>>�� �$��&�ג8V~��R��W�p��^���h^���t��h� ��:+� 61@A���g6�sFF�`vsJ;i���U����Y��4�6�O���=C��eR�j0�[�`8�C�VAX: k����&��-a_5�U��c���$�H�J��6��f������ʌ1!6��2�n���s�+�  .߆Ư.��N#Ȉy7����(��/��!<����%)Ըf�`ޓBV���	�S����d���h��m-랥�u
���%m�Im�	�ݞ�MP�Ƿ&��|S�#�{��̔p}qs�^�_���:L��H��nD�1w��Z��Y⡙� 쵃�Ǡ$�����5��Cp�8�י��gh�0�&\DtkQ������,�rx�5B��+��������_0