��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�"��F9s�`&���a�oq���F�g�O�]�<ݲ����eCL��D���{�5��8̝DFI��Zp\m|Q��
�}�6C���UnF:<�jΈ�2�����<����sf�k��,jڙ�����2��X��Ss�HL��	�������+g?���N�Ż�����|�v7�{M��VNB
��Rs�゙�Ld\��X�'��R :�J���^�����kMkx�Q���3!P}�e���Z�Y?.�U{�RP	�)��lI{tI(S
7ZF7��R:]��Ѥ�>aE�+``غ����%E_;��p�H�9�`��A�g�(V�����oI=�H���$���u�5�q�
�f?嘜U��u���K�P_���57��m�4�m��̷h���ߎ����i�&��O���8�.U�����B�7���N���S�q8Ks{��T
9`p��� ��a��މ��/�띳�����sU����鞓��d��O���Hƹ*�R�a����85��Q2�\�iXf�vh��U#8��f�[��K��ˉ�����@��G/���j��f��r��]m(�λ�="F��x�������M8X�,��R��ԑ;P�D�qΕ�P���Jd�6q��C���V$��(��of1}���Oj���"�f�ך�>b�5�6�R��
L�~~eP�U�mP��^f��(Ϫ$�����O�6��[�. ���\Dd�]*S=C�.���0)����DY��]-���UcQ�gq�ɟ��i�����h��)*�C���̬��� �m�v8�k��oF]�Ma�E���@-P�T�5����b�M���=˓��Q<��Y �<�p�b���2,}�������t���%��A������7�w���V7���6��&�x�7]'�n�$�����E���t�g�ui4a/�e/vg}9́�:�}s�*U9 |�|sT��*}��ұ,>7+�,�&��B�`У�c��^��\�*�
{����O�/9��a�
�.�HW<��!�m�'�>�)>vq"��0oz[c��N]���c� ߫uF��r�J�
��J���+��^���*a���|O�����-���x���V_�w��0T�0�E Y��
��"(�Di� �s�(t��W�r��>��5�Ќ�2�ݔQ�:X9��d#Ŋ�$���dC�A��ڮ����!�fe��w�ɥ��r�����JԾ���s��'W���R�N�(۪�H��vp._�O�.!Щe�A�6o��X��ҲWC�oiqS�,���ő{7Ԏ8�50.��G��~l�8�ڃ><��_�xm�.xvN:��-��ۉ����
w�n<`�ee���A��ׯ����El��J3Sԍ��c��'u�����z�yj���
t.Җ-��+�>x�$םl{z;|ޠ�,
ύU���)�㌯i��I
�^��$Y���4k�!Z�W�Ͷȥ�«X��0�֒xaXG�l��_�����x<�'�;59��#��m�_7P��g�zI�ח"R�o%�ԕؒ�9I��xL$�wo��7ٸ��:�.=_�x�P��6������ǐ�D�i�<n��/��<�����C�,V?NK��^0���5Ց:08�V�r���z�����ź����>g�V019y��_��}��h?�k�~������3��x�ʉR>�J ��Q�7�9i���\�E��T���3?�e��M\��6�j,�R�x�> �5����)�D=B�n?̝��Xb�����ﲉ��;1v�1f���`�%�()���x/ �^�;ƽ�z�U�}t;�w��1e���P�P��K�`R�I狵�7s����ʩ�F�S��]G��$X>��X3��c�sH�0�H:u8�{���.�.�`	4A��	�K��J��b l���S�����C�Thk^��
Tj������.̼m�6�`��cv�-��߽_�d_9����3E�TiX��L,�����-2N�$v"*a���xn|��N�[Z��ͯ�HK@����Y�>�b��=�r�Us'?`�Ei�R�n���X����k,�s��/Ƀ�-:;���1_z�Ӣ���� �&i����2ua�Ş3į�hð> 1�mm�90W0��SZ�puP�2/궪 �.���U�1�z+�ۂ4�(�6r�[&�W���4�3M�&�H�g[��SP*�(P�@ZubPէt��K���}��S�Ə���a�g{|N�"��J[�O��9u �B~��������
w�^�?Q�!6Զ�㔬R2u$M�+v����X�OU�L �U9�o��"-������t�U��@Y�J�vj���mb��z-üM�a�����P6,k��y�x=���${��5k*8m�lQHMg���x�ȁ}U��gLۊF�����MR(�(y��E�_wg[�D���?G���,�|:f,KS�M�%�+3��~M���	�Ȗ+GZT� )�Z�v��z���u֓&�5��E���7�]�:���}���Y��*s���6��. ��H/�C�����L����BN��'�����x�g�k�ޚ��_���.���!����z���SE��
�2�Zl��������C3���ÈگG֏�����吨��5�_��I@(ķLaʗ�Sȏ���n�o*	�G��쉛��9���^p�Yo"o���)T�u�d;�n�'��\0�E���l�J}�N����X��:�0���D�#�K:���'}�9��Y�6sa.Xv�K=�7�Cw�xSL3*r�^r�kI+x[nj�"~����8Z�"�O���f���ê����Sąmlh7�M\\p�4����;&p�%�*��&E�&�8x��Lv"o�2x&�Z��pǼz�АY�\��QE6��8N箜��Zf�YI����'��x�ɛrX����-����\Ԧ�f,*�v����.�Mr��]����V�Qg]���y/!�o�î�Y_�K�A��h���v���~���2�VWu@'9�+�,�h�|��碑�֯�ߪ����fm�'�3nߡ��������NF�f��[Xq4�;�,y�ߣ��s������[M����-:|A4:�d�����H�[����r
���hg3
���.�wY?"~)d��㪘�1(T~
�E1ðlr�Y�T�8=���Ъ�G��#j>�hV3-�2����":��,G
ر���(����ܶ�N�.S�(�L�;b�T�Y�Z��F蕂�y�:$�֒{�$�S'��k=L�E.E�ir+<����ҚUe! ��T��g�U�-����6u���������?���-��|���[��`��x�* ��j#�ӟ��~HU�j�p��^`'`%�+��
?fԗQZe�',�o��ұK��x������M|6mK�	�e{O�uRy�0�����f�������7i���¤I܏.�j̫�1v� �$��au{^��

�w�MU�����n�}��Q�9���~F/tx�?�Y��F�u��ݖ��� �g��3J5�bg0H�Z�Ʊ{7f��cW.ͤ��o|s��� կ,� �{8X���q9.�����c�?��L�A���_j��b�r>�+���ШѠ�3r]F���t��S�`7�i�Q!�I����)���T本�{�d)�Av8�?�_+��oN�L �������U����qJ�����9����/�6�˟�nAN2E�p%��ݙe���vG"��8�RH�R�~���A>��Lb�\v�tX�!o��*��$�Rb27�pe�}���'����x�ԣ9�矉H��	V�ء�^��p���٭T|�˺�n�6��د{p�G5|SL�m/��݅M+�O<��xajf~��6�Q�~��qʃ�ֻꂔ,q\*���1p�ܭ[��%mԽ�.��n�w@���_�΍`�n�=�Χ��i����v#*�H<��ii��?% ��/Xa�hS�w �0�@0�(�,N}�7�X���L�3�l�HMB'�A�W�R�;��h� `��J
��K\0)�fMF�ވ6��5��(p+yl/[Uk��8�L�Z)s�ϛ! �[������q'jT!�����h�~&_t�K��#�5=xb�M�
��xL�y���"�vp���ь�Ž�_ �����y�ǩqF��Y�^7��V��<��JW�0���)�e�-nR��bXB��ⵯ���n��B�#�6��$��H���b,�޶�e�!��u�"K��z�����0ˇu4��Fk9�q�5���ƻ��[�΅m��*k��;��Y�\)*
����P�t���4Dq�V��	d~=�Z�rn�����签��'��wϥ�����5"�������n�LI��bd�і$���d5Md�9m��f����k��}��g�9:��=�+�(m�*6h G=��&ښ6�4�f\J`^��EJsJ��?�=��r�Q�pګ���L]'
�+�yew�:nE�;�w@G�,ʹ�5���E��.��7/�$��ʾ�J��S��(1�M�Z�D��^2�fd��2ꂙ�P�=Od2@�\��+y�W?[�A"C�6�>ݳ��4=�\K��	g�C���j};6[af��G�/��!��۞ګ���vy����ӏ���\�iK�sE �0�����G:d�
3��4���:T&���:��(Z2�������(�L�2�HE>���馎q��M�7>�*D��xiV �c�\�Ƃ���C�x���-ޘ����K2�e�_��f-~� ���2�>-��Խg�j8[o��g
��c�3�f���|�iUv�3_�x���Y�5������V!q!m&�Z#iw	G�y�!��յY��񺋵v�ᓔ����$\3]1؊&l�]�}?v^=O�j̺sa{nf]\�J��A��2ď��c-�&���#!Y��a���rG]=��v�K����rY<3��{�!�H�jg�^�_�-�z$�N����+�Y$�M�ԅ�*�e��)��J��ѹ���c�v^�����+D�:T/L�@i>�����sÈ��W/�c5��u���e�ϡ�S�����͊��G~3�k�k�wt�p#Кʴ2 ��R1���zР$/�N���J�b7K~82o:7:~_��r	�<�
~W-����5O}&Yp��%`�)��WWd��k	/���:�v0�*��ֿ'���ya=�)^Y��#���]�H�kн�V"Y�LG�Gv��aĩH��%�o�39j�����W��"
s��t���\��Y�~4u�D4��E�Ý�O��l�uN�Y	c���j�+1ǍO�#X`�s��%�?_~R3��8;ƻg�'����RT��ᕞHoK�QsS���I4��`e�y���֯� a����H�'��H��K<�bTSgT�E��Kj5bD��A%fA�_�����#��$:�#�Io����_�5h�{n��8�
Z�L�9G?�mA�=/w��so��\�T$[�acRq���'�ӹ�����h��9�0�_�z�c��l�Gb����������-!.�w�v�(�����y?���0k5�*e������� �|����Su�`�م�Y�x���/�7F!�Eya��ؔ��$�a"7>����BlNໞt���1�N��_h�jNi�֨��}�
�{�wL�(W���*[�0����
R�~���� �B�$>T�I	_ir���YX5��̶㥚�[��B+���Or)���Ƽ�h��4��@���?Ƕ�ެ�i޵�Ǒ9^�F��L��iM����6s���e��.�����0Ai�d|X��n�7-C��gZ��9=:�O�0q&.{�A=D/U`/&mZKhx?H���Z.����	_H$�݅�������%��z�ӂ
̔њ8�|t�^�ZA�U�.p�1�P��%oςB�&F{�L����N��݌���c�'#A��g�þ�7Z��5����E� �j�9_�� 0:�.�N�z<,���Βm��{��d`�&��:�=�ze�����ռ#jy�����I���H����3����v��Ҫ^~6��5l:�J�A𠄛��vXP����m#���1�F���`5��!Sb�(�'�~�]�נ�/F�p�ɇ]z4�X��6q$�9��)U�=zM1S��C�?l1�X�jG�Wc��k����ճUt[sPc��S��Em�p߽�l�j]�ʰ���֍�����V��J����2�gf]��5ڏ/Ƿ�+,%~حj��K�SF�-��u*�6�2Os]��p.�۹oi��O�uǙ|�zN��p���9wfv=�;�s	=�k���Xh=xU�P&��
�O�uȉ�V�`&�mߔ�}Qނ�����K鳔���R�����?����̺WN���c�B��D�$i#ssq�8��V�^.iF"�tbbm����(A�7~�4"c��<nA����Ա�c�����Hl�X�h�
����AdQt)j��?2�t�}��p1NZ��Ӭ���G-(O�[ �y��y�t��\���r�0q�$(�ɣ��`^%/�������%�{y���~���D�_������>h��(0�ƪu��MU
L�&D<��Y���Tuk� h/)��{T]�@���;:���]�rG�C_SK��B�|o����H[���;q�m_�g�`yU�U���>���r��_&��1��b��Fʱ���d�4�-l����H���3��,6u�蠠���<��M����^�*��� ��j��Z�nE���v0F�#�X��]�e��P��H�˸>;g+�D�$V���豀Ygw�!�e ���Uh~���oZq����nތ�^�(b<�s�3���b^H���H�8s�����;Ҁ[s5ڥƛ*��GjGpuݢ�ʍm��>��Wn+��#���^
�����-�^�nu�^��?�2���m�pw0�5�[sP�A[�ur�pfG$��d;���S���1����Ԟ�@]i�pա�\G�=}��P;]��onݐw��;j�ϗ��ۮ~���{E���(�GW��$
��S�i���,�掔���nV�t]�~�`b�D	�,�aERS;�g�ç�_c'j�`#�)hdtA�WR0���O���>|�v6dhf�~��zc��п���JF����f���"D��z�=��*,��۶)1~�}3L9��2����
9w@�IЁ��*����KSy�HA���$J�T�Z���a�!9SR����2et��1��.SMsc0�!���ʑ5��^̲��<&�����ת�3gp���@w�ަE�K���5��p���q��B=�w>E�:5����e.�1�;`��C[]��Iu�r$&>����if�S�t�h�gK_�V"���՗nR�}6wb$�"�x_�缷(�*7����d��S�!�Z;���;�4���I|Jq����,�O��M�E�L�����k�3���G�:)T>F.r��J�r��$���[�u������b`8�@�0�a��[��=S�j����P��#�l� C�I> +#��