��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|e����M`p��L}a�1���mq�ݭ
�:ث+�n���M�B��7�jŽ+�"��Kk��։`��X�z�1�i��J���e��4Z5���C�&�⒇L��禭�c.Ę���\��9�^�+����Ƈ!6A����`2����<^���4E���l���V��W�����.��`3��ϴbg��R.���,-k���*;�pͽ�̀XjD�tn�lt��f:�s)ĉ���Nk�����?I�B����x�O�zhe3�!�ZO�x����\ ���63�c#��~6w���vG�B�W��	H�8=B���Jg��^���Yf�h_���`���-���)��P/�X�u�Q,�ᦫX �op�g�Z��؂"��	K\�D�������lJ�n�#׹9�f.�m�~��0�V��i�=ֈ "�4�����;�o�%��_j����KC���-PT��`wl��֯��"�f9�}n�N�z��U��cqIAğھ���{�{����|.E0}I�a��Em�A�i�Q�����5�����\xq�uAt�p�V9%*~XΒG�"੉�����,&������N�=W˯ �.zo��5�&g���ª�B�I�0��o#���60� ��꽰[b��u��E�`�! ���\�a���{]�!��,�e�Z+TVw)�$I�2N�S�5�|A%6X7�M��� �1I�ݒ0W�@6�|P��x=Hz���UY��{���N������NQ���P��f���a)3^3��� |/94'.I�P:��m�ϵq��`������<=�D7�ny������e�?{�>�u-	sg��$������QY��&�u�Dw#��8��]+ ��_x�S��#�
3�JHYPR�,D���������{�˖0C=��^c�<OM����q��P�Uu���'"F�Tev��UG�e�d��R����/�
�i�r���`N���\��{�Rx�?	��k�#�������yl=R�=�ݤ��x<M���nZօ�rN�3G��uB���K9^�����r$GBj��![�{g���uv�5�3��X˙
��좤 l��UY� )�y��t΀	�	�j���#�8�?b�֪�i.8>C��J�(�f!]'��4]��U����E���8��L�>E-������/�A��)Si���5{gL��^U�C5xH�̈v�r�'޸�"�)W!e�'e��V�s��P
��7��H�J2�\����z.v���ߴ�U3'�n�r���=.�f%F��+����i����\�=�� ���f����#�� ��=���!�y���I��G�%E󫙯ykzd�;-�q_�%2�~E�x� �ZjXlN�7^o�iQ�N��i�C��R�k��N�D�=e3�t������Y�y!�3�#��e��\#8�\<s�ԌoQ�`e�X�����¥K����{c� ̾^��2�^�&�LE\�I�'P��I�N8�OY��<M��{;��DB�NOkV�SX}��G���.ӯ�y"͡�D������p /�_ ��A��o�B�zN^��:O��S9~X*����H��;=��}�H�� sh�}����^���v-Y^�c����+�;70�	N�p5�`��ګk_5Z�/�s`lF���w֋ж�Fl���+�4���D(u+O�hg�x�ǍI���6~A#z���^�
�o���g�V��k�����D�]����=ƣN�c:+td3FY���8z����H8�x�^,�nT��Z4cZ�a����#������EUDL4�
���y�d�8�Q�<�N�ZԽ�ù(�8R�ru��
�jЦ&_^��k�K�V�&�:FE���$F�8�?�"}��PY>���f#hX\�5���#y���qn#4�q��s�b��Nn� );3�O�ĺu�IU�f�Q��[o�O>�巋����O=�횅J�|����tq~#�<��c,�"�䎽)�/2r:��X��O͵D8���if�N�Z���}��fx�"��y,<�,�KSw��%���*'��=��g.�P��:���{����ͼ�݁�HU�:@"�VI+�xR�������"�v��$��go�>���H!A�@�ר.}mbs�oe���v��'qeX�υ��#�U`�W0�Q�(�U�D�����CO�?�1�C.I}�L�D(��PmOu>��K.d؇4åe�1lA�������������=�k�W4D��f-V����󁽹p ��i�*#Z�� W���q��o1-l'�c�XZ]c�R\h���ó�IE��X}��C���M�laL�m0ןlT���wfQGj��>5��|1���T��(k�E4ڴ�#��>�4�[�2��V%8�Э"�< B�gu��Rq�:k�P����M��;ؤ~y�����虎�l�PӸ)�LU�eģ�Ѓw�����d�Wqu��eA���p�I*�`;l�I��7\�L*�$4���!�j�R���m�X�»�Gɗ�H���W�!vpq�̿���.cJu,
�h4�Õ�%�}��g��pm�|�8_<��at�ܜӎ��� ]˚�����k6�"R�`�ɖ@�}�d�-0�c�Q�(�>/��3$�cc_\)��k�d��`��ۯ-a�2��`��Z]z4�vK�R��J��
?bŻQK���U��*۸pt���`� U���[�6����1Be����$yQ
��@�e}�b��u����!�߲߱�E�	DJW��P���K+�}p��xE�%���9����E_BWS�Ԯu��T��;����(�j�RxZ�m�l�׷?K�Z8��ec����8�5��Й��v��\0!�;A��+Fv�x��m����x��O�/(�@��c߿a�&Oǜy5,��S5�'��G_�h��j��"�G�0��-����:��>�sQ����ڭ�t{��oGW݃g5/r����U����77	��׃4�����@Fϩ�{~?�UbHI�� /$΃A��v@��e�A��!����&�<�ۖ��0��AVl���exRVao͟3�Fg׬'u7<�m!���uW�K�}����]<�ڶs=�c�خ�O���y]�aD�D\��������.��Y󞕚oglX��J�iL8e^z>�B:�+���4���Ch�6�)�Fhu=_�z:W+	lW��O1B�g��_�.n�||����M���()����]�j�}�RI�4�b4�� M&�쾑��`� E�'���xO��,]���|Qmr����l�1AQ�#�B"yA��,�[z滲���x�l��`v=5�����@S,H�M�K����e��SB�v2�{����~y|(�Rw���<�p�Ao ъ����c�(~�[���%j�Jdr�\Ζ��k��Fy�K��f?���i���s{j[/�8L��{��<��>�L�$���ގn��R
�4�\Vyoڐ����+}�5:X.1����]��"�����E���tIɫ��u2xu�w�T,�]l�#
ygI�؅�m���	^��L2����%�n���7�w���b@=��h
tA�z_+#vD\�,�	���v�088��V���X*��(@���Ĥ]V���M� (oĨ7r���ۀ����� �yBeUZ/(�^������� Ϻ�֣J�K�L9v����Mr�����%b�#����!$�s]���h#�޾����JE�L̔o�oOd��a��<�
E 7N���R��-��f>��p0cr����m����z)^)H�	ێ�L6�B[�-�D�QK������B/Q������0\:�X��rv�{���N���ic>�M�N�_m���~{%s���e=J�D��C^19*-[�`���U%�^pHzǄZ����I�O��(�<��0���z���LH.���<�ԵQa���v=?Nag%�hN[*�h��1�`��J�+b�੧5���B�Dt�,M�\��蝇��80����
�����D����z� /���aPw��/�~�_��qZQ �U?LF���Ӛ�����R���;n�]�0[&�o��ΫW� ܓ�1Y�X-ߥO��������݃�7p��Z�*�L��f ����`q��l��3���J�sj�=T8����3#���p�eK�PA����]~��b���x^0»�u˟e��	g��0��;�.�{ȿs�Ĳ��O���!���}���~O�ˬ���T�V=B�k�u�=U�=R����f��p�u�+}�/�{ʑ����_����Ɲ_A�\��(E*=uݩc��W*��Sk2��5xR�qQ��I�>�n�� 2�*8�(�Z+Y��/�tތ�?���d�m���f�8��U,�}E��"B_�d���`�6q��ˮ.)��-���ڶ��e��D�#�@M�XLd�1'c�9s��TA�iX������ȓ��h�L*�#«9l���C,-$ �<�WXr�-�!�����d|�q��д[�hջ����f_���2� HY���y;gG��%vp��]�oj�ژ�SY���Å�7��Jǖ�,���^f��zU(��pL�:p����%�GN�V��P��c����)�|�>#�E7�DP6�ڦF[x��~��-Uf���*���t�Κ�Lr�8����}���BU�>=�K�<�0H�v�T~4� �m�Q�2�L�p��%@���ŔƑ#t�� {�b0-W1�
.3�cf�+/�3�Z�8�K��ߘ�{KAF�\�N3z-�!�!0�����'|�O�������Hg}1�^/��d�s��veb����L/�����sKu������h����br̴X��8!?8�ܖ�;۳���چ�EFE�΍�D]�a�Xm����4]e���c�MGv��d-��Du^�e��6��,�$z�ᴑ����qx��vf�?���Th�����ޜO���������"���&;�xa����X�� `�Gb��a��s��TG�LC'��8��-]���,A�ܚ�w�=v�A�	�8$`�p݇�~eXN��r7h8�3u:��s��H6kO"8$O4IX�G�N�[K��%�_�-�f4�sH�L=r�5W��IE�c��O���c��;��:�k��^��"'!*I�!�� `�	��$�0<0a�1B��K���(�F�����PM�.|n���7õ&�5���rMw�'N�K��|ojɷ�.6l�lw���1ݭsD2
-��Q E�'�xaY���I���(��`=xߝ�z|ߠ�����v��Me���_�/d�r05<���F�U	�8j����'�գR�-+X[�m���̝�_0h"��=�c���G<cR�K�t�*J�N���4+O�������jI�v�y*�F�w��g �I�`�3:�&��]6uk'�<����~KM���<��}X5�#���������6�����j�ey@��}�k��'*�\@����?���PS��f�P�'-&�R8�c>��Q������jg�|��@�cM$�/=�`�s��O�x��L��w+�}IM�q����+����J���C{a�i�g%�I�h7�mQgKh��Ұ.�(%�kz��Hc�����^�y����}(U��B��.��Tzo��.y➍��AƒKE�Ve��2l��Tq���{Ny��h�WZ1	���G�|���C ̓�a����Gv�Ǩ�E0��q�V���/I7����,\9:�l��fj��"fd��ɑ9�I�3I�j���Sۀ�&����y!]VXx��&zG�:�y���45��N	|B��v7*�m D��r*�@gL=<�I����T812�n��e��5��qG���RP��,���gCیU/��S��A.�m]`rw!E��M�<��i��;��X�hq8�`��Td�]��4��/�툦?����8+��j�US���z�hMx�W���{0�e��*P������~�r�C\���8�LO���o�5By��c���V�6�2�٢`��H���MU���M��ī9����?|l4�l�J��/A�����a��;4��
R��C�4�+b
G���N��bIyH�o~C �˓^�8c|�)X���j�����Ɉ[o_���#�<�9�+�g6��]з��6҄�7�q�~�q���%��f��,�����^���u��F�T�:��)VZ�! H/*��a�
�8�p�����#�����l����u�TX��}
ܙc��ˀ=-��FP�P0�S�4���!49�7/�ڼ�]�U���@7,;��m��P���u��L�?x�O,�>h�z�5�#mm���\�=��&c\ e0z��Tˁ�Y�F��f�����DMV������u ��������f�݅˘�%�+�l~�M}�M��WR����~��֏��?F�����,z�^W�����������$���qe~��.�}�e�Sl��y�]{��G�Q+w�&�OE��6�+�U�7:66٭�9dgsf.��'��t:�H7_0ó��_fO�2r�f���Ү�3痙͘��>��A����n���QY ��x�v��Lb��~!�H�K��W	�	�@P�'�Q���%؝=V���.���C�@g�x������5�w�uR����,�,ԇ&W�$�W�I�gF�x����}>n�U�h��P�n� Gi2x)j���M�_\�٦��e�/�L�vc D~�/n��?�,Ll�%`Q��%� N�qϴ�#��ek{|݆W/�v�ٮ�A.����qӁ\�6J{�b1╷���/̦aג�������oQ`@ ��s)���b��C�z�O�X�"5��2I�`y=d���������oy�w<Yj�A�&;��4 8!��w�S�����M�/�'��J{Z{R݌y�d��#�'(<
D��"�:���>
������;Y�1f�D�������G��8�~�4h�n)X�{^v�*��9��t(H��5Z�k�:#Y���[o̶Ѫ���S�ۮ��.�@su9�?98�uRdk�(G�d3���
eT�w�l�Z[#��f�(I����e�gV�H��ҳ ?Ɠ��2����O)	��ya�S�-�«�a�d��$�p3���6�5�ˊ�N�q���� 22;�IS�G���1ȼ+ߴ�,l,1��Ћ���VmK�q���N��J+�,��x�I�j�=[�����l�m:k��A��a|�!��pGoWB#
l�J�g�x�,��[��n�#ې�b�*������c%��0��B����9[	�.�4��[Mn`�1���*P͔�wT��������b����5K�Fϼnd������eNp���X�o-}x'E��7}��o�U$I�c�y��;�/9b�5�'W�5�З-a΋������	��݃������pS�� :x,�?{�s�����{��T�;�*ǰ)��7{BsX6�|-F�lHX��������sɺi���Q6�̓����w}sf��|�u'7dͩ����K2�G�e�S�n�w�sz5'q��ߘ��L����)ΎJ���]K����r)2r&A��4S/�@C��9��R���	����0܀X���C��"|���kĭ��������oI¹�4knƦ�C���.y?8x��Y�#�LM���`�dDwGX�Ʈ�����������]�H��҇���'�M��Ee��xq%�$m&�_ȼ@(%�:��-�l&���ihL;�N�F.�[��%C�e�B��S�?��a�<;�Ҕ�2�&O������Y	��U{Ko��3�
q�ƶX_n���P�OKSͨ�1��'�^��v }��D�Sxe{��Z��� � 6ڌn_^���~�����
�I�o����վ�WEL���]ӷ��s=�\�n%cS��tq��9�W��s�{�x���!r{)t���R�G �`�4�ByN��u������W��pUcNs��5�,=a���Z�Qaé.$/\(��9���.���H�J��G�$~����}��9P�'�����JF'��$Ő:B�dkQ����
;Y)87��%��
�TZ�ZZ�:`��O&���~3x����e�~	�KO�ɻ�
��	����y`�Ђ2_�עN�#�G��Kf*ݞ+?�G�1�#|��o@,�݅�S,���$ԧ70O^R�����(��ݺ�!
���Et.�$�1X��]����:^D{_]&�I���B���xF�G����+�wOh��_m�������v_o1�W��2���.Z��&+��-�6&0�-Sѣ�r���Z5t3�O�Q�| ]��)����6��B�ӈL5��^�:{�{s��0Rr_(��<��1��3�g����0R�%�,��)��(��a&�f�ő�J�)eڼj����/z���;��Q�B��h�|�(�%*m�*�>I[]�#���`	jr��F�V�Ҷ$�L^�NJ溹:���2}A��*�%��b�ȟV&����F���1p���1��-&'�U�$|�.��W2ҫ{/U2���E�nu~�m�9�N�|��(����A��	�Z�k�OS8Am$�j��õnL{�F���*�I
JU0�3\Zo��b�9/��;E�(M+O�B���#3ɾ��:7@y��1�ܾ��(�Od&l�;��`]l�o�6�J*l���F��j�>z����Tƴ�D��r	����o�*F�����<�U����I"d�-�
:���i4�x���FO��C��'��b�D�3(=��4ʳ{���ڇL�ʂ:��%�_-?ޣ��zQ|q���H��R����$�}.�%0�U�ϋ�����(�Mz=����HIA} �j/�cȻ�\h�@��O?xO�]�J�*�Ⳕ�H�mG�+OkȞ·z��.��c���"�/r��Tj�},8���	�D�/M}!/E)H~q~������"�6�/��&dN�-���í��&$��0p��B|=�A<J$��1o)tA�B�'�Z�Ծ��V��_֘������>XO�ɸ-XY�pG��Fٰ�.����K�����/�4��(�-a�6Y��\��^!��V��# ����8S}�t?��"�f?���M�l����)a��;��uS�bD�P�K��u:f�o�ok����	��գ����4B��<)h�6\yny��XͳǟmW3&OH�R7�l�L&-�R���Z�w|c>��������T�D��`br���P8�c����$��!:$�5�_u��$��nZ������n�lE�15ƹ�c�5|���v۸�*S��<��3�<�Jgɣ#._g�'�!����g�J���\���j����	0���l�I��sX!���I�}���l�T�u�Ӆ��)�/MJ_�� K��8w��P6HY�C��q݋�&k��olsQ�
�
�~@����֯�����/��DZY;^>�Xɧ��������(}UBS���es݋�D\-�eO>qF�o���תK 2))Eg���R����{��^JCL'r�.�I6�SEzt��;���b��q�a��Ў��ޓ&qo3�������V���h0jnY`�qx>���\�꠾�T1y���;|RM|)�v$V�i�dj����,ԗ�6k�Ƅ2�T��М�Q= �WF��2�
Cx��+Y���+wr6̱��7S���!��|p|�"8��R!��i���G�`Bɫ}{��� ��\�7'1�~���l?}O�}*ά�}��[��K���T�t��g���v�;�	�$����IhZ^���e~kD���KoN�Q>�~����\�]�����&O���eC���S��{.�Ӝ�1�9r4y�g���|l��d
<�.�
kˆ�Z+�(��.4�XItIs/S�{��1(��t30w��,�% }�Q��b*"���UeJX-�Ff���~Ӵ6�R�?[_��@�F�ބH�ZO�C��	�qu�E4p����Ւ�~�<؇X�H����M�aR��{BCR)��,+��:��	�Z#�6B�LOC�=��#��0�}Aހ�on��LQA�Nu�'���չM��y�V�ZB_P���J�T��%6��4�-m��c9���w���CXW�	X#>ǔ�2M/	ʐ�߃F��(wk&�U#�i�ύHUȈ��c����$<A�z�2-�A>��\��ۛ�n�U"8�e~wi>���isS�*)��at��>:��<�ePU��*�^��Q}w*����iD1E��jf��T(D/-+�+�wՐ!�"� ?aѿ{"3[1��~�7F��«��近"f@���k�̯��s`��Q%���,*��/j�e:��O���МVJ*�D�j=�3{�#���Fet@���d��UrF��n�]�_eu||�O����!^�&����Q-�YWzUC���;�]������9e�rA������e,n(q��ߦ=�~�-bH�=�Z1���o%W5~+����hcj��5���}�7���˅b���Ma�Qѝ0�k��ה�!Y#�����Q��{������/V�Ȥ��鈬�|� <�>]6��b�.`�:�@T 0(7���4�k�l��0(ʌ�<��a�vc[o�	K���"F�L�j�NU��n��!��`Fĝ�`�{���(�ڏ�Kʄ�~t)��0�N�I�9��'��Y�!#���BD�,�{u���=j��(IP���\�-6Â?h�$���	��iX���u]0UP��_���Uro0M`F��'d�t��K=5@$�>�XS:���u�
�3�ǵ�����||��;�>^�m�%��g���5[:�h�q�!$�2��/O���d�	D�,Ú_��w���Ԁ烔hҒ�9}]����Z.���n��I�j�M��܊��}��2�U���JqR�O�h�)�@�6��erɩuDq�<�-
��:M�N�^vnj���Më|�9�o踔�r㕲�(��	�J�T? ���6��h�\U;����Cj(�H���4LN��6t���Z�S�G��.�?n�Nr��F0�Ce1���Z���+��ճ��z�ND΅��1�:yه�|o���A����n`��0!�������~EBQfS���if1�����Ē�79�a�D�;����莭�̿�M·�`�9�����:�
�32_s�M j�L��0�J��ʹ
-J��G��l�#Sl�K���'H_�Y=�ްkS\���-g�$�[)T!?��@��BU9�o�l��ia�LI������-s�,�wC�|4�{���Cq<Ύ�ehzf���6Z�^H������y���YL�ҩ��kς�R6O�\ǋӛ$�cJ�忿�����[��]Ĵ������|~f�ǫ�t ă�/֎��/-;����
�81&�����,�X���r��]m;z�*�הg���g�9W��:��u�w��o$��.���ȿ�x�9��6����s)�Y��sȒ��5�X*�w9N��eQ��$����F!bf1��y> �|�����ܹ��G#�%�.��U�&�����|z��LD�u�@
��T+&.X������`Hka>��ʩi\�E5|�U�6�ؼ�:�p�a�^�&�X��}��v���|�AM8���/n���9�D������nqɏ��������< x�ayt��&g�SxU�YI�8�QR}h������`_^f�T���d�r`ĵK�C~���g���a
���|���Y��I��196�N"�#���<���sKJ���C~��j���c���g7��r3+7�� UJVt��@$>����G��ʮ���kR:��q͢��"�λ^6'�oH��<��1�&{��3��9���[�]ᔌ�:��<�(8���^JӁ��31��$i[C
}� �Õ��	�����}�Z���8�7{=���{S.�l��������;HkI8�No���3�3p(y
<_Y�l�����0�x: #�l����r�5���v�9�gq�y�%��Br]�W!N�l��E�A�����M���e#��`X��`;R��R�ۛ��)%��J7�����#}ފ�KS���׭��2�<���2t#Cߏ�'GN�� I��R\�Gg%;�gbvq��ݰY�۹*d����Á���V��	ccpO�z~Db��7ub�qY~��m��0E�	�[X�<�e�G��DX�*�o��7��7.� iM���m:�p'������O=�F�ԏ�2W�\Tϡ�od|���˞��~�Z"��L`��N�%VV�{0_}1��gD�n»�*����5e�L=�k�
��8�����H2������*a�Љ����}�y�Y
�i�m�ߪ�o�oΟe�i�I)��΄��P��s����Lz��Un���Nml�QD��d��2:�v܅B��G��V�ȍO�a|V���O}/Ug�	pe6�`��u%K?���T���"v�Ưߩg��`�ʌ1�M�ciD�,�PN����4��@�w����IaD��u�'��@�K�\�����o-g�<&#c�r!�SA4� ׫�V��?%��W�j�u���|��99'i�֑�0@�N�&�)��J�8��`-����7T�� =�Ě7O�������g4�sU ��B��1Wd�y�_���3%ڧ*p�CڤX"E[�er��֦_��c'�ѡ��ʶ�`����*�3��,��[|���ig�V�'!p8�N�����_����x�#er�&*up'���X�*эF����vgd_���D]}�f[E`�����.�EC׳c5�3����(E�k�~l"��z�jA=θF�������n���$CD��#5W$qU��.I�j买r��
	�vjc�	`��=E�sP� ܛl�F�CQ�}��R�|�~v�!%��@��q�X����|�d�+�.פ~��L�`���V�z�ս�����O�VJ��	��޶'�'z�Jej�7�_E%�C7@���+��)�^�X��	á������8�v�R�#�Jvv2���#�֓���)][G��/?3�m":i�6��n��`���mqB �·ĢF���g��K���&좴ֹA�aI|�����N>�����1p���°g��,��+�[��@\!������L	y�Ja����Ȝ�a���e�ӓ)��	���#�����*�Wr� ����_��ug������L`t���nD챤�G�7ʠ�&��� �;.I�,Z�z6����G��_�[6r%�"n�T+w}# =|�<��t$c+ׅ��~əm���(t	��vK̍AI�HM����e�ۨ�['�`���A��fͺCWb�,�A��e'��-C���-�SY��'�3�Y5,* o��,*��N`���VZ#�s0� >[Y�wo���J��V@� fRZ����ob�_&�M�^����C���:���b׉;�1gc=D+���`)<f"�0c.���͙�xK�K��g4�[�T�ۖ<�dL߉��Kދq����Wذ�e�;�]�b���qG%��tV	K]�	R�r����!�u/8,>�f1�.W9��o�C�oա����#�$Q$�1��[\ָ��h��>�`�ѐ|�pr��s;�trP	[i=���<�śfV$���5�-?n�1:��� ���~ѼP/̨�@��m�M�WK9����d}5��B���'��Q�Z�%�%hy�M&�p;����)YJf��������T��g�<�~�U��Dj���NQ���84��E���MǱ/�H���Ȱ8�ÉHs;xɖ�lwN#�������i;���4"����5�sh҆*�lP�{:ypPw�]���@�[��	�*�3�� �AƷ���a���6���X<&&�F����D����KqY-���w%���sf�����3��%������)�
��b��l�x��Ym�̘�y�Z0S���d������H@L�<Qё���}Gf9t��������=u�H��m-jc���B��3F�kv=�V$�u�#�b��$���t�e]�S$�!n%�n�)X����Ho�b>��J��`�R��'��+`sA�>�l��/dH����W�
n�"�#���W��t�G���b�ib��32$ey�h+�@ČQc�T �]����o��=혵�|hl����fFY��k;(��jrITF"`v7����AC��'=[t�s=h1�Բ)C����h��Ȋ����jU
��f64Nb���j%�G��ɶ(CP�C����y��?a��H��xP�f�������c�MA�H��O��t��f#Y���dDH`{�qcW�L��a�	�u���C/ ��B�%ˊ=��}FfA]74��e��F}�y�� v��>��@�`3��w|4��q�j���ǍO��t�?U����<U4��k/����C�{t?x�6�h'����x�d��M"(���c%؄]\�y%5���]�Q��e��]��h���J��hq J	����u�O��/pG�+�s[��p.��|�X��1�S�jE��;�H�y�.�L�_�2��&,�4kx�A��GsU�����<DS�a��%|�xx�4�p !O�7:����
杹f�l��C��g�-�1Mi� M�h��vo�-�,���8w�k;��������,)Z��W��N)�&RF��5�"��,�� �~����^}�,���d�HF�|�H�5�#�����G�z,�9�V.������D3����h�
��$����cx�� ��~�7*�!�h�'^H5+UQ��|	�W%���M�t���u��.�W�a>K��� 2�%Ww�ך�	w�\ I�Q���B�`SV�!]i�f�`<���m3L��[���E3��Es�)4� [������]��^�X����$�'�∜�i4=��@�_Z�%ve��p�#���Dx$���a�3�q�73ly���S`�7��	S�ri52�TN��� �t�`d���@��t��8Az�U�`-C�D�	��0i��Jse���MdM�χ�;*�r�9�Z>�������C�x#��F.J*�X�F=�	���MrU�f�vL%��%ʴ(,
�A��j��@`����� _]���~vGk����F��t��҇5\D����-�g<���q'��Z~2���R���Fƍ��Q��r"V����w�?�컆r����ߏ,z�Kp;	v��9�|(��I�'�>n<�!�����R�/|��G��n:��a�Io�����ߵ�r�&����w=*ML�T���;Cj����]��P��Gz�6����
��<^#{�j'�YO�1���z�*��Љ$��U:�yJ�0�w�<5��<��s��|T2i���	��h�m��`w;���$>��V����G4�3��߾{�ՊnQ�a����XX����7�	<��/�^u�%�BP!
\��߮Y�|;�yIGڜ�sQ�Qp�j]�2��vm.U��eT���{�0��L�0]�	^j�:t���OI�6f_����}�7V�t�=W�U�MOr:'���Ö8����%��rU3`� �߆j�!�l'���rb6� �!�)��)��~,�>?+
Հ�j�a9�=m�S��ug�4�O�Y�'ݨD%�9-�����x_6�)���?qԺ�(az�>|[=D�O�����<�V�½�-����pY*v��W��6�9j���!:��JB��s�6j=r�1B�#���qE�R#z�`ƫ4 �,�:�
�iiY��0M�J�}y��s���2p����1�0�{�X�/��g+�����awE�$b�8Zr<�"H���>�p|4�.o�ݡM�xTbVuϸF��Gî�.}fWJ�W��w:AEg��󛣫Y�@������ˁL֥�S�
|���8ym�a�O�J��p���_��\��F�G|ni�X���\��sKY꧄���Ŀ��X{G7�o�vzQ㸍�JӮ��86�T�����\3~u��.#4�/���T�{�q���ܯC���)�tZ����	��J���b����e��K�l:�Ϧ��������&��r5f�M��������݌���@p
���sᥕN`B\��iV���a'�.w�$���@2A�޷��A,������D~=L�h�߸<���D,���ⴷ���!�:jl%�x� �n#^B3�mڠ��cM�^��Ҁ��7���qO�t�$a������8�xꢂi���0�`:���'>/1o�y\�j5�}�3�	.�g[z��p����?�+���Xh�������R�IYX��c�v�"Y0N�۫Z��p�M�|3���y�_�E(k�]�����=6U����12�%��!اZ����̣ʲp��SNe��5��0m
�̿���RQv��i�����t��8Ee����/}�5��Wl�ؾ��0�r���y�n8�h���I*�l6� ��~��1����g�����hVN����2��������Y���@��s��4kCp{:�/b���g�́���:���f��9Ȭl��,�Ze;�/H<U��r3��hr�$dY��|�g�rj���&J���L��:���c��F��r��B��l|�V/�6<I��)mM�� (�C7��#u��LY$��EZ�.NQC?gڦ#>���29��A����^�_J��<�u�h@r�]��h�s����� ��&B�;��ia@l�K�hh�+/}�_\���K"'8�o��z��W��Km��&��g�q�O;:�	�F;����x)z�GPF�=T1j�����0�p�NH�����
$�ڪ�8�-��M&hWxn
VbqγK���:�6x��7�����,9@t-�Z�tT�rn���I2wT��\�� ?�ͭ9�O&�$1%���[ӑ��瓵fŉ���
�2��WD\0E����ݍ�T��Rx��ԑ<:/�$o�A=�xx	�B��iJ[�x}e��e*W,a\��s���)��M#;3���e��� �j7Ҙ�zν���ݨ�&uۀ�����ϴ_��2��n��ő�U�5�%��6�Ml:id��e-0�l '�����k"�MJ�ȕvev��Õ������)�@�dH��$A
��*�LЬ�_k9z3V����;�^�KQ	1{	��hP��Ѕ�X�#wV���hƜXm]t5�3u�v��7���%Ka6��]F
C��xq��
�/�rl8"p]�Bs��!���@N�����5�*�����K�1���)��-̂u���s)�܅�h��;�TNO	i�һ��`D���Er�~V������_�W"��.��k��b6����ǉw=-td9��!��*�VD��')�� 748�{k_B�[�O�z��U��p�
�V� �ˮ?�2���L�
�o�ă��<�bx2s>>��5t�V ��3�#�Y��VL��������6�M�F���&��ʘou&�U���L2�W�<~5��k'�v�@Bi5��\��5#:f5���]i�!���`R}be�͖zk�%�";{�LJ�}����P|�A�3z����b|O�����Yu 6���l�.�ʒI��K)$�4���')-�qI`�K/�����GO�'�Ց�3_
8�f��Q��W�}F~��H��@4 �4(m��dJ���*!W�9���6Q�wG8W���5`=5`a�<�����;۫�OV�����^F��HT���ą��Z�7�c��� �|>W���y�&�'?��@i-z7e���� twG�+:�G[� ��_�L
�.��u�����iKN��	�#�g�F��r��z�ΰ2"sh�S��-�|_�T�����:2M[�s(cn�[��V���*�-/o�Zq2���i:Z7A"Ҋx9~ ���A�F��j�����DC�N;s�����q�L���Z�杲A��	�PS]�k���:ف[�I����D�@�S�4i�����$"��/�~��Ca�)A�Hd���׍�W�)�� |�G,�nK\�r>�9���n�g#��;h!s]���*ħ<)��Fd)z�\Fr��Z�$ ��S��z�>]�?v��?�n�z�YP�m4�D�I��e^��W�kwJ���?����D�q�*%}jT%b�Q�d���w�N0W�ekXѡ�b�F ȹ2u�or�ڪ �*K����@�����;� �(#�(�yzm� $��WFB�9���}�GP��� ��K.��q��^�U�W�U����>�
��寵�ꬋ�./�S�@�Jú�Z_�2��@R��l�ռR�F���3O�~�fATۈ,�o;���D>��
���+#�do��Z��Jۖ��N�I���H�21�%�<������Ofn	�"�cT��]ˊ��m��8�e������Jc]����@��<h
��rBUNI�o;�H�.�f��J�e�����d�;�65k&��rdʙ��A4������^�ǵ3(�,oK�*��i�a5n�	��2�"��K�~��%��ލL�YӻE�j��A>�T�F��CiW�w�%B�'�-�{�t�.�М���U�|�q��h˥�xK~d !nM�.BQ�s��0�,���1Us[U�w��6�7��'�����H]xY���x���m]T�o�<�E��+�m�j����G�~�����
3�+@��,�9��L��:!rj��7�ʥ�B_��^Y���g�پ��Y@9lu��}.��d�|����oe�a�r�����P�&m���;�UI4Q��pa�9�.}JY�BF��N�9)e:_�v1�jz��,�Wr�0�;M���sA���p��ݷ� ��hr�5)�M�!$��0.]ݖ�v�i
�	�n�T��Oc�E���|z��rOL��`$�0�Ogf��KND�r���q�+C��z�/I���աAjƣ�|A�� �<��ӊZ�FRL� ��]z}K�T&O{���]���0\ӓF��� ۡ�NCL���wl��W��w��1���a@{ː=�t��Ea"�����rԮ��D��A���#�)^��cY�&�H?�!��4G��W�Q�G���\1P���U�iA�b��չ�����./�F�<�Omg}ˤr�D��cX��Q�
T�ڄ/Sz���Y��w����Ɗ1S�P�Wz��3/�Y�V��A)Vr���<�ބ`��No��+�ѽ鰉�QK5I
U��O��pÊ&c3��}��Lc��W�B���uKD擪�-y't~�0�e��o�lZIsy>8�w���5Q\�;�ۄ�D�Q3+��
���
��T�[g �JF� g���rN��ڰ/mI��ͫ٧ۧ�j�� s���2�QS�e;m�+��m��a��=*���4U����&�.�	O�U	�p'A>~���2<;;�ӥ�nk���������Z�)زJ�>C�f�g�۷^�9Я����<%��r��]i_�u$ �^�\�:͵S�^�W�
�_I��Ú'�g��*%Gf�_je"��S.YC
ڦ�.#ٛ8l_
	���SbUj^���;�m�)�<NmlT���KL�,7����9h�;ԅ�=��m�Dʮ��;����F��k@���4d�j1�O|9\�r������zB��'�*s�(�f������W��
Ɏ��M�jN�^갾�c��7>-�`ԛI*�YEau���/
cs�42��0���Sw��G��Ϧ��ɩK�
,qȘp"A�����'.iX���%;F�d�\=:'&A�!�+-{�R��$e㲄@3�^鬛����u\�#��Ρ$�W��C�޿����ʑ��~�H��x�]/>����}���4���%u�Nr�p>�c�P	t��Ӽ�!A ��]�%=�CdN	��@�	*9���A$(wfm��@�ʆcb����Cꄫ2��p�ߙ��#ڼպe��ئ6d�M\W�>丧c.T�@�*Mj5x1'p�51^t�k�q�>�&��P�q{v�=``�jY�^�~�F}��J?�S̺J�b�a�v++Sc	ڹ���K}��*�4a.Q����{�i����W\ٻSt�DO�]Y��T�g�N���e��8�fI�����Q5Ub|���"@��;��8��}�f�J��
�y qE_M�g���W!h��������v_��ٿ�w@�c�3o9����57�F�\D:e5�w	��`&T�e`s���>�4+���V���ݧ���Į��G=N����;_��*DRq�w�����>%O��>I�)�J��
�Tr��w��ב,�=�/R��N�$(GDn��Hx�T��~Ǎ� �W�׭�%n���
����ܹ`s!ٽ��`��^7.ӝ�>]1�b��U���E1-�S<�z�jۯL� �h-WY�7,���\sXm���iB(f`_��G�'@"�ύ V�a��
iq�eNX�JXZ҇g-�@3�]Ih�#Ib��m"��K+J#��e�uBU �g��Z����C�=�sȌ8��Yh�2�m��Oj!���M�$�l�J�H�ZVS�|��H�������乸�����S+����׵��Q����b��E�
9{��(I[{D
�݂G�[v�07�5��'�F?��nf<�b�`����f�[�V _ϡ=�wڼ��3��<��z^@�[�I��bK�����Fj�P	u�-=4y#�*y'�D,-�,v&<<��g�n�APt9U��ݒOVJ�#� ��m���+
�{鶙�?�E������U�	��R�*�$��L�q��6�6���W�g���m��������b�ݔKO��+�#���oO1�"�x%w��N?i�tI�ғ�m������	6��r���yZh�P���%��-�(�Y"�1ڒ��*�>���@#�M�X�-�.C!�`��&�1�t��\�zӔC����8P��?�����.\���)T͕m/:$�2Ͳ� eǌF;��%����zr� d�Dq����qQ��"p(u�b30H9��K�kaN������~�-�f,ى��
o�`���Wm�s^�u�ˈ$?�Ww��F��n�$|�46�}����I��L�B��ڥ�}���E6�qqϲQvk2N"3��4�&���>,��l����e@� CT�3�r�'7X�y�+B?_���^��eA��Z���ܕ��n��N�i/��S��=O]1<�Ew�O�|��(�&�K���UtXC:��eO���+���F8�B.Yևp�&PMӴR���c=���}T�����1����� i����D�z=̄~L5�������[�Tu{���Wɖ!��w�����:�8��U�f�yMc���Elk�e�^��`N� ����-�Ѥ�o���S�91ES��!'�!k4bxs��E� z�z@!H����M���8�tv��� �����V~�\��1��-	�pe�[/��rs����J��@�w��W�1��b�)�����l�2�Z;W�~X��{O��,��c'��";�U���S/����[��3���|�0�
8.+C�6�/��@Έ�d����Z�f�uP�9:Յ`b� �g�/�j;�Q}�	Q��H�&,�Z�ܲ{=�2�!Yq�`O����}\�q�D1��@~��d�EzZ�)��	hh����`�:���X>n���e�{x����2��pM������b\Ƈ���P�wm���!���cB9�� ���xO�Js�=�7*Fms`&!:��߇3��������D���O3P�8�N�6&��6q[�Yr��M��U����@�͔t���"�����.��n��M�s�)CB"i}�ʠ�}�1�Z�G0�K�3� �֯]�uF��R�v웂��i�P�0���A*�?�>�U9���p
��Ros�{��{�/�*e@MY��$Z]�&�w=����s�k
���:��P�Ys��ݽm���/��P��(���r􉷐�&�Y3���aZ,lQ^�菍!�&O����)�Uj�%��[��ł���H5뒬��z�"�Q�I7T�i�f�&��X˜�Ysk�+c�՗�8�*�����j�������)&���UK��	�2������!z�::C�'��-T눧C
=��'����-%&�[ ��҆/����٪)zǧ��ᬊ~��P/?J��BO��~��T�;�[�y������f�����7�JL�����7�#�M��ֵ�Ŀ�֭���;�ɭ�xu�O(3���?j�('��\LBV����}7F�bg�[dK�����ԉT��h\�<R�cER���!����ܮ|��"��to��x/n>P�Y2�p4��8G?�a��31��!4����`l��� ���u��k�eK��8R���_^�m���h*\�<�JBՄ�*��e��M���@Ყ6��!�:�P��47N��&���,Ԣ� �����x	r��%��"ݷ��^�E�+Gϰ��c�X��)o��*���#9��YLFO3ݾ�'�<�f2�n���Yb��c��=���̽�F�Dwx�j�p�����u�,�s�	Pr�8˟�Y�s��]U�sE���{;�O�rh�d�r_��X�f�˷��W�&�qKw��k%>O�M0��"6���5�e:)� �B/��-_��{�~,׃�sn�>p���\jH�C�<kb�8My�w��N^�q���BtǤ�J���n���c����je\E��r��oa'�Ӿ�=�����$��b�$0�9�YOd��?Óz�k�_��:��Z*3˳ié:��=Ȣ}Zz�i�_���<��E�[�U��5
���IW#��������fݾh-DV�+R�'��t����0%/&�I��ڻ\�e�)���rb���� �m%���⢭�5-0 `��ۧ���܁��u����H�?�1�t���PH�A�'f�xV�1XO҄ȏ�7���k����8:��f���F��R�je���{�N�d����q%�sQ���0��ǅ��u<�D�;�ZEo������3���P�M��TH�Vfr�M��TeM7[I�e�$H�H�-�ͳ��rG������}#§Pl����#k��cRt0����C�W9n���Iꌏ�3	��	�1xX��e��C]�H�9	G�p�O ����6����e6��vNث [+p+�ޝu`�W,��=�]�Hh�v�:���8�-�̕\���$j�/�hڬ�[U��䴫��<KdtS�� �eh�gk�*�x�Rd�,'8��2���P`1�0�f^����+��C?�*��Ulg��({
����S(�&`�x0� �i�lM��@��G/hťS������x��YI3��Mc[^��l��?.�7��UY5�D�����f$k鲗�A�k}@@�vH����f�s��2�
S��9�����Ԑ ڔ�U�֬tL��x�k�o��U��y�e�y��C"5�4yI`���ܔ{jn�\8VJ�.�Q��c�+1��şI9��@�����yi<��O������⡤n$�k�G.	e:���N�PҢ�T�$���`BzV�a�q���YFfP#w�����Vg���� �3F�T<�_P
�~[G��]x(P����0�e�V�}VT��OX�ў�W۩���|��������k�����g������Z�C�\�����~^0��5��{�x4h�gx�t�ҍ�a����mLڑG��DZ0u��cK���yytI��	�/���c��E��/x�y�������aLV���ר�	t*rj<9��CrW.B(�U������i�'�1� _埼K~UQ<�T{�}c��aY�W#+�~��AEs�&4��g�� i�t3>����u��6C���t�;�RV�5���\���e���(��	�Ql�j�n���R�&�f]y��H�J����Q����Zj��qxsv��jôo�������F`^�������)>�˾��딥k�sA�H� ږ%}61F{�%*��C�x=��A��j����8ƃ�F�=���e��@ї	���tk'���7u��6���?�������ei~���M�~�3c�){R�SEL��_�f���ܐT�o2��D�\�����qj3�z��������)�G)�9&���2���\f�X�;�7����F��,�K#8Vsbw�xF�߭{��E�G�O�,s�4nP���cG�C����;S�n��P��𘦤1�����E��#��F�p)��l,T]q���5o�9[���^��H�*�n�W���0u���Ol��FG1��9d��?��X ���ߤ�Ƶ��;��7���{,�FYwLAT�I:no`cgZ��8��M�1/���������Y3�SL�c<gG�Tn-\Y����QƖ�r#��o�YE���4����q�oכQJj����7��^��
�Yg�i*�Z��
<T�Ӣ���z�)�]���E���C���ce��f!��gQ���Ғ"r��y.�˔~8�����f��D�=h��,�`���F19�d������nT�����x��8|0���L��h���V&)M-��6�Ϝ���"�l���t�Eie�	7��'�vi�;��\:�.si��P�{n�t���z�T͝�(U]�8�C̽�"�m�Fnj�;U�Kt�.H��!�h�,�ɠ�i4%���>t�8��y��?��d����_����U�y&[�q�ݣ'���VK�����4�g8E���Z�G���3Ō��Vi�{jPPO	-�M�۸��s�6k�@T����7^�x��(��mVQD�8J�|���(2���>CT���O_c��3���~�[)�	��C �˫��VM$4�G�N�!���x5W�h����}�^���� �(�P���2ʥ�dv��M&�p�;2�����n�}����*4��7]�SA��40;*�l⎏bRO��ܥ�v��f��o"�,G4�]A2����I��Z_��R��C5�<��f��	��9zY�i�;���8B�%�6� vݣx�4����2w0M�..GlԨѐҊs�4��)���@�
�{�Y#�\�J\J���P��(�G�[rk/���H���pK�Ld�y�5Ҩm*=�gEW�Ǖ��)=��/I�,�t���!ߡ��H8V�ko�H4��5�v
A��Im�*���{�;o�ɚ@f�{�z�<�����i����d���}.Zz�#��F04+(R��A_ț_�Ë��o1�8����S;�,Ǐ.k+Qx�b(>�r��ݱ"O% ب�E��?�ѠEY}r��3��%��B��p۴�rWu�y!Q.U��\�+��l0��z�џ�zr>�
��U-��"���P��!I�X۶t���xh�B~M��XE0/��H|��"e
[!O������i \��q;Ѐ��]$�B��*��������#�G�gbI<��{#E*�_&�/�f���lD�LU�д$'��o��q�����f�]#�3�.�<	�tK�.$�cכޠ� �T�\�h�b[kkB�N�_��#���|fG�N�P\�>�F���Ao�YK��Z�"'�Ӑ�ZSp�f7�Y�(�0i���(Va8� >Qbp�%��%�x��yc+����.DEv����U����#Kx�O��~K�f�YvS�J{������"�	A2+�5�s[r]P��,���\󖢟�"��X1.?R�h?o���ַ����_zYoIx�Tӫ�)���"lQ��j�-���y]�=|�y�\D�������)�u�1��,������HQ�Ա�%�o	M����{��)�{"[U��˂�L?���������^�0���F���!(�ڮZ>���U�ͺ�7(�]i0 6y1�vԁ&�j��ע;k9�P]I]*3��`����>¢s|J�>-��aG� �@�����@�1?�t>3 ~�Kv��>w�c�ûY��N���R�,��z��?�a>������rD6m~K?ȾT��	֝#�Ӣҕ�g��&��R`��2�j="5n��z8�X���"�,�UP�sjE�Jف�'�:E�q="�u��T���-�&_^�k+>{�`�_�3[N�P�9Dz	4��3cq_o�!�|S�������-j��8������U��Q���l�tm��{��r��4J�?p�E����K'�޷�/�a߸��c�0��\���)�|* �G~'A��� �DV�g��S�������!2w#��|����z�2�	�(S�V��j�a>���T�ݑ�N�Ĺ�j����b��O���&�1��R�Xm��$&uB��Sx�3�!�����+���RP�p�5����v��n?;�C����^V8tk��[�$���[�\;��ȅt�n���vBޡ��p��'���%���Nтn�DX�u��=����-����C�N�3��.�tT��d��)�ne��rZ��=$�T�"i]�ⳘK��a8�fM@��i�Z�͉3;_m�%��`���#�I\Uj��-�m�)C�|V5bK��_�l��ېlg������F�L�r2&$�+�ҙ�������ZL������!�T�r�%w|����ޙ����\�E]��!H�.�S'&�	�`�P-!�-j�_���x��hff��[585^���e�hst9���k0�{�I;�J��<s��fw������Vj��#V��LD)�����!/����O��� ��.:��#��#�À�UA�t���"E����О�O�Ⱦ��0#S��R�<�3\����B�t&�M���X��+�)"�N�se3hE�ǿ�o�Z"	o[���PUZ�y��l ����ZD%p��﮵�l�P���mvHֶ ��y����Hךּ=��ƽ��z~�
t�S���ݕ�2����ے�"����BU�*'=V�i�"ٲ^%��R^�]~c��{P�Z0lՊ�����"Ǟ��t�0ʏߋ��^��|v�9�9���"̞��� 0edty6�V�/�}�ɏ�֋�W�001��f��?��f�<z��16J�OU�4�̣_�������iI�5����z�"�ŧ-�,��y�ʗ��SM��ރ���*L����$���^�MBhE�w'����p�-dw|v�7@��o������S*����>!�Y����4�����<�����0������-����� D�q�R5���D��F��I�hE���VQ�b��).ǘ�~Pq�|��z�ՌO�˅[�)�W.���zR��j̫�{�m��}r�G���e@��L�4"�I�|�I�����H�ݓ6F�vTIjMhFҰ��
�G��W?���AUք�_(9!!R��A�ˏ[�4��P42��XZ�
�@[����~w5���u�yW��\�D{���؆��8ڷjaY�sv!��E��Q���O�iI3`�kl�'�
������k��L7+0�en)���\���F?��Rqӿ��iQ�m�g��<�($��2cnp��)�D3�Ɩ[Fɍ�h�&�h�>>j��>ps݇x���ǅ �lsY�Y�bYH�C s�	l�v�Bc�i*��rmn��Y��|�Ȅ;t=qm��O�W�䝰��{o��zD�r'NH�T�
b `��%3Y�����Y��!�g�UHΰ>�)�_]�Gi�,�u� Ϻ��a�x�v��n������b��3�i��� ��`�v���PkƓ��։��p���Z>����)����A7��e��G��^aؽ|t�'�@��b<�X	�9�ĐL��I?]5�|��?��}�(n���Aa�os�f�R�9	8��z��&f���ZQWЊ�{�15k7)H��]&���Y)Ÿ��u���>�[�������7�i2���L��͊N=6�)����>ue7��*��R����i8D��y�|˽ض�RI�,�bO/A)y��7�y�V~���U�P�q��?��'�15mb�P��=����ڲ�C��pBA�F��^�gh`[�så/��J�ԃ�^�dr! �� �8��pW�ۉF� t^�Ey=�b��k�P�Z�iRC��-�ȡ�m�:�fB� ���5#�(v1Xe緰� ���(�w}��Y�