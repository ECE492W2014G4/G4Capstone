��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P��v�"<ߞ��&'��k%P碶�R�ӣ�sĞ������FY&v�h��aJ���q�[��6��58�}������u� �-Ǐ��L��ݡ��w��V
�q�tf���2͠�ϫRTŨ�x���L�@�w%����W�& ���1�Ѿ��C�Xh����`8�8Kޓ���O��$$Є��^���<�4�4z��vZ����w��b�cLi�Ο�G�C�6j�**�uÜdѷ�LV�Fd��Zɠ㋤9����+�62bmW*1:g!�n����x�g*�jb��'��6a(�I�m�N�>�
Y���J��bނ��ykc>S��UYHZ)�&>$(%�;ٕ����N�|I+f�|����+Bw����+B����4!TvΡT�+~�':��|:P-n494��w+R��$����� �&����9,;e���l�1��t{=��*݃�p�!�Y��Pjtm��8W���u+)@�
�03��E�Ԟ pL����w/I����fRl�!�s�� ��)�
�^|Ï$��bu�;zOǍ��N�+�5n$�.7}��p��Q"���O�(��A|^ĉ�����c��T�^����;��
k�ߗ�r���I�m�z2������t����|\�B_�M����ڦD`ROZ��}뢾Z2��6���l�4�M��vm��?F�?��hH���-ؾ������R���$�~WD|#��o�\eUEo�Քq:$]�/T���
D6Rhh˭�����V!R8���������t2ӞN�>x���;���l&�B�˳�9>�K}}-��!������maQaW�␯U�nsF֢T���R���z����1?�����<�*���Gv�3L�������W�Y��13o!p�1&(�\�[�	ب��v���%�M�Zm	g��A�:Q�_�<�s���3M��?QLgt�$H�𒳨[�ɼ|m=���(	���
��w]��SF�r���0�a������U���K̋ w\(�uJ}�Y&�NY�}�}���
�_Q[։M��w�(ʣi�~�x�u�J3�}=���v�"<ʘ���Yuѻ�E+'�$�p.Dl��#$�d�7���]�F�l.�M+��ty1 �ċ�Ѷc�L=�;�!�8���%x��$��� �\?�������T;�+����.S�HLZ��3D&��~q]�Y<gx`�#Q�q;������z-07#������H�"��S�HW��"�ܵ~C�&-���p��]R���/=�Fj�iU����=��Eκ��4��?`,�5}vgXC�XYT��bE�x�^ѧ��|[��`�}J����>�T����A5����!�Ár��{S1���͖B��)�sVN;Fk�w�_
�{׿� 4.�%�h8s�P��C���I��}��U\�Jt!D���Qp^�D���V�3PN%ĖI����,N�j���鲴�v�c�Q1d��pp&]A�V+�i�������*U+�Q�G���x��y"�^>����/:0*�CQ
Δ��}<�B �C��͛	C��
Pc�D��GL�KW�懓�s~t�Z܄�EP=���06�p֛E���	��5.)m`���ǋ��r7����X����3�Z�!
K��V�`���0yFga���h���Sm��F��<�tĶ%'ޣڥ������R�U�䊘z���i��:Mhz�p�߲1�na�ŀ<D�������}��R���}m*�z�����Rk��3���m�?�-���tk{��?�Iu�|J�8I�ޚR0:��R+��kx �ܵ���˸I/�;Ɗr�S��PӬ�m�$Bx(���#�n`�k�������z��Ey(0u��'P����V$!�pk����V+ZLs�?1��W����ɿ`��B�`��P]Ȍt^*��Phx��J�=�'\[ƴ:k���$�n,y�(�_�<���; �u���?��hN�r m�!���HQ���]
�����Si�s�1m���1�sɃ�F�f�W��EB���=W�>�g���4�Q�W�n,Tk$?��"�73�d�Ҕ��͍�Y9M�Z�qGlC������C	q��:7��7B���4�s'��Iid��pCCL�k�%+������]����=�q�z�~��	#j���!�c6ϙ�2f=�pB�zް����#& Gɿ7��ZPo�c�&#�i4I��1���4wK��S.�Pe����+oG�L�
���V��k~��+�L�ح籧�YM�4�l<x�x��BI�������.��)X�(r�+,9�391����ƞ�=OȢ��䗒J��Q��gɝ.M}�tw��ޕ.q�Ƽ��[�UV���j��'Q?w��a���VlaHO��v���kދ��~�$���!ۦ 4&:����n�.�t���L���v�U5*��$(ӶR�+,�V��ns�\��������[93BD\�(FwV�ǧ��)���]콸Q�Rd���0OI^ba�_hP��^.I�g�&s?aM�J� R!�� $�B�( ���c���K(�Hp��HBCA�QݓY�y�+�����~u�3+d��~�}[����8R��ςEv"�\F�q(P�h��{�J?����~��i�{X�X����>V���L����|P[�h �&���8�U�W>��b�.p��vE8C�0��@��69t�1�􎿢{�󱌥?�hQ�>� 8�C�����'�m���Sݭ���Q'R�m�[֭nA9uOSͮ5&�w\�uS�dgwhs,lMt��d��{�H��<,��Z�������W��R����>�<^*��?UB�;���Jb�b@Ș�������H�ӑ�!Bp�������I)%�n%��p7$ ��ygEeEt��M���vr�[3��3�L%*��a϶s��r�9Y�k�3�����/�n'�|98�E9���?qq[j0�]�p���FӒ^z|=y�
���w��r)�"���}���
��	u�O[[����*���Z�O$��Ց�5ƶ��>7Ϫ�U��<��:�?�)�VѢ	X���Lo>�P8�[_Ì�gL\0�q¬�!,#���woi_`�^�
ʕ�xd;)�g��R���62S�Xr�v��܁�=��S��x|̥U3±�ؘ�}���z}7����٭�~�/8����%�\v���P��S��6�T����3�$,�CD0ʍ��&��C�� L<+1 Ծ�Goa�ޑZ�1�8'�̔�
���Ժ�C�W��~I��*���:IɎ��s);�	Z�1S|שM�NJ�Xaxo��z���ke쫘r� &k-��6Rz_x�F��=e�"y�Y8����
o�9߭ټ�^G,�n6�������Ѥ�)Z�I'�P�;�|��cu4~a�CBp�.x~�j�U&n_,�鮙G�,D��@���怒��g�LYǟ0���&'㿩��tXd��/u�fŭ�����18M�+!4��ҕ�L9�b���ڠ����*^>���%�o���s�3�4�r�I��io�4h�?3�d�%�Y��%-�@0���,�bhT"'���뭴��(�y=�,r�b�TLk"�/�4������<��\�
}��lU�=k��N�*����1�H]�Y��BH�[b(H-�̦h7��>A�P"��x��.�����|������3�u�sC�H�UŁtڱ�2´� 0�r��]v�}��(�������v�"�O�g:ƩmD�_ƒT"3h���O�~��	���4@7;�Ԩr�|��rfh��[<���=�׎Z�I��� �.4�9�<��r���Y:0dr�xpY��ڐZt�#2_/ǒxKT9�􅘱&�n9^+�נϭ�9��]	]���.��@����׺w���0�q�+ūʪ�A%��5S��&�GL*��nFV:�0�/�ج��%H�4��re�i�zXRFg�<��n�N�'��|��+&��?s��& \��8�Dݽt0=:l��{+T�Ίr+��Vd��l`��lMu�~��8�zM�	��`�Xr!���#�����CS��ӗU��^  4-U"�O���&�"1�w�(@�K�4��~3IhlL��q���W@�?�����c������Q����ez�c<a�ZJD��-l\@32���}�jJ�X�p`�ݘ7	o�s�L��ջ�2�~n<�%��U�N��\Jf����?�c=���8����RD�vG�ඪ��Z���v��%A�DJ��+�%C���Ə�M���n�y&�<*��ժ@ws ���jM��U���'v$���|����a��#��fYC��%��xQ�
���}�k#�OW��5�H�X�c�)��ǥKhq��K!A��ke['�|���j�����[8�+�ol� ��-S����k���>���`��-�;�(�
����l��l��"��%?i H=�o��*�^�d�B���>!"|��TQ��R\~̽�{��!pNP��X�;�ҍ�1&hZju� ��w��~��J+�fhI0Wmt��1G�Q
J5�.-���7��f����id�vG)RA�ɫ�$���f�u|ܥ�����i��MPN��]zQs�I���k�F�-J���-�Mn��Ųr$�$����A���7�%�e��ࡌ�7����k}�RV���0�F�D��n�/��'"G+��{��V��2A����7��T�x6Yũ��-��"`�A�Һ���6�=H�;c����yض$h[jØ�[�c��2���$a/]W�Hh��(f�E->3P��p�bߓ�T�80"�=��Bcg@8��Ú���3�a΃��t��6I��v�6��Z��N>��}�6��}ן��^�Agf��*�}v��8��#X9�>�G��b��5�h�9�I2���ȓ[��U��y:�����.[z��>a� �r%� �56q�O�bsu +�k���Sf��%�^��-Eq��^qR��R)r>F�THc��������"�r@��*Tɘo��w7�{��������wx���j������὜��&>-�ϸ>�c�H�3x;��u��,�;�n��&��U��1a�����m+U�6�i�2߶<�?vgX>��U"��'ZO���t���UMQ@�	.��;"��7 iL� ���+pWe��m�eq|`/�Y�r�MF|6VHg�;y��yX�L����)lS�7�'��Z/��� �[������RH�ߋ�_�~AvB+�r+Q#����Fh�M��O'���T�Nr�����WY]�aQ�������#L�BB��ŽFb�'|�.0+��e�� >�|\�}�L���g%��gX��F�w<�>�_>���0`����}ג:Mv�X5, ����~o�n�D]���rf *Qe�F���A�tϾU���s���W#�p�z�
�)M�9)a]ߴ��o���,�.O9k�J���F�!����>�)T���V�f�s��t��q�!
	9�o,c�ĥ����܃-��8%N��Db$�Լy�c�1���7a�#������s��s���k2�1�;{�A_�ćSLte�K�9x������[i�ż?5�ա��@�i��� �h��e�0[���J����W�YN��W�}�l5��0~i�r7�c�B�CgLUK�f�t�q.ʅl�kY�.�?A������!A�$�'T%O+`�m+%����si.g�� ��GH�x��9���¡ҙ�4;h�e�1�t�b;�e/W�+Ոʟ���h�7w�/���ۏf���1����-��R���[��Ɉ2x1-P�c��_�ziei��Pg%�i��굷���L��0d�ڝ0���J���m�ѡ��9���#�w�f�f�Z�M��7��~��=�g}k��8�}����)�Ŧ���Jr�tĆ\2=�����n�m���if�F�z��4�ޠ1�Q�9d��ꟿ���nP	�.}���άN=$Ǻ�SG��nE���=�R�3�K 1�&VD߭��BB�*;�=&���(hI1�]ﲮ�b<*�!�4��z����6/�Br�X �o����N�\��ڤ�wI0��e�SmmPen�*��	���X�鹐��Hզ��U�e<ڱR����K
��X`z"�32sE=9���	]�p�<A����N����9�"~=B\��Ph�u�+��P�6�9²�T^���v�z�n�G�M{�y6����1�زw&���G��(��]�$���%��٘��\�������k�l��2QH)�lo��Y��&&���oq�㇤��<�Fh���a~��p�x]
�x��['�!�U������z���_^Zp�D�Ub�W���[�H��1�#z����Ro�I嵞���ב�"��L]K��c�rrR3��#UQD�t��ɇ���'92)j/�l�9��7`�Jg:މ�k�<7䒷H��NWs�f_B��)rj�X� �g#���Q�������>Ñ���D_�(!^�0� �p�1BO���Q��;�3�`%čM�ˊd^��������9�P�6�p�!�jy�1�a�,�c�@r��1 >�zX8� �7��<}�V��$<��E,����ʸ���EUTϓhM�rnA#���5^�$��b`P1�|���߆�4j���cG�rA�y+:�m����U���C���1�Zq K��89��P޲ �}�`C2(Od/9/JZu�3��r�����`�?hI��$|� !��)-1�DE�/�cxI3������處�s(�c(�ݷ*�O�����0���rY�;��̂���,V"�L�:�1�x���e����(Ad��@_o�ԡ�ɇ��>aO!<�G�MwP%�� ��2�/E��/�޼�XR�q��˺��A����>y�M/��w^ufB`�Y���_pU��NN8��И��ܭ���i�~$ۜI)�%�v���`�����{�����@)ֆ�i5��f��;D����H��__�xۑ`0���C�Eud ����M/���Ӷ�������(ձ�9�u`ܕ�9�Y'@.�7�B���!LǑ9��j���K�KS��]GB���"F��<P���E�_���A����@U%��&8���%�R�*!K�7���
N��*��# ��E��F�c�VVӛ��(L�y[F�w<� �F���n3U)��j��P[�~�T�.����0��9�Cr�gUV��+��q/�Ba~������=��j�[?�TC����(<�&���E�@���l��� �q뼾M�bٌ��.�e��,+�ৌu�֠�ڛ�'�[��'�\����������z�	V���bB���G�����4�� n�N�����ʈ �W7�P�B�0��C��U��Jv� �~K��1w{U#�6
���9j��:�Ar�߮ږT����w�L"�x	�2� 	��)-��)�\8�H��ƾN3�B�Y
ǠP�U���A:<sqv���LV6��h�(0h{�'?JJ�P��z���$V�I�\[��Q4� =T��"�X��?������ۜ�F��G�Y�޳�;wA���dF�P���po�Z�Q����8ge�F�P#���Z��T_:�`�KB"�O��D�s��Y��bt�r ���?�2�UiN-!�ؽ�J�	-�K�K�Y�]��&��yy�3��5�̭y�sV@t�w@2M�f���S���	�����,3�SwAA�J���:�}J��
��"`b�e!�Jt{�ï+�ז-a�|�l�	�����޴j���.�Z	1� 4��������M��)�9���0}%Z?�q=C���L��z"O�vr�	��l�Zl���#��ݵ��4�?!Ƣ����͊0F��a��=����8��5���+���1bψ���k�!Em�MB�T��7y�곲*�����h��w�8W$r)���B���'�	� -E�K�*O	��]@�K:Z}�ٙ9�i�ؘ`����,>!u,��E�K�%���Hyc(��T�ت��-��/�YB��ym�˂��K�WL���A�"r��^�s�q�iP</���;x�~"�R�|��5f̷u+��0�$$.z��u���� �vn�2i+}�]"� ���ʸ��[�#��|/��
ߘz؃�O~�Ѕ/(οJ矢�������]��]^�l$0V3�V����
�R�U|$l�i^g�M���V�җkUg��=�Q��;o��ɔQ��l�����3��	�	ў��0��Ĝp�+k�_޵\ȇ�.��N��T�>��y7�lzD���9�mTt@j��z�`��*ʗ��.���{b�G��
�K<��U�7\c�% 	�y�\�"����i?3n� FM��h��;�h��sRa$:>4��_�E�/eV�k�u��BC��G�K�>e� �P���+��e���\���k+���`
z���v=U�����mћ��=h�դ�s��W��P���m�V~2��"G��NE�jMRk)�C�싃��}��DU�==����n8�j(��d�7l�q�Dmn��aP�C��C�>l� �3����$\a�Ϣ�>��3L\8��$�"�r��4��~����C�S�KH��E��h��������B�D������`uZi �woՙ�Ũ��}���ރ-WW��jjo*�e^�'g��uo �z������u�h�J�7�Ro�|Jި�j5rÅ��t�z�>1;=?s�A���DN��X~��W'e��s�)���:�u�ٔ��_ :87�v��ع����ɟ�ΐR�+n,Ȉ�Hq>������iM�ϗ=�P���M��[Ea�%�Mz��j�'2&���M��ܴ�X��t�MB�q �B�]���o�x�;ΨW��L�u�^N��5�m$A�⁘M��
g�"��әD��Q2�
���[,��N���|Q\�,v	T�k�,��|�}����!��%'vN0�$���~�Clvj>���|.��x�"S�����+��Nm2�X�{b��1��?�#0