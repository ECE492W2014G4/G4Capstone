��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P��v�"<ߞ��&'��k%P碶�R�ӣ�sĞ������FY&�E������z��*.7G������ .��] *�ʧÀ��FF��j9�kH��<������rl�
�h�5���2er8��97#G|�	p���Q6�4�v���&�'u@�Ix����m�?+aS���"��~qXCɶ��}��F>�=i��d�B9����J���B(1f /K��qr�z��n�\D�Z^�cm�E��j@�@���߇
�t_� 댵�6з�r���7�7u(�g�Y���|��#K"'V
؆��������)?Gv$�_w�^T�?�]��q�I��̨-	@����:�o��7foD0��'[�hj��^؞�����qg�{{"��?Lv�B&[gݸGQ��DP�����DY0	_K��ME])ѓl�ɋ��M�6ejM��ji�j�S�u�@�?�v�<��Ht����Qwh6�
v���ը�yV����߾^-&��/�t�x�
���U��h��ser���p@pl�����,Vceq'.8�.����Q�w��6jA�F�FkY��_"CL�o���ɲ_"x�s��Q���ɭ��s�`O%�G<y��鋝���>º�%Ia6�uh3������ �! ;��8|PL!s/����jj�,X3֓��-�#�U&L&l'��\J�Xș���Fc��[����A�k|-k��t�k�8-�xG�W�z�ĘaT!���&~`�Sp���ʌ&���q_vĩ8��R��?,�����ِ��'�/�ŗ�o�����R�<i���JؤS�A���t���s�I����C��ǩ���m��<�#	�1A�<;3kV���N%Z @^i|V�Adh��V?��
s��2(͗ڗ�d����u�m��e��~'8�t���uk���gx
en�~Q}��� ���5�:�o�qq�R+���a�c�=���0��أ��80N�i��~ ��.�Ԫ��e[�^�,ʓi�~���g$lB`
�r
6��uQ�LڏY+�1tm��['=���I��4�N��;]�-���WӔsΒ{�.�em�o��l�vV{J�[]J�K`bN�$�����]��	�)��󉾬E5/����&oB 'YM�����t�\��[�}��0%�[�yvQ��"g(W�At&��٩�o�S��r�d$K�Shu �U������k�i�z��<��h]�^u5D�Z���Ec�G+J5���+/Ga��3/+i�O-��G5E'$��sF�QI`�{ttDHXv��Uv�P6@���Z+7��k�۞Q���~��$�G_?N��o55��`9fg8�DJ��e�������������Ia�%gڋjg�wђW�W�io*q�K$�f����A�]���^�TsW�4W��F����,�㊎��>��RsV)*oXQ�{?�ʕ���Byt����w��@��!gde.[m�aA��v�=�i��{7���U��$sU�i�v� �#�iAU6�v�f��?k�0�J�Jb<by���DF���C��A�[+��,Z<�[2���#Cσ���i�z�5 ��k��U��y���,�i9�l��4x��!�rsᨲ�r3J͟��ܮv����ڌ��PLZ�`���+��>U���>ٔ�oכ:���v�UO���@���R�o3��L��kz��J/6U
�h�"�GQ�5�
:GT��p�%u����X}`�.�C�Z�TN*�R7�c7H� S'_��䅱
�q�����d�U�ퟻ���^x��6���o|pKy�(���r�����:�/4�{+��?Se_��m7��ֲ����z�!-���,ZF���i��$(�|�u�4���(����� ��7�aI�Ɂ��U��l����ܳ�y��>Ǜ �����gch�\�y/&�)��-�����߱�f�	�j�F��CD���W<�z��Y��8,4>�U�H��������m�����ɼr�a%<i�eLa�K�f��mg�zjuSƇ���z�`���Mab���1L�*�JU?���M��i��R�h�*������4�J�7���eE�X��87�e�ޠ���F��Jv.�*vM�
9\�i3[�o"��?nv���"+�	�=u��>���$�D/����'�6��e�8K�8{L��
c��|���_�+�H�<0�Q�A�|�Xl�#]ì�g�tG����-�]e�F����1���
��n��UL���u�{ �\�O�p}	�H�D�)2gᤰ�W�x�������~ز�V�ђ� �w��g��p9�]�����u�0��|����:�o!�7,�/��A��ǡ����5��m��ۇ��WW�2�����Lz�s��,���53�@	��]�P��O�3�9O1�
��@L��M)44�}��L&dW�Rl��j���l�����{��-h� j�Ӈ`�!�M���6��ԛs(��#_���B����
�d���� y-���C�u�r�)_d4�,��Ed\=�bM�n���8�k?���\\������v�)z,�����Y?��=�N�6�@�� *��/�,~_zE�Y�'����4k��]��HDf�7�qga��&�U@�2Y˰Rz����!�\_h�ǃ�	�6&�Ⱥ_~��a�1x�Rjs�w��l*���ꎹ�ݰO�Q<37qZ�f����Y�X��ju0�+S��$s��/������W���)�à���e�R�M�ɯK�0�<� ����^)�\�l��=�W�}��e��w���pc���+���.��b�%դL�z���{nP��D�����5��	H =z�bµ\�sy�T�ӵ0���B�H.�`0��Mpc�n��R�Ii��\�鑴O���H]���*H�媺�M�8L�?[)<Y{��v�-���֓ݏ@�[�=�߯p�y��@�1$�'u���l��ryvm�x]�,��aO8cZ���u��w2-"��y����@�~��J�Mc��έ��\2��E�����K`��[ [��2"aj���+7��f�D�h>7��Z�iG�~L�2���)[�� �HqVg�~��Zz*re�,!�ta�:|VƼ�$A*{	d6f߭'��62E�������g��\B��^���;�.��#�;�!�_��-S��z�uf��%�;Ӵ��v+a8�=$KPH�5Y�>���ͥ,q.�p7��m�и�*L�{��"cI��ɽ�Ġ�5�eم2�5Ln�-��S����:c�m�>��r/�\��6:�ʄV����g���|l����ˉ�9N,Xy�1�'�H��ʋ��T�JQվ��٧�v���[�u����0e[��n�3t!^��)V�[I��Ј�5ɣ��&�P:mò��'�����i�}����'\�[���=��o_�� �&�`4G|@T��E��җ؛8�ʮuq��hu�����JmH�v��!�N��-PX��1�p��w��s|�@����+�����C��G���D��j�amE��O�h+��������	�� �B�X��Ce��kJX;��i8ڌ��G��	(�-Pie���H�CY�A9q�#�A��A��]���^t���L���<��U��W�@�e�&?}Ջ|��  \��0�8T��j��ri�Ŏ0�Pe������?ڹIt���Z��-^{%h+|���F�`�Oj�@��[$v#���(��������&`C���+����3+Hc<����DwZ
f�l�L�;�j(\x0`b���d�jD����{y�%��0g#8ƌ���#���u�Lۛ��a�|�^��V2���U��������߉��eU�>t��iN��Tm�����Y����'A�h�ԭ�W��}�V\y*�|�4�a&��^x�Cf���ZD��փ��[��6O�÷�nH�� ��-E֯q3̯LXE��S��;9X{	�~����\2��t怯w�M�����<����C`�ۆ`���V�S�C��[��3 h��%�6:������O.��b�Ǵg������3c\���gf����G��LU�2.+����\&5��7����b���5��p���-`	ˤbb�A��{6_t�V�y�UY�D�<�K,TϷ߁�W~(�����;b�ӯ���^�����ء�E��As³j8�d����������cxȑ��T\d��¤Q�J�J��Cۃ��+�*��la�Y�@q�[��l�Ҹo�|���`��k��tQl��PJe��l"Z���4�ߧ�E|�����[��(�+�^V�P���p���Ǯ����Ӫ�О��:O�C����Y$� ��Y�nJD�r�+ٓ@R����S�O�yT�h�֚Q�O	VT	S=���a�}As4dV���GG:-���q��6��[f�&�&�
��#%�g�ޡ�����U�
r(�����v>^؁��8���brn"r�̫!U1N(�������#��0�.�Ln ��yHRh:`�bcG��ˁ���� RS����C�~nwi@2N��^+��,�4ɲWظ]����d/3~��hH�_���*��(�&v8��i�u�S�i�-M�eZ��+�"�DR�=���f��3�)��?�'��J��I�m�!����	�ۂr�wܨX��eoa+J�T�,ҕ�8T���v�F��R��U�X`κ6�a�v}Oɽ�'e��f�<yA:~�D�`������s�Xn�@=Y�^1=w������!�U�^j��=6LVg7��c� v?�z�e��7���J��V�����Ьteޗ��3���XX(��|w��Z&�>ǈ��q��Ͳ�$�p?�D�}Mt�>�+�+I�u�ܜ�s�Ҁ�b#4�۲׮�v��Jr�)^5&R�na�7�����¹�t4�'�AN#����Ŏ���)7�����B8�ϫ�x�^��.!��Θg��)�B,��l��/�����4��r���g�v#��Ké��%��0Q
Ñ�����I�#�����0�����-$�� ��x1��xQ<]�Mc8���N���I����K,ĕQ��=�O����4�7���ެ���lܮ�;ˀ�՞#g8�e�zRP

�wd�g�:�&+ب7�3�E�  h�C�Jo��C����h7K�5=�C�h��6���n���١�n6���Yo^�@���0	iH�Q٤�99�݆�����VҲ�=⚷���=��;��C��q!���s ���lmR	��Y�~o[��[Q�Q�Q����٬
ү�U+	�`�a�+�l���oK�U���F���b��؊M]��ԥ�a�^�n�	����Q��/��Z������!3}�L�*$��T	L?���1�	��W����}���1ߞ�U�P}�G �Н`G�}ڒ�H�P��"Y,��=�\ȇ.=7�㫺k���@!��5ļ��9禟�;��4�e�{�M��F)!���$���,8{a���J=��#�����y��t�b|#%#}��`��X>.�z�)�&V�5�&�9~���v��C\R�o<�K�*_e�K2֜����K��.�����-}Vf��caGy���DU����G�G����� �NkS�"B=8���j�@yZ;#&<8aO�41����(�S����	�\�[���ߺ㦤a��Q�6�-�y��Iġ�V�z��yR��l\�ev�.��a?����%T��9���OmKO�@ b:�z�ː�7�����?�_0�f������X
�q�1ߧr(��H�s� ڔ�⟸-S|v�n�-J`"7�r�����kܥL�v�D	cGX�٨_6V�H.�;���%���BB����]QT���7C��k��a$����Sb�S�'�h��3�]?pS�C�W��(�/�y����������ض($nJޢ�p��Nǣ��S>��<}���o���cx����=�#���Ьq6̭A����n���/�`)�u���<<cA"4џ\�B
)u�<�R�(�k#fO�$1���n��5�"��	v��φB�7����k���w�6K7ľ�Jt�2��I�Q�a�iĒ7�v��ۈ2�����QiC�U�S�
����q��	f��/�a���=},�SŐ{�O�6��2ۦMy��N��XP"� [���HA:����{Q4�f?��� _b
P����+nn�z���:_4\������դF��j;�)��wRB�ʰ�����w�b%&�w$��H�b��%���]��~���)�����(F@-!��|��3w�%��'c�Pd��JG������q^"�����Ռ�Q��Z�d�^����*J�U{��#\��r]�o��fiW$ú8���4&�
�T� lߘV � p��n�R��4���I��G̱5$:W\�yN��,hj�O�>UteW���ʦ��N��f,��7����%v��V8�h�p���f�w4X�1׀���gc�Z��|��{Y��m���0�f��i����ob5k����$D�����3ӓ �z���<�̀����%CF��zA��m���3(���e��b��p�G�����Lhk�Ë�4���S���>/bW�3��Uؿ�o�q���ʫ���H¡0�{1��	mp�!\^7�#GPј
on�y��[QY�ja0={ث�FC���Ѧ�4)PH���q���]ӁT	4Z�t��~�z�k�Sd�y�����a�����8��@��cSD�{��� ���k=��X�-r7��]O7*B�@�Dm�Ə3�(�$����Y���3?"bU4�5��"��tw���C���T���C�$���m
�/�I�B�y�����?�s�@oA���,�!�x�GÜ^֐f�"�j�O :�uU|�Z�e�BP0*_v��ݳ��kr/�>L~����|ua0��&��(i���1�ψ(�F�!]˙x����-�(���>i)w�ϸ�,p��4��M��З�$nFx��?�@��U��G�ǮI���nd��q�fԎ�����8�8�l̐��&+�v��<�p�һ$҄�\�Z>�&e3�_�����%\�eC�*���d!����ϖ5�B�P�ͫG�Ƅ��* 4d/0л4�ᖰ��w3עE���p�Q��7����@߰(ӹ�$�@��mW�<���{��J�{r}OkZ�R�t%s�2��E�/�W���؁�<�-���XN�`>�\�vş# ���.��ǈXHS��×������vW-�f���m�Ѱ/^�� ��Ӛ��@
���(R�<�ھAj�7ȷ�V�`@��M�P(���J�a�P3@��Q�~��Y�ZWu�#�h;{fx�d��{[0��I�0D;���K)�n;�+���8����K4*[���?�[n�S?V���x�ݚ��C��,�r,U7s'�*)
sǳ>No�?���P-4�$C�>�Yp&QD���2N�����‐(A�84�9�\r(�CU*�^*&�%�ɗǗ�!���߫�M�<`N��_V����	Q#r�� �s��G��nG�)�#�9��dEk�l�������XXڦq��@˥Gs��09�����Y�p�39��zGv� =�Ji�����rz_��V��w$��)�n���^�()Y|��:t�Ǹ�����#��(7��Y7��e[E�G��^[��jYF 	a\���q`QN("����xKx�/��X5��ᆤ��k�r3}q0)_������+u`�3�Z� O�6+.��|��֝�|�n{�z8�hC�G�8cؗ�t8���?��W��q��/>9�ܼ*���~���p�H5>�/?�v���Z���#�� tP�H���$���*��_�B��S���͍^��|3=�$��d��'�-����Й������߀�t��L��K߈#���y��Rٰ
O!N;�gn�jy	/�H����A`*R���)Iݒ{��E������e��6�4� ��Ѐ0� T�Ia;eg~
sE{�}:�+Ԁ��h�Ԉ�K����0|�C�]���ud��j��sY��{CNG�SN��F��.�}�3�SyF5GփA���Ȯ_�>�{�uk��Ky_):WB�D�"QB-�J#]���/��W�� qE�E!C��p+,U���*�S<O,�Y墵�t>��~и��gbP�iS�[7�yS�����<Ӓ{�>���.zS*y%Pz���ad�S.S4<Z�5+���9�YP�V�0PiPȲh'M��к8K��h�İ���k�؀Qu�F?>�9�� ���ݧn�������5:d�e8��u[R��n%�`Wj^[>�?JK���wo����w-��͋g�Y㙶D��{c�� ���^ )��P����.��h�t&l�c�)�m��+������{�)N����hM�1'�Ōx�܊�W��G�H�kݧ�d�;��b�E�e�{mq���	%��Ye���R^Jh�:�D���-�Bk`T����O�^��g�����"o|�:�%w���d���yɕ����t���t���B��	��ȅ0�?)���j�(B��������zZ�}D9��̳tuG&��**�'�-�$�/O�S�]�a�ܧ���@nMuZ��<V8��&L�\��
���~A���ӟ�Ξ/����$,����w�ل�H$�y�}o��y��nϯ9������YB%��� ��ɣ`r�R/N1��qi�{נ���<��J�Xx��d�h[^�ѡʭpd^����G� ?�9ӂ5��+�wE�ʎ��R�=�5�(�Y��9}']0f�QX�c K�)D�����,�u��N��j��d+t�Hd��ν�3�%*����|C�[��AS�v�������b$���v����&�l�b���x<�}�i^�r�F.��)�����gX۴�q(��5SN[���(P�$̳�p�򠐝�d��FRsu���