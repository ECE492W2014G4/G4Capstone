��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>��`HX����5a8Sjf\�|Vv �|�
���ۇ��������)��T�'�L�3*�51?+"�W������7���׷� Y�[�}nP=�PyW'���J14��qKxW�୽�V����+)Ό���-�o(��Q��`�`߱��H=%]�ȗj�u)9P��?L\�Y��rq�+W�||ꅡ]����Ҿ�G��=����`��	�*d��y��z����'ݤ�ֿ|�TI�7x\���B���挪}wNlR�p����\S�l����&Fǁ�`>���Z��K��EN
���4�ȸ��2�^������o��$[�5J2��.~��\N��r�8 3k�~E�F�%���p���:��:H�%9�χ�H��SHg�7Д[v룕�Ɉ�x��Z�S�9ͭ3u�.d/�0W�͛�B��U	�Tq0&Lxs�aQ|�yk��8z~d]j�V�}�~����@i��Y���"��t?��yz�ذ_b7)��Ar
���Bu\�J�9k?cY2* |��Jw����0s ��\�l��|IR
K��w���V6����H�Z�!���r����&.n��Z.�����L���d9Lmq\��%3_�E�ڜg�b��u�l���ez��"�4�O;�E���*]hҞ�b#)��9G)�H!rX�(���e�+
w)~"c-��
F��ݣ@aߥm7=`���S���/mŔ�21���%=�vL���e�T'T�8���j�p*PA��z��iob���o������C`��� ARR{�_���x�%�S��u/A�G8�Vf���T�Y2�����7�f'_>����E&��G�x��׍:��q�S�%b[�ٱI�W(y� �m>|��%3��E�t�|D������ל�r�C`~ʶ����dd���"~��){[[����T�to�Q�
�Ó!�U�x_��M�z�!����1s;)��<S.�(�T�ѯZO�*�������7F��.��x ��* eʿ$H�#3Y��	��J��k���N�\TZ+v(�U�);��{��<mg˖v���}"��F|Y�V����G���u"R�ԉ��g�Av�
$n�C0H�c[p,ٗ|�����e��?쓪jG�p+p�rif���>�Yd
�)���m�#���07fj�E+�'����,.X�l�� }����5ᆪ�{M�[4?d�	�S��"vW8ƿ��Oz�?N5��±4���?���?���$�N���B$�	��Wu��+X�8eK*�>>,�ū�i�q�ȗ��(��i8[-C�J�S�y�c�z5s���QA/�E�c��I� �O�d��0��/"� �c�+��8Z�����Z"
(�����q ����/E7;�@iY�X�^,��N[ �?����R[ذ�!���03����S.�nq��D���S��a��]9��e#F�%�����p�'i�$�e�L�Ũ_�"0C�H����-xX1�!��6C�x?^��6@A-~X�Ŵ@�	Q
���+uq4�J����pj*�B���l>T��TC<�OBI"On�st^����7��Zy�bBmM;7�	����5��Ǌ|HΖ��~IDEss�ML�~��c@����ҍ��+�)�M�]X����T4j�O�3�-+��B�F@>��r�lE��:V:yE���4���96�������Q����y�|��e��#x����b����-�?oa��߭f[�� 7)��iX��V�7�rBN��Bb�阣�i
|C�c2х��<��^Ͳ	���.H��we�	3� �����n�p<'��� �"!��Z����"N)��oD�lPU�ѥ�s����R � {�b��I*��͎�����CdIהh��M?������[����i�p�'��?ދ2*_�ߡ5�����`�I[�^�eɼ���4~�!̿��+��@��ץ�z��I��A��4�`��� �R긷:d��Q#�}e?� o;�^`$/@2YJ�5��;Cz����Y%6��V���Ou}���i��]"�(��SB��.�Ė���H�"({��Hb�u��c�Q^hPWm�(�jd1���ыٛ�A<X�,��!����{�J�szD�)wV������mo ���N[Q�[C�����v _��JA��L��Y�-,�$�[�2a����NT�7����_��ð�����=k����pN%u����W�x�$Tn�涥vUg6%�/���Z6��c����l�Z�C�ֽ��I� 0R�]���uSڂ�����%#-~�Yb(S���Y����՟�G�ѫg�'�O�����}������=���i�t�.�.nP�&V��=����bx¡ez	��&�FG�|K-��M�u|���(,��;�n�����`��޵9�LS�������a��9�J,5���	'p���o5��<)��4�\�d�mUuy��2�梢��=R8�vl�����p�w�9g�y��H�/����7�Be��B1��e�O�:/����Bl�RT/o�١8U���f��b>��G�-�j���5ƫ�^+�~�W���ϯ��=u����H�P���ָq�!�[��tuW���>����C�1~FICZ��Q��bx@4}A���R� I e����q�)%Èp�c� I���.D�}*@�|q���58��[:�3��>3lM�tjvZ�l��^2'Eg���QLm>x�)������&̅�l	0��b�e�y����)�ŸhΞce��Z���龔��P��L���A�.0�0�V���&`����X/�h ��>;�F�M�wT�Z�W�?��/O�k�ʙV����n�c�e�����Wޮ��o��IU5��%��40[��gՊѽڴ^�q�\��i�-���62��36J��>T�عV`T���X����7:Q��u�H��Ӂ|��2N���:+?Q�J��ܽ�����B�ӌ�Q����������#Z�P�e�K#�~N0��Th�Ť������ݏ�C���X
���9w���>dsAÒV{&�����X���L1���j0!�?G;��]��q2C]5̣��k�{#��NYf��Z=����{�AA��mT,�e/�����SaV1�NP��ɵ+���,���:3��J�a�О�^����?���TO��>`ϕT�Xu�����	��4�V:5�<�x%�$j���h������(v<�&��)V�����N5�F6K�>�M��3c0��	:��é���Y��9 �2g���T�j��8�� s�[�Ҷ�q�uh��x����)��l�hO0� ��� w]Z�O�=�qے����?��5��-�4kB��#ֈ��-'�ۼ\��K���m���u̐Lt�����S@�M�	aN�e���y~d����b��\j��|C������{�2ZK��!~�+�3b"�D����l��#������7��%����J��X���#ϣ>^k��?��<���/�/�@R�0��'c�.�`�j]��ւ2�p}�)�~�u��Z�2��p0�f��������32����m�~;�.4�������C��9��j�[=���9W)r��l�����KGbp�]�/U��x'c#] X5�1���TљE>�D�Қ�g������|_�D�8v(*[�Ev8�݋�3�M	ض�wɬ�����\�@Ң�"ht��T���unc3hv=���׺aЖ-ǹ���Y���Uם�����"�}%_{���t�_P�'X��� ,ú�n��/~".%+]!>PL ���9�d�	Q�R�	�+��I���#$��.���]^c�BY)Ũ�g�|�lm�NjVSc7|�
��p��7�L���9���ݖ����RA�� �8��B2o��nQ�D`A��1�2C�"Dɹ�Ax\�q������\pfNW�b��%���oz�!+���;N�"^�2��<�^�vȗ�^3۩���垈�m$�L׭0�Z2���iy��g\�b^��缩���+UMv*u�3h?^-��o���Z~��mtP�X�6N�V38��3Olp���T!qY����܆�Xm��1v>J�@�w �}�v҅�@�d޷��m�kV�uS;���m���V	���.�(��#��}��zw�2�3�$��#�j~i��CP]���:~1E���������^�!�dK�H��"��43&�ג�Ϥ�4=����JA�-��٭�.g�6���[�bؠ�3D��Yu�#�3�x�Gx�%%~E�u����i�aX���ɫ.r�����lݟ���ڕnS�����u@���IB�E��^6����r# o�����a��ܼ4����J�����}��?��NN\SZs�0ww��K�y�v .)N�N�0�w�b̐z#��g����W�(��$�2_h�0�Z��]���>�j���Kq
?�(�B�K:��u������������	p�K}F�g�j�F�Y�+e^��+���ݙ�w-QZ�	�@Q������X]<)f��;�Rz�3�\��o��9jYEq�n>Q߻��*�So�;�k"��=��퀤Œ�� q���3�:/1�x+��O��ξ[�L?�b����lEty�Kӿ�7��;��i��$t\�-�I���vm�̩G+i/;s�����@I��>:U����bPu����,�� �Rn�7�p�0�2�Q�˹�7{V/U���*�l�)�$�v ��1�����@��I(eQi�U���Ck&������qo)j��e�p���1IL�f 6"�����2�R�]�����Z3(�8U=�q�u����8`���<��k|L�
~��	�&��c�K�{�.����&CK���,�.��~��~5}���B�3�'vh���y���G��3�`�2��Y�ϊ�,�w�Ï�g[-���A��?<f�?��4�rj>v�e��Ґ�);�<�T�E��8����>��	�h�!�	R�,�wx�#��h���7	hP��A��>��?�Dl�SsЫ�3ɔ�ρ2��y�~�������bj|��@��(4��y|q���ǥ��I��,���\��3����.!f����6�<S��6V��3�����Һp���m+1D�{���G�;h�L�N}�Zlx������0^]�0��H�Vö������!+a����Oys�T�%- ���0�I���ű��A���B&9����dl��i���k좧q�7ڇ�j�j��NcTvr��V��f�U���C2|/S�Y������2���q��H��m�k��JP��²�V�l����!&��XQ��U%�>��~@�Kn"��s��v�G�O�I��M�73U>V-���З�#RS]��ճ�?j�"G^.%���7ΌKȌ��%�y:5B�5�d��<&~����=�s<Y��X��M�ٱ(�r������3[d��
��*i��6e�G��Gʁx�$_�wǸ&�xQ���Ru3)�Xr(�O�8�SR
Xf��*�#�'����r>2�9�W_�A�D�z]a�)�Ͻ,Dh�4���FZ�9����#�%��ǚ<�S�����5�.x�%e?�x�{��A�L��ж>_�f�Oma��ںr���C�"�T�U��^��N\»7Rۥ og�-�i3P�'a��PX�Y��=m$�u��L��bB�U�C#%�����'&�6�>	�f��komYdUӬՁ�e�!���~%���SGZQ`a��O�{��I��졬(�;@%��"`�8F��HyjG���a�v�[-�A0����@�"��#
�(��[�RgC�Uv��ý�+3xz�~#caF�@�<��'E��p�cy���p�a����Tk�$�l�]N��4uHq:�@)z#G9���wk�F]!� mr��cR̋��I�dYXvJ��7|%b���(�$�\4$i�#2�tP�Ȏh��GH�t�/��?�%{�������>�ē!���7����_܅Wm�]�(~�Ҹ�M���/[�__nƓ��$�Kn
l�rJZ��^�V�&�]T]!=N� Ml�I0vo�f1S<�6�`	V������S��7m��U]��Ղ��P�5�B_�==�3PX�٨��X�*c(�E����9s�!���Kf���Y����Ҙ������ʶ�����{�lM@>̈X���L�	a���'�ҸЗM�A�� ���ߒ��_�ryB�'�q~sY8�Q�J<ӟp<������*�:����-�O��*UVv\���Hw9c��RU����4���K��B�����9D��od���4�;'�M�%�u��h��ôn>8_�0�9s�өX���m���iZ�ޙ#�1H �����g8ʙ�ˑ5�+1b?^9�Y� �ftbZ���:Y�x�*?�;�h��+Z0A��v{�;\��m7�o����m�ٕ�ة�}����zF�I�Y)����)�m#sd��%On��]�)�Yy7��[�����YQ���P��`�\ Ĭ���ox�����f���H�����QK�d���6��G�td�q�����wzs0��|{�r(�e�X�2A%[8�]仩�"n4���ŋ 6�
^�e��9!z���C^�b��Ax��Klg������J}��<c�d+�orb�ɮ}fi��h�����k?�j����-��EC����..�k��:R�
�A�ȷDJT��X5��`I���\���7��|�}���)����3�|bLo>-)t�J?�(���9wzP���U	�|}�t9�;Am��gR6�G]�L�U�n�"�{����ͧ�LR�����+WB_� Fo{"I���[�g�\�����o�4�7i�B4Acs���2�Qe7y�ˎ��ۄ2CRCKa�2��l�=s;���m�KST�?��P��G{����O�s��#:~�����=Rr5���'"������i%�G 闋� ��W����vNnE_F�w�b����[8B�{��Ϟ���:��u�;�2����i��&���
���4����JC�\����`	w-���۩�_� /0�D5w��l���ust��"g�AM�Լ$^J��7��T\�կ���iX�m�/��;r�q_燠m66wC���ts��+d��k4����4,傢u"���!s0_�W��j�WE��!��o�'�xJj���	���_��u�h�x?�ߩbŗ�++$��1fQ���U=טm帠Cu{�.n*𦊶6=ȦTd��@,��3ȃ�=৛�/���r$�Gʰmt���-لv0<װ_'�ٹ"u���*m����*ip���;X2sNM�^��n gx^F��:+ ��>~$�j�E�e�RC�.���u��0�aba Vd	I�6#��B8خh�����K?�^���Dp׹T$j
D��[�>�m���=�br�n��̅�|Ӽ��ղ��4�i��(!&�D����6*�_��N��)�
�ti&�3�P�-����X.�R��QCe�Q�3C���\���&� �1����)[YR ����Ř�ë]����h/��%���:�3��w���џv�?Z �j���}2x�4���\~�@�����bRS/=#��fܐD|�Et��۴�.Fi0H�}�0�\���	�����}���67]�w���Ҷ���z�Gc�͎��U�>m
"]*�g7��_�^����;}S����	]=�x�y�+0l���h�4~�^49�Y�󹧥봻��/t�,%�<� �ɺZ�"��(�z��u�T)���g�֭��|��6��d��Ůu��|n��l�-N�4�.�M��p7�L
�u�D�Z�u�1�����V��{:P_4'�V�/�܉���יd|��1�9�5��{�u�\e��6M�a��S�����	��h�i�C`�NƙMOw��U��20ۛ+H����� ��r�ZBV�D�u"��9����HD �-�u��w�L_]{���eo����=�yCH�c\�>�2�|RV�����7�%A����Z�n��Y��N;;Z��6�5zJi���������Su?X*�g͛$u�?k3���?�7��EY34�%��a�ڂ��;_����I����}9�{�9:AO����- �Y�pY�|q�j�r`�-����5|�էeKG7���P�A�Mʮ�LY��M8Uˀ��'T�akƮvOզCC�t�a��qxSG�0o�O����@S��E^�^�-C,��؆����D`nJKl]�S�$�/�%��ft�K�)-�M~@�ln��C�+�i�t`�C�U@}���9�r҇��.D#��H�|-v��@.�w��4Lq�zmh�D�|��lU���O��@6�����z5��S�C���^�X��}��K�;��p�gM�D`�0�h��(IV��/�论T�P���<$���PC��ux�ɽEE?��w9���ڏm�hS�#��ָ������x�$a��z<�z�3S�w�p���ҥ�:� ���Ju�"�~f�c�	j[�a���;����_�tɯ��U�t�|I�rM-�	��ua��x�%J��A"�<�:��&0͋���|<k[ä�"�D����pku���~�&�� ?�;��-�j�&�ni�7����,�=Lx��[��K���,xQ6�[�F�����3����� �K\�?�u6@u�q��C�I�':��5���q:0m�W3��"��-FZ�aP��
��t�օ���r� I��c\��#�ɍ� N�����}�����K��-7�ϗϢA��x<�`xC�7��$� ���S&��<y���d�>�ޠ�gb���&;1� �f���v7Y:��(��a3Ҍ.i��{�yE��đ9���}en7f,�<����	��Ш�[�Km�1.|�(�w�i�.OM�I}s���ht�c�D����v�K���=e�I[�v'K�ws��)�Z_߬��@@�S��q}QΘû�7��l�\qx���qI��S����s�� ��KF�6��u��w ��;�ɸ�#t/� �����4+��E��߰�"���Ԏ;���
i�*�@���/��H��P��ٟڽl�e��I��}I��&74�m�'�n��ƒ�C�y��r5�V�����D���I��}�q��O�-��&�@��D]���?(,n����w�u;�"'�/ i��!�Jѳ�D$q(�7jCB����mK~R����J��ޯ�����58BbɈl��~5_�͂����Z��'v�#J�"2� �XE>���Q�a��]m�w	���u��#�k>���1�J���g{��3HӉ���i<!���Ĝ��^�~��[�/�w�t��eiz�и��s���(#5�c��Qi�9���@��V�p���
�	����5���ʴ�ܹ�silْ�3m��uF}��j���%���_��֮4�õ\Ϛ#�:y��g�X�R�F��ߐ��@'޿�Ph��:���W�t��A�C�{r~ʊ�"6��� �~|��[���$�K^�;�����p���+>j)��0+F��L�7yA�Т$��٫LnN�@�����N��������Y�h��L�LI[���vr�P��8=�22���,?��#'��&g�o��Li� �3Z���:�!�&J�&�}Kz侘�T��2F�P�h��r~'��˵c<R FS"����k�������8�|�X&��M5��C*�3�m��U���7�t48ȩL��8�p�N��' VY�u��ݞ���6kg12N}7����l�Q\U
z�Y����Lq̸<�c�ÈBo�h2%%�Vmv��G����O�P>E}NR7H�_cP��f�z+�pj(��=����#u��"-%�`i�NE��ڔ<��#�h; ��W����c2���W��`�2�iL,�#x��	�4F�|r�s�v��;���*�D0�N��x�0�][��}��M\T�OĲR,hkH7��F!H8���%T.J�S^8�=S��I<A������d'ycs6WҘ��
��5���a(��Qs5u6����F�K�L�N�T�S΍�z+Օ:��%X��均|�}Z��n�~|�C��j2�a�v��D@#Q��tF`��h�]ܗ�q8��3��=o6HN뙞�^�qVx}�OHV��I��"�G_F���*�z�&�m��-�����K�Ι!�Ϧ���.����!?��8��$ش�P�FR�}��O�`�Ȓ��Jl
`E��Bm��p�Y�2��}��w���C���86���uf�����!m�� 3'��N�nN3�%E�� � L[k&2.<�(Q�[����z����Y�W��ք�q��&��>	�C�"Qoй1�o� ��8���h�g�[$�]p��� B����O&|�W$���]	�����`�Q�U�|��]���n�� �v���Z撶����?R�G�~���1
0�څRP!�+4� �v�D�eW��	S����[YiӠ�	���@�<���»b���8���=�_V1+�9�tꀴ��{��9�Y:�s.Bz���-~5�u-UrH������p�
��r�����z�K��=ʐ�v��|Wr���'��#lE�s;|�;ȕ�����g۩ C�EK}�V80�m���YV�^��N�%v85]��6���u���˓