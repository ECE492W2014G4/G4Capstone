��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�"��F9s�`&���a�oq���F�g�O�]�<ݲ����eCL��D���{�5��8̝DFI��Zp\m|Q��
�}�6C���UnF:<�jΈ�2�����<����sf�k��,jڙ�����2��X��Ss�HL��	�������+g?���N�Ż�����|�v7�{M��VNB
��Rs�゙�Ld\��X�'��R :�J���^�����kMkx�Q���3!P}�e���Z�Y?.�U{�RP	�)��lI{tI(S
7ZF�I��!X3�.k�(w�q���ⓟA�G����Қ(�G�0�H˝�u��8��.�J�U�S�G��{��ʓ�	8ycn�����e�6��X��嫎��X��8j}}�Db��+��]n�
q8�]�&�G��s�-y�\+����u�~��W]ż&��gC��u	6��_~�h����ܔ��F爫{IA�tr
^'���8J>_���!��c�{������w	p���z�Yl{�S#�3ְ������i��7{�`��L����L���1F�K��A�����H*�G��0( 7<��L�(�*�=�M��)n������!��Zc�:��"W=~�~�T�8=>F3"P��
 ��Z���IL�v7ņ.,ko���X��>A��ϑ�`�-�ȓ"��|�=(fqg	՘'�iK���t������n�C�����Z�p䱼���R��DG��H6͉����;.� ���\|���"5�iHc[�pI�ٵ|d�{��+JvR�ev��>�<����n�8�߬˕5T��*$Ac�0��g����>�)
�qk 4eƯ��Ϙ��$�)�5I@�oT�����J$Z={����1�����?���~Ac�
v�'
*=Ql�+�w�aOB��.���Gb҆_�����|���z�d�o,v�2�Q/���@0JX6���l��VD�$C�$֧���+�Q1��kcD��Lc���>d�����Cr��p��F���'Z�4F����@A�YK�����`�QwD
���?{�\�ɸ�a5@Ʒ�©��4/��]�jm�����ҙބ�rHZ?^ͭ��w��j�I	�g��	Z��K���^��K�"y�EX��zm�8y�A��4b��M`�jq�N�EZJ�Q��ھwrlR���Z_���m4$RI���#�EY2�sʪT�5&xq�3�B˹%��!��}�LE��h��陟k�)z'o�iU�����v��`OZ _�0��J����7D�hQ� �apo��B�Yμşv�dv,�]��H��8�R��(m6Qi�^�ٱ��DC���t@9پ+!G;�/}�R�Z�s뱷<�?�p�`��b.���(]�,MP��������5��l���m ���j��2��0J"�M��"m��zFN��f�˺���Dq"{%�
8��V%D��L�QJ�V�X�A�Q�$��"�J��������^��I�]�ZOo�si�dIS���Z�|�p�r"yrJ�<��1y�}�whΚ��<�#4�.��F���w�qל�Ʀ�?j��<Fbi���>��3��+g��+����	,m��[{�d�e��f?��(&Cj�FPp�T��,�p�t3Ď�'N�"�����A��A���V6S�`�8�
��>�p�����5Zxc��}�h��V���\���۲:����͗D�����U�{��-�_��{����
������~�,P�\�Q���R����`���o+t����|�8�7N��r��~� ���i$�t�*?��(���D�C��V�L�=�us�������M
s)�4:�&�����ыS�Pe������Ѕ9���'�{G�^S���Bs��X����M~��f���sgǖ!������lʴ�#�I�����I�K��[��P8��"4�:�����eǛ3��Js��e�ϋ�v���%�(�i��K_��\6�{��^(t$�NnB��@�7{D�5�$��( Z��F�9��;N
Ց���ɫ�Cx?��}-p���s5NwX�]!qB��܎�w�{�4 �E*)oz]ߘ 8mn�;�6�ԙ� �������t���Y��>c�A�WP'���DB��:����Ē%��"���J�I�Dj�Y�5�� `B�R�߄����5�q���^R�iR��(�Xf���)u���m�9�+��q�J1�ۄQ��*+y��ܣ4��<���B՛9˂��b���� <�L8T����f��'�4*=�Ogi�,�t�jߏw�H�\\�P~�7�`�dR?	H�a0�J�<���f' (7��ȟ�%`&,k�)I.�k��p�>��:q���/
}p��k�움�5��m���&���/ȕ�����d��ذ	����>b�ht���Fg͒��g�N�\�̇�r�3��v�'
���v�[r�>.?�侞�{����+Z��L�J����'<��*��uQVt%�{�gd^̐��"��7�����"�C^����X'ی �5�oX3=���s7�ܐ� C$��Iڑ�C��~ğ�~i�!�ʣ-;��JG�ٶ �9|!����A�9An������3�1�'<��J}�]?�T��E|.=�m�r�|�����0�#�O�kQ��ZwЮ�����&h���������4D<Tcݺ@�����n��'G�S�7M�NμL|��G����`=L���gJ��W�CXG	��2���wt��E._^|�$`Ŵg�+H�R/C�6A7�bz�e >DT�L��	��,9�Xm�����7i��8�'�u�'EI���Y�uVV����G[	�5D�P�cc&�������������{۟h�o�ʽ��@�n��:Z,(����i�+��%�MC=š�x�N%��E�*94�F^h��H������G����2X"J�c�A£���<P �I��m"ϰ��>� ]EX1��{wX�`��%I�l$_ܭ��vi��5��H��Dԛ!�p_����gqc�{���yƋ�_�A��H���T�v#f���e ���&vG���hN�����xb�������2Er�����I����F����ID�ǘ��	�>���I�~�SU&K�܁���Xg�,�EK��x�(��}aw��d��F/Z
R��.�ʗ'`���w���+������$t�����!�S 󔔷hl{q���w�7��}��^�&Α1�e�̥?�&�������'Z���}��7�"q�,��KU�S�:%q�u2�u&CL�Z�K��^���鰄x,��	]�5q%0Qp����4�p�)���<�>�-D$B�(�=������΄�j�d-�e���"�W9.K�
G՝��耤��D��bF���^��c�^�(��	R+�c��=;��4�s�/��v��D���$�4�����*'"R���ΞE�,���R��Tx,ۢ��bD9�Ԍ�,0���{�WDw�H:���l���ָ�݃O�埚Rkg�h���ϊ�v��E�Z໅�mq=JjLɫòĻB�E;�K�����U��mm�_�G�^E��H�T󋍷3t�l�t�6�^؜��;>P���'akn"P#����|Ǥ���؟KQ�f�2~m�h��7K�)A��=�t�n
�6�:<��޹����k$ϔ��i������	 ����q+U�Pj)
�.KS�[��K�+e"��C+乮ďGA�Z1OYQ+�?��nϮ{N,4j�i�L!��Z`��߿�����Hn4!��P|��e���r�#.e��SvߖN����_kő�4�l;�ٝ������(+_3I��H��mC*ڻ�P.�C�5�\Ġ|4v���4���U؉q��&zRz��Aq��+z}��f-���j/�T�\�h���̘Ơ^:�/6+p�LX�a�2=6�=�'oKNJ�P��P�O�Z1��!�P����i~��i�%f�[����ͪ��7mA��nm�X}p��I~��;F1z�ݷ@��r��|z���Q鸰���<��j�����3^�r>V��K�����vR�[�8��PN�n��R�����������2���kM��"��� ��̐d�QtvK�Z���^�܈��g��n(�R%'�QP�:��m��]���4�+�*�g�B�8"U8@P���չ0)뙮p�:��H�;H�t�C	����:��h�t��W3Ni�N/m����$��08ʳ<YQ(�
bk|T�0�Ԣp������AZ��Y��o�g�:G���ii���$C��V�8���,�D��x|�z�����sԿpV�9M�����0f'gj�|eox�����R��"��(��Bd#\A�E�v�j���;�ϐ$��?jL�@�i3�I/YϘ@D��������&K���/9�[�*�H�ʐ1��G9W������A�U��g~ ��X��]�6i�)������fT�^y�?[���̽q��a��*Q|B9B�Nl,ٞ�������jx�X�yz����Wu�j��\2.W�MDJ����?�O6���@ll�$�B7�Q`P��ˬ�^r%ɟ�R�T 	m�H��Ys> �r��j@X�7�1�l$�!w��))MLMWZ_�J�W*Zjd�����C%����;���߬f���	�_�/���C�qJTH+k�?\�r��a��fpq_���d�`-�$S�K�<U����}����/P��`2�R�S��BV��$����F�h�q�?e���H�CL���̚��3�>HpuS�3L�Y!W�V�>q���BX3b���\��c�Q�#�ߛ���V���KߟA_�����p��G�cPW����+�Kd���hv���� ����Vڵ��˹��hn��J6=dUG�<��u��$S�<���\	I��K�C�aϴ�z>} ��+��p��z�Z*BT汬x_�������L<��`i2�Hb�c��m]�`�o�AB�����G̬��^9��i$���+c`�+ZQ0�j�G�[Tb|*܄YkV��C�X �7�ֵ��:�o�->����U0�k؏�o/�Jۘ��-r-�b	�����$���L}�H���̌�b����Rqc���B���cB�Y_�aM�өt��eX�T�BS_q�q��]�:AM����R8��_��
��e�k�'�r�u��/���#蔈K��J��Y�6�*~i��Qӭmr�;f�+��C�ӭ*�\��2(�%���}�wҧY���k�g){��p\,�<`\�j���j0m�x�z��֚�ʒzL����rr�����q���2��dEY����I��'���ˆet%A�^Wz����S���s	�|��HV���5f�brϑ���F�s
�%��gy�mTx��(�`!,9��o.F������n-�9m�u*����Pd����-^|�X�n������^��k�� v���W��Cx$�:(4�"���=eZ :�.���v	�S��U��ދ��`�X�{��EFHan-�B�[�Aċ���:���C��f �ce���F�@�痴��O��'��pL�QVHէi(�R����Y�����y$�M|� ������v��%�T�\��|%j�&�Ug%ӮGH;�Y�h�����@�����`��j=�+>�8e�����3TT�(������+]��Odd�4%����\%<��|����Ǵ]k���?�j)��"�$�o�|��&�����Ef���S?��5��^��n$.�V>�2��oO�y��d�e,>j�.�![ �4�b�(�c����.8����J�({��E�U��=}�4�@Һ�{����YP�,�:ds�tK���*��lY<3l~�(@�-Z�l�Y�mH�Zł��9�7p1Ix���F�p
}�Ay��'/Lq�Q�ƠusMʭi%PU�E��@{3�^iu����t�n�d���4�4f2��T��Yd�1�,�D8)&оf0��
w^`��-�`F�4?��ԙ������|J���Q�g�W���(�|z�B�K�%ԙL��ъS5�|�@]�ڎImI�@���|�:>�E䊿�s:����r��#���+Y#�#_��sѹ��[{sWG#�9;�0j	�:F����ۯiU�R���q�����t�&W���w�Ѹ��;�����a���z�Ǚ��|-u�a�c��a���� v:��X�!�{)4J"W�O���B�cTn�~*ˠ�7����Քf#��n?����q��+R � ��L�{@���h"M��j��!���c�0�Y�����ZS��&�ÐYي���qY5��X<�v��� c���̀6��)��0Vt�jǨ����Iؑ�>W�A�$����@�ЪѪp5�=��W;�l�,��8s��O{i5��'�s`g��x�ٿ���pB�e�~��3�[5���>��O6�W �u�x�僾:����v-gl#�'i��%�d���zi�$gmD���b��|�ʙu���k_naL���۶��'4����X(��Lp4�|N>%��9;~A�
ē��̽��t���j��}E���%���:��Vy��`����,ӣs�Y�3�ȌJ��;c�8�L.�R������cfo#��������2ޛֳ�3��ܸy��nXOQs�̺��8-�Q��3���{C=����Mˤ�6Oi`�ξڽ%ah�3�����#	�k���V����s��v~�#C�
x�:m�1s��,)j\��n���^��O�i5���/�ŉGTt)-�����"����V �N��x3�#|`].?x�i�d;J������&Q��#"��6���|(���9����o�����B@��󾃀BV�F�n�@�Z��8��E���B��P)F��HY	l�YF�`�Ω5*ecm(<pM�d�&�-�ti}��?�0��%��԰x�{�y��3�QJ�����HUfy;9@0����>�)��}r$��_۞����x���7��ؗ����]H��$�V��E�ů�T�<-6����d [����
� 3�W������2m�v��7Z	|e�)��5Z�fX��m�8����J��p�w�G�dH+���.C �^�C�5�:[	Z>#��o�{F׆&��	T�}�a������g��l�&/E��nI)��4�H<��*U\��eD��g;�+Z����C9��p>H���_D+x�� ��ok�@?1���?1���ݟ��r��i��[�H�@�d�"�h�I>��ݴa��
���.�H&N�%����~
b�:֠�34����@u�_��OU��S�#>�g��^�
"@��o�J�OQd)n��I��J�7�S�J�ǌ���R>k�%�X��<Y�����2��7��|��h�t
ӛ|z̞�v���p	��S|�J�ZP=�5���,���� ��%N����:�^�8�87DA�Pi�\�iLvB0�|�TܫU��$xBT����[��B�eQ�2������;� ���o��^���_��'W4Z����`
�)��Xa��l�s���@ӯI>k����X�A����[�D�B��j^�
�\��:Bh��&� a��F��k��Z>0�fW?��t� bP�l��w��(Ѳ/������b�A�)ȋ~�(q��B�,3��A��o�����@���,������9R����2^[��!o>���Q~4��e����|�8�0#7G�;��z����bH����-�
�������e]�F�u�KF+�(A���ZJ�¯'�D/W�7�Tz��Yqy(k}��k�#�	�����y�0������X�?��e{v�R�t��jg���	@M!�-{�Λ�a�&� @�m���ړ�u�D�uL��c�W�����`���!F�:IAID���#�q��V`���m����r�lb�L���s��:��5��GU�M�Z�9bq�`�m2�*ה��Զ�oo���S�&(U1���!sx���5�XqEX �3��-�g=�	�@�Q,�&:L"ԩ�JG��*h'R2o��tܪ׮ �^��f�9P��[9��z���V��:�F̣�b�D�e������\A~
�\t��iB��s"9YI��5�v>�bgig������@��deلwc�*S*z,Y�2���N��pUT��I_]��Onx�U�B���]hEc��C�M�� ���/��e��0�B0T�~oe�[����iYApUJ��ٷ�s�l�����d�`+b�5�y�_n;�Q8�+��q �#�b��N�Qջz3� ˢ+���1�^EWvF�1C�&֔HN=���"#s(捰���&q�F�s1K�7J��]�L��?�0�Ek>cz��S��뻳��\6\%Ȗ$"pz��7E`��a������ű�]�>�b�kZ\$��X�dobv�ן��ҏd�y)cC���T��!Mg{N[W�sm�3�p�椟����KF���@z�����p�,�l5	�yO߫|�b�ܽ�+��g�ڛ����е�K��"��28B�Q���SSmJ\ד��n������X�F��x�:�J9x�`󤫈rƔ��y���-:�i�ĳ5�W�!R�RCF���mu�C�S¥�0�>q�H�ײDfdm��
��SK���o���D�V2^.�M�gUF=P�q!ԡ�.?�,�bS7�q�00ӈ������[ߗ֡{������F}��@��x1Z�d2�E�����<�y�؎�j
��v�U�},���Y4>Z�"q�Ȱ�"��z:������U6���:�^�b��/>� u�f��(�F��M̋Go�i�PL�Uu?T��\8�)��=�k�Ӳ�
t��	6���F|���M��x�y?ll�y܄�˩��Q���ɦצuG���� :� Ys�a7>�>��,���ٗ%E-kaI�S�#�&V4�a����,N�i���aH=�������д�-��f���k!!f�8�r���3T�sZ�RC�e;��v���n�F��
UGN�]x�Y��H=�J~��މߟ2^! ���P��䦋Ĕ�%��n������Q&i߃�s���-�Y��t�@������Y-Hj��o�#��X�&擒^��6�~>��gVT��[��t@*Ƈ�\�c�vA3��.�*�ov���\`�=)�F��t.�� )�Θ�|�ۄ~.�-�А,���D���\���&�)���_���-����I��"�%a{�k�k<��?������lISⳛ�ۊ�=%I�9�A���7婏�
Qe�����dj�&H9�U�FbV�bs��#�2|:��e@'�Lۤ���+�H�D9_�N��rzJ�E�1[�6&g�|0�0n�wc�K�G\�ۤtE�q����#�,P� �����<���%Z6O���d` � ��PYq��f����Z8���7��eI��E���yXP�'�e"�� �I���ᑲ��<M�o�p����CT?����ܖ����n�̂�,��a�M��"V�dv7R/�:r���NYe�jI$\j][j������c[���<Ab��V�}��\����I'#�+��j����L���MG�z�1/`|Q�LG�zT����(PĴ]N��6k+}n��G��A��Q��sY��������� �Ӂ�o�G^8{�o=��T��-�����ٯ�������]�������}d��l�vdXp�:>*c�ǜ*|���hF��\�U��e��QS��
��!������4�k�$����� �C/�G��Hd�\�#}��U�?k��sV�p����r�d�Gxp��5Zs�]F�3L���F��3n�[��0J�˓�rC;���j�������鐩�TmS�M�[h$��>2�g$��N��� {�d&;��uݸՉ2�$�֩�$7%���i2H��	+~��KV�A��ػF+tZ��&� Xi��u�W�� ���
���@���$xc�q� ;�6��w�p����p-"`����@��%?��2lp�Oh�}�5ނS�(��k�r�ajLf��G���3���y��`����M�6�`�����N&��)X�``sBT�ZVe���E~r� �������`2�B�$U�.�/��cy�u?����\X�c��i�˛t�ѝ����}yD=Q<螄$�CY�1{�ఞ��y;���H �����i�؞h��� ]?f#$���!w��D��-"�\QS�l���&��D#�e��*����?��V��X�W5Л�	N���Q�f[xe�&<í��r��x� a�Ul��&�`��x���B��=�P���Z?(����!�� Տ�Nj��"8��2�w9��m�3�j`���T�g�wظ's��
��?���Du��&�e��4�"�"2�Kd�ܥ]4��g�GS�-|$����g���᯿>˔�u�L��`w�b�*d����1��x��+�y|��50	S�Ԍ�t��v�ϴJ�J�i�:S^2ZL�e�Pm�<+i8�P�����#�%���5��8�]�/D�XtAR��:�]�?؏��Jy�H䁂Ϧ9���.�j�\	�9_�o �n�q��k����c������D^_@��`y�����bQi9NE���l��6|��gJ��w���m�}h�y�2WKg oe<���>�|�� �%�6���=�D�C�5��v�=�;b@>�*��yT(�r>\���D5�.�A'Ϲg��,m(*��c��~�鹐sL�7x�w
�kb����n��������t\8��Bw)m�D�x���l�Y*1�"ֺ�9�hݗ"����:}�uG�)��&��?<L��v��9j�?{��̀�睾B�x�pI�+��K�K?+���.;��J'� ƾ��it+s|�i�<x��X8��*@���6���9���F��`�̚�V����p��0s�5�W���x�f����OB�K���b-hE����nD�n�!�쀁�Ð����ݙ��9��f��z�~�����	yuqz{�C���X5����#\���]KuB��H��|:���c��*	�떯�Z�I��OW�m��w~�u��7ʙ۾W�M�X��EN��D�F����u)Vx��O�U��E��l�O�:�����Mʽ��}����N�%ɑX5=�u� A�wn�$�x�t��U��®�R:�f��h�- �(t�Z��,?�IՕR��h=<2�Ss�B��t{ӊ>%��-������~(�y��>-�Hr���g�78vE���#�WBwx!������t\���E��7ou}�.7��8��:j���'7�-9:-Z��&��K��R��Oy��67�5.,�rC a�~v&���˻�N�I�}�[��x��q��"W<x�}P�,�|�����D(�Yu����B��Q�>��-��dzO/H9�X�4�Q_�S�kx����5��и�ҏp%`�I���>`���s7Kp�t�+*���$<N�^����sG`S�"u�8H�AygmX�����*�!B}�lÄ�klt�	��m���vS �s:�s�3�����4p�Q�ó� M��t�%`��B����GGf���!�p�Jid�	�	�ֶ1OI� �{�VUUe|��eL�jI��42���1�e��b �v���̍��BoW'K�ss䖝�$���%������w���i�.����1;U��c�.�b��$N%R���!9���Y�,�/(�s�x��!w�t�@.2�_��ۗ���B��|ۣ�<�v$��Y�I0v:��rQ9�m���}ŭ�MF��ЃJB%����@�>���"��f�w5ĥF��C����'�]��P�'՞�N0x������*�+1��@Ǵ���"l��&�F?QkYW?�!��ك�t�ێ`G,��P�N���E#�I#��]�g?�X��6��[�>��@�JS
��!x�쬘�0�M��9ݭ�Ŝ����|����Q$�iY�ъ�7R��W�<�QvW(�1�-��c�za��S�Ƶ+s@��d�/ynq��KT�N����QB�6Ռq�ߜ�����I�7N����YQ^,/w��&�N�U��������ԧé�CPl�'���_�Q���	�g�dx��U�p`\n'���;3ӹL���;��P9NO)������W�k�,ǰd]�U�k�ͻ�u'�3ٝ���.��S@�ă���r= �r��h/W�F������,���!���πg��0��tc?h�]������uI k|��R*M�x'����W��w��EZ9'�O3�s;�\j��N�_�2�#�I8�ctrn薟��B�ceM*Э�KUv�\������8~�ҊG8�Z��,�>\i*ڈ�%��*q]���6��;�SOM��r�����I)@�Ur�5��JO*����sĵ��O���?���tJ[J~ǷgM�O"��8C�[jN�FC�9?�B��D�s}����j��dU�q��>���,	M��VR���@`��Ϟ}����kR4X{BT�@׻< `��à�{c!��Y���:��Sא�y`�q��d��$�Z����D�O���sMO�����������P
�*�o�w��(����m������l3�n�*�".�[]7h�F�im���Cܦ�p�>0K̈́�:RZ��h���4�0��� r���*|p~Y��n�bIsj�&}R]Q���/�
i��5:�.*OtM��2�;�5�� `�r{Ӹ�!��R�Fh�Z�R�l<�Dr&,EM�0MP9I)5+��+� �:�&�GmNà>�o�T�l�r m���!�1����<��{�.!?']Vt�l �B�tCIT�nk��4��}�u>��s�/d��䧙�ݻ����������Dyɬh~�!~y���靦I�%YW�k5~��y_b
��F��k�zwŪ01�Hw���w����hN!�`[_Y�ZB�?�s�Kq���凧� �&���Ǘ��.E�t�+v��J�>>�%W���ަzq�$������Sjh&�D�d�Co'�K�V��7�De�s�uV{o���P�JKW�$�Q�c���mao|����=���1�=�
���[�Fn�쬗q�(�io�W$�9h~.����4?�
ڢs�q#Bd�����Ƌg�\N�V�����r�*�l���9�kףxmEDK�'m%��h(�������1�r�x � �OIFaZ�.K��M��$������V��
���4��Y֒@G�0Ym���=z����z~Noݑ�A���˧(�����9��T����rLU;��@�@Z�������W��'�4rd�������tD�Y��s�0
�=r�<�� �R��5ǫ>;�]��.v{�xZ�n��-8��*��B����:��Մ���#>d뎩 [��x��s.�˧�c���=���0?�@�B��O^G�]��N�'�!���)�o���7.Z�F��
�]�翭W�c;�B�Auy�_䐧��$@�+�jd"����Υy$� ,��?�X&I�sF�ٔ�%N;�k0|�)���v�=P�LO��>L��7haD��.��h�H�����V�G�u����-Y�G��b�	8�Ğ���Q;�u�� !��gFj� �Ȉ� ��Sm�x�Jt7�i'd)f�j�x;�b���md��_N���-ӻŇ1���������	F:��۸ Ⴙu��˔��2�|3�`��*t�'����v�|���I"��~����G�g�睿tB�$����z*_��x��;^���	ԝ�<I���ï�	��+&�l3i�l�7�;�ҿ����R��e��m������k�g5�	�E����&�GF���o׳��������]�9,̴��Y&n����Cv�C�$�&y�܍���K����*�xH��X*>���!s�Oԡ�T7��a����%�O�%�� �0.j��8*6��g��d?��E}�/�a�a��@.�g�����"�c2��[~ܛ��hH��,�E/� ج%=���K�*�Ѓ|'L��p"�b"{����\��Hջ��M-g��K�$�X)�w�C��ɢ�E7���/qj�CĖ ?�3��"}�A�b�_$�{>w^��/�~�	6,��RurD�G�aSC�ω�]:�r:G�qbӿ��"��f�^��5��BEw"c��e��p�`���I�	⨨�%��!���ɪ쵍G�j�4�`�LS�zFu�!��Ӵ4��N��1�i��d�	/��B�[�Q�q8t#YV9���	[V��_�Բ��p��:D�)n�h�Hc��j�f� �!s��;��Lό+�
؛�'��`�����k��W�� k�_ �5в�'x9Uz��_`!��ׄ�Rb+�gU�'�0���x
�Ղh�	�3'�8G��yo�o��T�F�7T	6�ֶ�%�1�<9�o���F�9цv�#���ad�8^1?{�Ȃ�����/K�]�Dӈ��%�C��:�d�y���X�� ?&�*�Izz�!����CF���3\vK�x�x'd%�S͈��t��ʗ�a*�O��<?��Rl�y�z/Ҕ�ҹ�_�E��B�¯��L��-\bC9�l�%�X1s��}9��� `2��qмTNo�*Sj��BHJ�`)�I�#HΪ:�9��Y����K*t&�X;�ʊ� �{�i���jptQX�CM�h�\?Y��j��8'�m��-}!����F�Qx��MR�?o��;0ت,�k6��JxZh� �Y�C/�Y����27ޛ�׹���T�fa�'i��ւl�Y1CIlƷ�5�`Ȓ�rR��:�եE,>�~��k,wɺ9�� ��me73"��;g,"%���ȵ�F���φax�A�]ä�LoD�%��*�5�J�qf���c*=�����8N)~ц}�%�}ʰ��y޵4ꁘ�R���y�^�s���мƪ'N8���C������)ׂ�T�2Mk䴰����G�٦�߯O�|����h��W�p�+F�+z�D���0qT�b"�W�qӎ���芝Z��*��y��� sz*��	����F{����ĔO�U� ����-��W�궪�
B�]�0����}�9N���@���]��H\���P���],䚆�C��x��o^�ڂ�%�:�M5	0�|��ķ��:�s/0���ū�?�X/��z�R��Y �����$r:�ʯ����M��d������w�R|�J����L�H1p����� �;K)����-pfT��aמy��e�Q��fWF�`�WPH��J�J�
dl_�?$о<4��ȑH^*����:h�$<ٔ����J�T�=��K�P:\���7=>)|>�y��eE�����������߂@�H��e
�{8�{h�b�Y`D#����q2)Cs[�V�P��8�`d�N�~Gt]�@����Z�+i�:� �G7����510s�wJ4 k$�ḧ́�p�Zں�(�Ԍr,.t��$&�³Kl	��Ĥ�{��('�2 ��?� n?�RHqwxY��C��T��k
C��ҟ_/x8&x�?���)��-����z<J%J�� ��
ʠpe���4��f[ſTUY_om|_�*�V�v�c�tQ�5�Q�FA���I��Si�Ԁo)�X���"�B̀53�Ү��n�Z鸍������x��K�g�~9�� 5M����z���DB~5��������S��E/�/`�R�F��I�53I�h���]��5�lFdaɠ���.����C{U��Q�o�������1es/u.!+������w��ɲ��3B2�3c�z��i�G��i�0:$�$��]�8�쪽]8	X��.��!�{S�_@�0��[ta�	|��t���2�9F��
[/ͻ�[�"D�� �ma	$
�M�8�HT�ʠ��Es���-NpSA�����JWf�F�8H4�@�'�!#���f�y]�t9�=k���9m�.^Ⱦ@� ���q����1߉V��5��\~�K���g頢�5��KIbNY�R0{i��	$yH!9�*��fw�����ԃ�+��%�e�:�,�V1���e|0ug��T9�đ��C� ��]��Iw�!�� ���c���zv��	���j���׵)':�c�ʚ�Q�(���F]��x܌Z��3F������k���Uo ����gc8"1\�~F��R�e>F��@7�l�_c�6,5���D{%��J�(Þ�u��*��%x��2>o5�W]ޖ�;f�ܩ��j�����)��=�=�W
s,8%Ӿ����ޔ�3�l����k8�F2}��K�ӟ��O���P���L������T�x/W��:��7��Xz]U-������(m��Q��`�	��v��SU�,�D�O݂^U��j���<ܓjE�iܬ(N1��2�������!�W#�D0���)��-��'ۯ>�oZ0��>�u��b1��#���t2W�����B&l�Yƫ׽{�_p�>8��X�kQ�T�ǿ��|���
)�?�������Pg�j��ț�]��0m{T�,�u��6z��·�3��~�Z4��c� 1U؜ �
rtn~�~�2����R�¢A8H]6g"���HdR1��w�&=��k# �?��m�L���K�s�o������MJǻ6�O�j"�̣̠m*�k���t�umV�Ty��o�S�"#��o*|�M�rS+pz*Xi困)D��'[�w���=��a���P-F�!�S��)��x��^
x7�ƦȌ�mW�_T���.u�mo�s-�y��<�h%�v������e�ܑ��x��'i�]��E��r�&�[6s2[��
lH�p/$Y���-�����3�\�;���@��@-:�՟p�/�>��?|>�:y�E3-�ޛ�b�5�٨��[��}϶[՝[��Y� �
1@�2�J�4����fM�?h���=	`��KjMM xo�d&��~�
ª7�����/�U�}���_��n)�V���x�\zf}ߒ�TaxX��b�y��c\ �]�ۀ{�v���E�F]�	|�F�����E���k���~��}�/㤫�ͱ�ߴ�E$tzH�6�4��\�=\�M�n�w�ۥ����_�i��J��bb'H�F�e`�_K�t��S�X��#$�>���X]��k��/������ƣ~�"��U���8����Q�n���;�y�uu���}�����*#�kSmV���W�*�dW��Ӓ����s�H\���d��)�r$�/k� �h�������Z�[|ߨڳ�r���T��HaBʞ����R�^@�56_�S�c@��Jo���IcK��KUPrY�A�#H�G57s#ű韠9�>�n���J5�%D[��/�/E}�����5Z���6��U��K�ρ����������%�:(U��s��A�Նl�zk
> �e{�GL���4������S����#wB=@0iT�F���馕a�����5|N�cSF��~.� �G�j��cA������l��j��H
ƵkF����"����h��+V!��;V��`���n�@��a'f��H�{�
'�8�T�ӕ��Z��c��Z/4.#&�I��\Ph���ڲ�6	;��R	��	�6�����u�std�m~�l�!ǩ���7FM��bp�_OgjԱ��o�wè|kӮ_�Z�KtJA�&T00)�&����B:qz��lȢ�9ڲ������%i�R�X7}�yU�g�f��.��	jN�@Ӯ?(v�P�����U''�1\jN�:�3\��~�hf�n_6s	������Wgl�x7C6�Q>qCB��8t��?g�)����SŽ� @=�U��G�Re�p�a,�n��k����`����|�4v�����!��b�Lm�W���lۋ�:f�=�Y��h ��;�f��f�����u�qM~��x.ԝ�#h Z �{u���+ܞ-ݴ����Hi��¹}u�}A�`��"�`0M�����w>�p ��K'��-+韒��Q����Jq���GZ]z"O���y��Q���3w��	��9l��]dX	����xQ����H�xq�5�r?%w.����߮�"{���9L�$,��z8�7I�,��R�Զ�}}��Tj)��zFg'Z&y8�H�ca�y���-�ϱ������X��Q]Y�oˠR�O��М��ɯ�޿s�2�u#�qd�I�M%�C!������0|{��O��Pl��F16�e�R���b�*���/��g�s���x�T���p�7Ӂ���Gq�RS�@FW�Z D���C����=�h��L�s��f��c�f��˻��W:EWi�dkܚ��˲y��X����tlW�R��yȽa�@G�t��F���ѧ��|�����'���V�
�D����fY�]�wT:u�BS`A���~('(�q�ލ��^5e��tB�si�܁[;����y�f��W�F�ʤs�1�H�;��`zh�ɜJ�M�!�?�j/��LZ]�%nQ�4�o^n#�_�K*}5��\t��g�y0����!%;0��#/c��6��:�Hs��b�5�%�	}�o ��ö���y�� 刞�/��3�W�1��@�-9G�Lt����C�[e"�L�Y�Cթ�P3�H�� ]�u�H3mU�t=��ǒ�?/Ѥ]Nx""���̆��>�
_^�Alf9��Zܢ�	���Fw�@�Z�G�m�H�@�X߾�q��Ņ�\Dw	;�,W��3{��Q�^��H:,˰�]��nm^����&f�?Lk�w�M �~��<��(����|�0ް|!���?vO��wwLZ��V=F&����1҃��h}=d�܌��7Y}�]=ɉ��K�HJW����/B���=j��B� {�Y6���V.�1��dZ��NB[p��mH����*����������P'�F$۰�)hֳM�P���`��5Rq��Y���L�s������hm���5&����ٸ2vq�B���1��c��Dʐw���~)3��ą�U)�7
O�O &+δ��!x����jX2�f<(U	}�
������� �����W"|#\���;Z�ʛ��d��fP?���Ը���2���@F��F�!% p�MO��*,;�Et��neu�L�e��gJ}{�ݸ�h��V��&��~v��ߏ�$�7��B�o��˺D94ء�2���7��է86��j4 _�I�i}MC$�"ᨿ��&+�)��H�F&�e����>�.�:�#�F4�"o6�P����F�ى�V�`aw���r�ΣF������R�8�zF; a���� hC��l�D-���o�8P;����^�c=Q�P�t)XAn�	���j��I����$J���7�dY��E\�|}�u�J��Y���x����B
��/�,s��&���<M�x�3bA�(s���dZ"�l�gZ��+��Wiz	W�%)&Y��ꎿ��d���FJ�g5X.>�%��w"Ԟ��P�/��|����[��@PN�E��ucT69�4<����̑��/,���Z�`r�����a �w�}�*���K��h_�9f�m��+�d�Y��0�c���q?͒��?�^� m�3��z��JAD<������܌�'P�:�a%:/;��'�
+�}Y�ZSdm������cv��:��o�_L�g���]��o��@���[���b����7���H�9h��9�z�#ۖ�F_�/�G�ƋF��OK�_^�,Si�(�YM���"��ކ��~����i�jٗ$��;�䠓[A�^8^��7ރ���]}�
h{����t�� ME�͛�O ����y?�w�s��/
��;���^&B7G�sg��)=�TH�m8(�:���ͤݼ����v�i��bj�z�BJ����=� R��e�R���Ȟ���AZ��{�Q��͇�&k��q5!�-q�P�D_(�F��od�F��q���^�iحSA�ۯ���謅G՚#r����t�+�������t'�������ZQ���Ē8	Nj�k-_�qx�V����\8����W��'K�e$,H�i���F���U+N��hm�����װN'���[�'>q s���ͤq�Y�߅��ţ��r��2O�kq% �r,���t�2,��v�W�"h1|�<�d�u�_�qX���g2X	�|K̄:W�Y���� �u���=eN�)53�g�1*��V�z5^���(��_noз��4��~���j����P�����"�1Dk~@���i�2&�/�A�����lVZ�n�%?�D�W������^��0̱Т��[�-v�z��أ�R4��KuX�p��9ݠ��bv����br�z"5�}ڒ�T2��mƵ(zߢ��dxlmRs��1�	�=݈T����M�M�_�����IW�HT�}�KH� �CLo��� �+�(6��dq��?�tų?Q�aY���
�?k샜�� U��B�M�[hP,�N���LG��rCgo���8�ة:Ė�9�_.������=g#�Kh"���+�w
��?Z�~�����/u_�u����aJsˈ ���r�2�u�|����h�1�붴�$��`p�&# _8@����:Dy�9V��@�� &)����o!8��#��fn-�ۈ�s�e~�	�IQ�G-LQ|7~�¾��9�+h�4�Gp��os��� :p�e�����P8��C��
�7�G��p��CF+���t��T�^5i��.�,�*KZ�1��כMtg}I�g���a�j(#��$+T��g:�^V��	��]������S�<˱����`2�^����\��YƔ�u����:Β�_�5D๖J�wT�6K����������V{G/O�/�B�ك_��.����v��6pi+Q���`$D3`�#/��WW�L<�J>ÍWG}�?lb�[�z�漓�h��Ϫ�A;�b��|��2xr��|o�E�Cy�SG/���cS�X�㢳�򽐛@;(h��fI�cw�V�vL��;����i��>��$���6�*q��E�C3"- 7��-=�h��i�*���tJi�����^��v�e	2�(^��B����P8�R�=��iZW�q��5���j�l���G�2�!/i�;D��䴫�ƐD6@�J�q�}2y�R�_�Xz2���j�@�
�o 2����䖰��w��S�P�}xx���^���w3B��G\ҋ�����y,���6���O	��VK_qҥ)(����s�E!��)�X�l	a������f,��*"ϻR�z��qhԱK>��J典3j9?�E��#�-�Ro�|O ��9 R0�V���C>�}a�t�;�.{̳1p�����j�mu���[��hLwLXq�����2?a��'8'ԓaKc��0\����*�pV�E�`���T��C����?�AuZ��ra*J-��5h�^
N��kؼ�N�ip�^ԇ�������co�ۤb�Ke�@&�_��0�d�ׅ0@�D����#����yo��Н���.h�ڜm�����w�_�G�/����-���|�[�d"����d(����W1ܾi#�J�xc�(�Gh�v.�2�)�P��E�P�uJ]<T�Q�QE���Y����y�޳�(NO��i��	!�|���M�n^o~�55lr�}=��[�/��߮	�R#���	]�����׸�,*��OX������O��REs���և�?�t>	�LR>j&�y��+���e������ӕ�y7��&qme��6$و�r07�X���H�L��ma�*	p~��1����yj���.Z,���җ������H�*N鐥�܀~s�.b��H�wѝ����P�`9N(Af���נ��+���
.+�~0G휅�0G;a�e�T��Lߑ.οfa�N����+7�m9�Ԙq�2��%�	l��-)�ak3Be!�"6 ۷9�R��@����]��8h���Q#^�E#��h��O�ɥ�D��q8�wX�%Hn� w��×�?s}?�~�ǚcX�������������X�ם�+b���� '�zd� �b,���j��2���Z������l���U&�;y��C�;�G�u���� ��|�X̼J�� {���ݙ���:�n�����1����~6&/��%��c��Q��ST��Fo��#Z_0 3�F��N���0���6	d�ʶ�r�NHAW��sa���A��Wl��T8U3	�}�7
����<�k�-��� ��\��	�����<r��a[���<��"�H�Mٙ��ԍ��0�P���6�9K7Zڔ$��S�,A ���s�}k�,X�]k{�+� ����n��8C7
�S�F�<���=�37Sr�8�Ý�sRc:��/Fأ;�$���!h��d�y�t�I�:V���H�����}�[�'�VјB.�w��储��w�S��2Vu���.K�W\	|��V��"�E\
a��h�f7�����ף���"��(�h���Qc��MF}��3k̐�le����BNx�iE�4�E��Bev����މ����N�A��ǿ8���_E����3\�4��>��w�d�����UYɅ&�)��):@|�e؆Z������K�D'�:��T���dѧǁY��e��t�����OѬsF�G�Fӎ���5Hx�_/_=�(��Է���K��D���L������:����߱���fty�ue�l��XbY����֞�C��\t�
{�S��~�_��4�Ж2c+sG�U�:V����=����TY\��+E�W��d��pR}�8/�O�'���W��E�v�+�éP=?^����E��o�э�l�Hy7��޹���x�A�0e� �z��U*W<Va��,���fwY	x%��~����mĘ��$���FХ�ՀRmp!zQAv&��Wws���l��z����l�h�n>���y��6z}/|�v�/��er��Q0�@=�Jk�q�p0��?DpM��]�4��pǰ�.�j��"EwO���'��
T:$X�˩N�,�=� ��ȷH gʛ��������zw���@�w0=I�l}�i+�A7��#]�Sf�Sk�),qr�=�Gj�oBw�<R̦@R���I��k���k���F��>����ңn�����}����^�Z[U��*j��_F���v�*�T�Qy�ؔ�8l�9�D�l�b����Y�X�ST�#��~�N��=���7A���,��AI G���O��)���Ư1����Tû�C�i�ٴ�H�ò�[�o�9�*%eQ�5�d]rAlՊs��Z�^'���#���GQ7\��1o8Y���>a��s&���r5�_�y��5�ڐ��������)w�'ۃ����=!#V�;�a���e {g�I�4-l��{Åȷ˛tm���>��M�Ȇ�_iK�E�:���hSd��w��q��JN�6���<�y��U�I� �g����E���}[��=5\�J�t�J�B�K��
Łd/o�WeX�d�� ���A!��[m��T�H����n�� M�E��T�*��٦�����aƨ�&��E¨���/7[S���a��?)x�Oc�a���Z��):-\�>���u�
D�H�������++n��>��ċ�#ʇE�'i�պ�/L*dUݺL��f������oA�Ⱥ�@�7���hS��n��>j):E��
:��T�M�"�_·����˒��%&GT�~=�zf^
S_��W�������Α��5~��<�[z<�f'>f�������h��V>��Z�9��N�]bT{ז����}UiI�MRɘEF.BR��hPu/^�7�m�?%V:�Hڲїf$4��M��pT��*���
���e؅��k�,��(_���Υ�y���gv_�V�n������%�,�r6��,��~��K����~�}�B{�|���;X/3L���AYû8xAr�F�-��f�v����0Lmn:+Q����� �\��>J�d+����j���V�� 5okŢVRHk���V����Z��[Y�k�T)&�`������)R�cE��^��H�!`[�
���!����1��:S["��xlݷ4��'�a��-]P@X�n����MQm�{��kSE=��p������}�#�B���k
I~1���DG�ƪ�G�x�V[��M]��嗍R�M'�-���t�g8�DT��6N|����Yא�\�f�GTI�.����@^9AA����虇4�'+Ͼg��O��]�\����UB��A��W�\�����U�~V,`Д�F	����d����+�s��D(Ӷ�S��b1��2uG3������k�l��G�-�7��B\���h��`�!�����W���N�
.J�M��,$�^v������J��S����aQ_��3;�����ۧ4g�v�N"����H��=�)���P�p��Y1j���]�Uۡ���Mq�a���=�8f��@�=���vc��h��W	<_y5u׏��Т�F&S�~�W?<��`P18�bxIl����xU@��W�E������(�]�I�.��cP��B2O՛6�����(��*>�J�e��w����G0�?�D)p�BT	'6�1'������2���b����ڡѲ;�.��߀\��	eV��t�F l�Ip��j|
r��R�G��|�[��r�>�$�1�8��g����Տj��Z��1	u����ӳ]��o�*�t�mY�h�)�gǊ��U���9Y,{꪿��#����k�(*6#�hD��"���4/}1�Na��E�c`���J
A�u�>��`(��S�u'עq �Ngc����Ҟ���z##�� �V������\�SQ"��n�$��,
�oP����<I�%�E�Az��Y�x�ד��)�7�#�w�k��&����zG;���h$�S�n��T���.�-��(�q�I�h=~{�-%*�|k[��4oc6��S
����9J���|��&R '��rM�;�b��P�4�,�~���6���G<�DJ�Bn�E����s������� �P��m�L���Nx�R���y���CR�z|$X���QKF�K����1�I��
��,筿�}%gx���*]�������Bke'��w�F���4�mm��XbO�6aO�5�f;��nRG�ܼ��z&���8��GKՐ�eg����(�C�w�2�E>��|CC��_�V����ΖK_��]��GE�n\������tg�LR;9�Y@3�I����5Q	Hݱ�3���_����d�ϴ�]2 B���*N'۠Q�<��;���u�}n�	�w��x��� m��.x*���)�����_�"�u_&9��
���x�i�aS�r���-:&��uv*��%FB=� ��*+�J	@���y�=l��.N�N���0V2�Yı��9 ��½>��"��;T��'�s��dyE�@d@�<5�K-!�l}>h���� HY{L�u�n�	ݠK/c́���Թ�,R+����(� <��D��?����ΪxS#�0�����iH,l�厂#¨Ť��:����?�V%o��딎���?a�C���6g�����0l�����THWn�)�M��Z���K~�s�³�|/�������@��F�H��&���}J�cXy4xnb�@Ъ|���Pbǋ�]&ŻXt�oM�W�C�4�7���~��5
�׿�`6ƍ6H:5�B!�'<<6�/��=�Hq�1�+�Ӣ���.�*�v�G_�ER]=ns���~�� &����TE:�&�G�&e���6"�&�ԕ+���
�ꎄĸ���}�i��{��mK������I���rKX�7����� y��?KO���c�9����[L2��c���g����&�ܐ�8�Κ~�`�Kj�شuBg��/ �>D�s[�;Βj��]���t띙o{ן#'�H�k�βr%�$�^�E��������b��*�N�t�rt��~]���o)�~�������x�>�;�{H� �o϶���6�g��
5��IQU���}i�Ȩ8�;�ʭ�b�O{A�Q�_E��_���Nre�h~b+�"HN+~B�r����W� ����#f# e{g���zI�����C��t��2t
N�F�eu|O���G��~�S<��Ŗ"5Д���� �G�L�Ȃ��YR�v4љ)^��kxH���Ά]B�j=�;�:ԑSa}�R���y�'�vt���f�Xe��:��M�z��>* �#���T!��
� ��)q^��m;a�������}�?�l�q斓j����(*�̎�*z_{��c��zhߣ�$}��Z�K��B���I'D���},+WvEb#�o��!"�������i8`�c..l��2����q�ѱ���Բ�t��,'a���1�쿱�+Н���zI�	
0���&.C0ww���FxLf3���}�`���IJ�O�R�=^�P��>zG��WW�|
|�����n�ٹ�G����!��T�c������4��qG��D�HX���mhxq������Tۊۜ[	4��V��*>IUX�� �H�R�'V���w�QIwH��.�4*��Æ6L �����������CORW[���5p^3Ey�h8;��ghkPr��b�걁=�aO�8$1+1�-��8���-_q(c�=��$[���K��9��iv\�׸��CDF!�H�v�qI��_9�xոV��UB��s�r_�M��
�AOB��C{��)dm>�+>�N���#4�
�\6��$s :�k���7�t>�wq�o*�'�H�j�&j$��Vk��r�r`v�3�9�q���oYe�.W'�\�X�h��ˢk�]0���/K~bjA98tب��P#Z����S'����{�#�,Y"�s�S�X�O^��{W��
��V�s�hpm���2�;�\��}��	d�r��Ɨ;��)}/M|8F1�9�8����{���y�8�%N����*��@W=��<Z�ϓ��6�5%�d���t�΃^�{����Jb{�Cr$�h�����`��RĲa�\�P�$����R�xG�^Uf���m>��;��J�><���֩���9T�L�҄�V7�ּݫ�_y\$ɹ�$�#!����)rsD�cn�:1��^���~��߃��K�0���V�pH�ij��,�.��zy��'N=l�����o"	~最�G�S/�8��s�l�3�3j�w��uO��q�>7U?@!p%?�Yp״Ut�˽?W�8��%=���8ި�s�a:<�N��f��+y�WG�B��K?�A�u�}��^pA���\ ��3bP���XF��o%��c���k蠊x�Ur��$�y�i68`���d��m��,�Dz}����k�KQ`�x�h"]]�4��s2�8Fx�tUtV��zw�U9|1�-xT�'�|vh}?�̙�d�fŷ�d���S+�
Q��0���>��e��?��3�+��	�ь&���J��>���	����'����އ3a�G�����4i)�ET�����]uV����؃`�}��y�{�O��{�.i�M��
��NU�Ϩ��TJ������{tw��!u�,y�)0�އ�[`��=0��ߦz?�"/�c�8s<��B��bL��Q�����/gMxv#x����������bn�'�Uz��>4��w�M���5j����G�^|u��eO�\�v���V�*޶YT�u�7�{F�KB��������q�IQ����C!����i*���"�{�t[�K�Pz���B%-�rH���AY9Қ�LdĂ4���!�]��>?���F�{��u�}�s�R�Ft�A��WV�^��D���O��R�i�@���u���g�[B��������Q�MX���!%ﯼ��Y�~�7 ��C}� {�a�c���
.z�zP�Z���
����l�y&���'�V�O��^R�K�$����v����j&�&�ִ]���oBdN����с�r��8� IB���m��I�?>��?��"9�����h����N�$�e2i��14tc��)b6��K->�|������1+�M,��n�*�}H�l����4��b��ޯG���N�{S{�S��%m��aH��˧8G>+-
Gde��V�	Z�K����u�Z��@�r�ٗ���[�8TܪV#�pG�|6[�"�ނ�7�J�h�vF�.)wBzX�� a'.�jTd���#K�aN=2�ʜ�clB�����3To��uр^�޲N*t��ɼ1���dP�R���rI�o�Nw�淞6��Ur�%8�I��4�l�U�E];�@i���(O�IJ�ܬ��X�������*��xpߧp�����8�ƺF���D �#*���==!�Ӆl�ǿ��{ʴ��k6ή�o���x�#�B�;D.�N�K~�����լ-G�Ў�N|��H�lJw�ll	s�]K�%�}��#��e[��K ��,..$̹�3<(m)�<i��v��� $�m���6gb�O6O�$��f M� �1åy湝�35(�1
Q�أ�Y�ͼ�Ȩ�o��v~>���(mr��(�MFy��,I_f���Gcޮ�<e���%����Rg�HYx)�,wq�O�"�:c�g����4��`�E|d+|�@���S������_ɥxB�xN���l�B�Y?��"C�(���7Y�C�n;'k��Cp?��v��<�enG|�X��ۛYbHY>�}�s��\��F$�Z̩��3i{~8g[�D���Gy{:%�vt�����碎u�]�sO�K�+�dRKkɃC�0�T���&7��(s�CA���������S�v������'�A[�>����K=ӾQW�?������G=�L�K)fqtz,�da˩�����
�f=��)���;�DW��H�va5�֩�]�$��gA5�0<||YjJ%a�2���V��:]�5=�\`1oV����~>��yַ6U��{��G4�H���+�R�h8ΐ�6�+&���㠘c�f�+G:~UȐ>[��Ͳ�`�q`pS�K������S�~ލQ�iCt�#!Po�Jzq��w������EJ��t�fȯ|���M9�\�O��y���Z��`���г�ْa���7Ͳ��ֆ�����0Q����\R�Yv�r�G�a]+���ΓTߟ�c:ia�w3'�csܹٳ��/�WOoKZ� M1�[5�gd�:�L���� $��!2kKz� [jr���^��,�F�f�h��L�Ơ]�ײ}�#�E�3&Nss������$X ,xfz��|�W�w'�l��ˎE�P"Oh0il5�]�:�p��`o�P\ޞ�������%�z�b���V�81¹��h�!���eȜ�B�ݣ�o#��d�\|���%�y�<��6�I���d�cQ��/�*���Mޜ&6/_p�r��+D���ܡ��:���?W��g��I}%ۏ��G�GCs@��vX!˥��7^�UWK���fM)cT�QV�x�q��;��f�v)S����k�ub ؃[Ca�!c�<@�09�� ўe�g,o���)��1*H�;~C��B�����퇊�2�Y�*e���K���げ���ʳ�ܩ�J.vL�$`�u{���m<ݐ]s�A5]E��y�㎉P���ɀ����A�y�z��c!���zJ1�s��o8El\��J,3�W��. x�jFsFЫ�����Lȕ�je���d���=p�X=��=�jb�ȅ/��0`_	�f��p<�/�Uv	��+�@�Ն������q���"Uq���x������>�$8��U��]���pT�\R�VK��WX�X���/���g��f"?�m�LqU}�0�E���u�E�&p�;����c���3j��ۡ��ذN���^�y�DyE�� #4s���g0�lK�L�i��u�})��~���E��L��]b+�n���ם6�1��}8H���,�'kx��x���� �'��F��e_C�I(Qh�B�%�q]��ȅcAWR��͹Ҿ똨���o����*�H4U�sZ�����%(�B*/
)$���)܃W��A���k�� �9�4?��FW�����\U��G/�&0 �B�Vy%2�Р?�(��3��s۷�^���F)ڋ�����yeRGoٹ������ң>F
2���E;�j��	%�ںcJ&��S��~ ���xQƋ��ju2�����S�EGs�׷�6�,�%��h�Z��mW�o}-e���7��D�g�ﱝ�W��B#-�_���|�@���Q7���c���̣�_h^	1�E��ƞ�4�K��_�Q���[g�����Ő����a��vݡ�:�+=�lk�7�=���"�;��O��l�/W�m߇��M�Ğ w�+�'L��.O��qM����S���_�{d�M�F%�����B���<�̘ )���;��v������P؅'�M���q<9=�_��� yN�;���Z�	n�ŷjs�Zb�C��${�E�ô���-sL��W �/�ԩ&�YD��:�Y#xۚ}P���w���R1⇳�X�I�>[�w]��~��D��8���K��ÐdQ-��ͬ�B���u����~�EV>���-]����v�|p9��kW`����!A��
�,P$6���ֆ=)�2�~���8i�0d*��А���C��g�_��j���Z��O��J�(�qn���>����
3��hlA�ZX�2������ң�i�2b�%�#����t�2W���p�?��D���!�����m�k:�7d�F�lt�ǩ <�䛲P�F,?�LĒ����y�r��R��ʗ[��$� Y3����)�?����a;���uDA�<��^[1�ŏ��o�J��"fm���R���MP�|�!6#�����!~Q ���޹B� �h���¨ت����x�8�D>�W��>!w�8���z����52A�� ���CYyT�][Nq���"�ՠ�m��Ҙ��Y�O����Ͼ�*L=���|����t�[���;��Y�8<�bރr�LҒyJ�R?S���'����)��<̐��7��Y�{9%�|K.��.gΨ�c���Gr؀��a��I���_�Q)��9�p���EgPsa,� ��F$>�(�'�mJ$P�S f�� �ȳd"�qS���_�T�C^8�m�~�(�r���������'��}��=��)+���^"�fEE$Vi_����uc\	�v��%y��N���¼8r��ǚ�-B<��y�@�#�1��(�K��f���ω/��M?(��Xl�&[p���A��c;���@zPOe�$ux�"� f+��x��/���U��7�jh�Agq�ˋ^�����;����c�m�oC74E����z�rV�%�{��1����%�q4�G� ��ew�Cw�o�yd���x�B�����V�$��&%JrF�A+�����.��?1fæ	p���6�}Fv�� ���	@�[ PyS6@� ��r�쬝v����h���!.�=���~�8f�	D�,����g}�X.I�«Z��%Nc��'!G��E߅��ޤ+��!E��u%�	����G��;
Η΍�p�3X/�f��E��q	�Ɠ�S;Ts�2��KL�!Q�B#�lYc%����mO�Q���p߉�2��Ң |�XP2<X���>"|L������A�F+IJ�  ô*��be$�F��v�Z6���\��Rz(��k��zs�A�^����
Y`�[[���� �����<4*->3a���n�@��Wm��<��Pن�qs��@Dȋa��$[<}Mj0BI-��`�E����Y��dߡ>��5s�?H_
)<;�)|�1I��&pS�C���z����Z��i�U�2����?BQ��j����-	&�ԫ\)I��ʼp���8-�;����j�yB
�}G��e�wT^�|���f���ʏvLE�tԲ��WRC���-�88�H���:���d I����?�^�3$b��	�)���>L87-�M�ާ�9М`q|&�V�D�ؔj��P�JT�־Q&W4���b��������&k���Z��k*m3?��E���7�MR����|}N�a3dF/��C4g����|�-d�og��b����e��5�)��m[]��5U}��U�����+G���9D(�-���0���G4�ID��;zi�wZx�f��$�ېd��8׶��-�M7.C?� �f�raAG#���nVR�2�����"	���ag�������m�@K�(MDö�`����m��5���I�U-6�P}����3(�'���
�fq�ָr1 �o�j.��=������]IZ���6��|A����S˄���b�?�(�.Q+.�'�����h���Or~��m܋A
:m��&���-;|���[q�]�a���Q���Hzcn������X��ܒ ��o} �N�f�t����G��*��5Ë����d��q�s��%���N�Ű?y��%zA��4�z6��$�[V�?У�^�vIT8�uW�H����������x��ܮ���X�2�e7V�,��Vp�r#b�3��"��:� ^�j��T�S��v��5�������v�s������p�X��ư����X�1��:-~H���>B�AO/��z��N�A6���'��ûa��j�<�n��Y��y��0�9,	�����	�9.n8�QM5=3��$����G��Ǎ%V� �SKo��/ǵ  /�ˣ��U5v�&�(�!i��Z4�H�mJ��Ϙ]FX!�� lN t�8���/�}��#ʣ���"�`�i-�-�>�#�*R:��1!�M��ɛf��cpbI"*�����2�ֶyP�_D��%FN�h��.�i�D"��7���#?���}%��`�a�+�r��/���W�;S��Mo��1q3�eX�GB-�w��?��<�x]?	Jol��7q�m�qZ)ʊk��@U�r�i��$%�y���¢t9���H-ZW�K�*�Ql��WS�؍	-���׬�Gt�����6p�aK�bw҈��Y>���"��(�����|g����y����<�H��0����%c4�X��>F�/-k��j&*^�E֟��.S	zd0H�{�۝������B1�����N߭� ��O������8��5�����7B���Q�ɢ�;��,=��U�I��Z�!('��Zb!�v�0a/��"@����DJ��8Tk�OY�Wi�ݗ���|�CB:CkS�^5�!�֋�Qu��U��=��m
�2��S�iѼkʯ�R20��,�F�ט抚=*. �ٓn-���Uv��hJ�N �Ӳu����W�f3��{�������A��'*�BZ
�'3'^���x恽�P\%9�����nǌ�i
�Q��^Uѽ)�锹��o�j�������R9؆gl[���	���xA\�ek��3;�g��h@��uV��vbl^n�k^��4���pP�:�v",���c�)�. '2��]_��Ѹ�%�G�[��6�!7�XP�6_`�l�V��p���Zr�N}iN!�'N7� $Y`�3Ak��J��N}#u��B<p��cn	M��5nM����h���b��.��4��P��[{r��5�P����A��U�  &U�E��K�iwmx��I����C$SK�+���]�F��O����X<�
�g��&^��
�*dJ�d������=��ʋ:�����c��	�� �3��܉��Hb*D� Ӆ�mf���*�;�5 �$��/-l�~����q^������V��?�䋮��\|�CIg�����H<��,8������l��De���N��i�F���sH��	���@����'�QD�9H�n?�K�X�N;�4a�vo��j���R�(�k��O��L�pDq����x�@����rɥ�� ��n}v���	���S�"��3�ަ���PMK��ƈIE�S8텮������sΌ��uU4N��3���e;N����$t���2@����B < ���\�3@�P�q<B�e0*�sz�TA�?��cYn�,c� �����p�{H��:Q��6hs�K��m>F��h"���{��@9o�u�%��v�/_�W���� �9̜������lq���|f�r�lNV��T��cu�X����K��F8 �7fiQXSN!��%�w��4�Z^���!����-�r-T�P^�T���V���S�lVN��x�1�O�zt�-����\�<<�]<Z/��XԪT��O���]8��unCu����%��Dˀw�!�o����"��j���YP_j�W�Uz?-�m-pij��,���T�uy�V�`��N��C�Q�����难rÙ��>ahG�n��=}�&�:�3�%�Șo��D�7��m"��ZR���-✷0�R���K�F����:�B��R��b�2�BPZC�Kh�j��~s�-D��B�?�䨓��R�1n#��o�{I�#6�O�n+�4�LhjD�b�U<�ջ��F�خ/FR$��V�/���u�ĵA q�È�ߑq ��'L��/R����
7����7W
�*>|��}��!��A��LxO�}-����CP���v1x @:� n!U]�XE`d)k}�x�l�W�g���@Nn�8�3�sKRy���!�'�o;����w#t�^W���Μ�Y&^9J��ȉJ<g>v�/����|NԎ��Ӻ����+�c�q��&kS�5�.�Il%<��\���#[�t�=$����O������<S� 0f#Kь�ATC&kUN�7�����#Q���c8?�ew�s���y���d�;�' h7v���	|��&K��Z� Mʁ���}����v��(