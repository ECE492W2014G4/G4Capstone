��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P��v�"<ߞ��&'��k%P碶�R�ӣ�sĞ������FY&ZQkƮq��=m?b�uм�8��ڡ���Z!G�l;E�R�aJ��4L"Ǭ�ù�fG�+�M�9m��(%$SX��n��q�2z@��4j�'NM1�b���A��NA*����B��y�`,���Tv#�~:����m��e���f}LE����Fr��D��*)/"��v�EwZZZ�PV���Фq�5�	����^�d|�:�"�{IQyp�����K0�7��ظ����Q�ի�SV�Ԥj�c�2�Ƙ�(
�^��]CPa����KCH�Z\��u�R����0T~z�-�Pzd��_T�َA�� 3ҡ0���r��<zd�W1��bf��w�L��o���E��:�* �T�%��;Yy�N����N���A��{(K�q&�D��X
[��k���ռ�oEQ���6R��8����	�Ot���l�<���L�,�H`�x�a���SZ��,���<��l�/��l��^�\�l��#�k��_�L�����[7�J0����؂p��)iG ĥC��)����T諒�"c���b�,�Đ�7j���������� >y̶��R�ȶ0jυ�OG=}í�7ǯ�PMQ�(��wx�5�Z���([_��Qn��1�ewm�1�Gs��V���L b�A�H�@���j�w�ݮ���������X4���d�E_.���낼���-C�F+���i�x�!s�K��3�3�A��g���Dc;�}h*û']G��T&p�*�V��A牍%(a���Z��p������.c͊q-�p�=A� ���x��;�V�D֑k�5d�磄��y^�༝W��U~O��r"�"���n���r�v��Z��C{��|�>�Ss��T.t��j����A��F.�_�mw5���\���JC�u����)#���� %���yjъ��,��^wK؅B4�YI���p�Ы�]@��\C��s3 ��m/xGk�/y��}�?x�����_z8V�W�G��9P�Q\^2�Ğ��kxp(��-^��\̶��&��!��Q��U u�"�?ڇ��Ut(��<�?�h�'�8[�?&_�ʓ��v8�.@~�V�c�Js���9k��{�c��i�l�l"��q�t:|�ƭkN�sL�%��6Of�+����F(%Rr��
#%�@�#������[�n=S�t?<)�p�0�Eᦴ��b3�K� P�ݹժ�ؐ�������� ��/���bOM9S���"�@ow~�U�_w�h�ک�7��"��P<���weâ�]��-E�k�ND?�oO�d]�x��4��`(�c����3�^|�&�7��C�!d2�W�.>u�.*E���6E�R���c��kP{N�d4��T�X�Yyj����fx�c/K���N���2.	x������9Q_Ѓ�4G}��	0:�4��۴&��)���	bW��7�Z�ȷ��I#K7�#c�ٽ[�:���B��}v|�M��eU��%����}=�A��r�b��'�	�T�zpz)��֦ICw�~�J���zc��^�ms}�70��w�{����q��d~.'+:-����. )��$��;�����;)������֘:;��L=-�ycGս��6��	B�V���Wƺ0
q1�����������*��3a����b�������9\��AȢ�[��)��l/��k9T�B[��5�3�����+��z�匋��3N���;;��o�*��b9#�L���*��izn�u�3@x�fD�`��
e����P���4�2Ɲ��Q,���&zܒ��6Tx`����nId���`��t�����.R��5��-Hf�-E�do�\���A���3�*�� �+�Q��0.����C�EPeP��`���^S^��������\�[�.�ڙ�p��8��+���Ƹ8D*	�NC����8�U�5g\&��Et�:Oe�e�����e��9g�A�B�/d[�gҒ��m�z�h����f���s�IQ2t}��{`c5"ɰ��֨V8~F�]b|�#QK�Ž�u*��L�gm���V2�d蟖��w�V�u6<�����W�a*Y?�;u�4�t����}RJ���>�����aL�d=�nMZ����D�E�i"�`�γLj�Xj��,kih��^�{�.�+����X0��I�o�"�]̩ˆ�K���D'�R��/�32Z��c�[� *��/8F���<*-���q,��瑴S�^{��7�_��G�C�Ѐ�/����� �<I��H��|�Z��dM5����=�9�tb�W�eZ]ke	�Y���� eE|��9��|M��+6��_��.�}b:�pd�Ȥ�L�����I���Bv�В�\
HZ`��g�S�~�NU]���*�g'E��%�Jni@���Q25i��wܥ�Z8��%F�n�G-gX6��<50.)JzT����4�0����Y�bD���ˀ�nZ"T�c�~#B�T�J��A�%F����#�o�B��_zO�nL
]��`��Z��K*��w�/��([�>\��:A���)8ۊ.�����z����Mw���+����'�D�|�>x�PD�(��&�P��H������@�PKy�E���Ɔ�6��͡���VM(v_:�nJ`���^��Ont�����Ƽ_6/�g�F��$*���v8ĄXwp���c�%�;��l+<$T<qw�3�w`BW����3?�B#n�o�Z��. ����Nm`�0�~���.��.-��;�'�'�WC|��		'O���t�"�gy;�G�f�H[b��������u�����G��.:4�/�L�wn����%�/,e��G����n�s�\�yp��\�����c͘H�9�K��6����";���#�_w]64V�����˕���O�����Ed���q³�������<ă;��Q6�U<'���F��e�!Q��Zϥj ~s���o:���H�ٶ�������pw�C����	t7X	(�;h󧮭��@_�2�c�j<��	Yj@�V�*�� ���TU���>x�m�0�q�{!)������o���;}T��)����q�63$�|�~�b��Ѻe`��7��2�{䒉�5m(��� 헏N�.�n2Ԅ�q*ғ-�x��Ry1ˣ%��ۇ�_)�(o�]�"y��d!_P��p)1}4-;iB�T	0r{�oy�q�n�:S��1
1�cK^�ޝ���zW�Z`Z�dg	�<ݩ�e�� A�gg+�gI�D\M��+'���^K_4������B�qv�A�����1�,���iNb˝�`��������ۉQ:�?�YV�T�{�4�QNQ,np-z�"Zg�gP��ڑ������^��0�S^��z ���k�M��6���z�
���O���.���y���gk�,%�� ��-� m�7o�W�E�.N��n��o���Mc=�#�1P�����x��4X.�|wk<��&�B�?8��%(���V�"��3�qͥ	%燝%IP/���>,\����ҋ�'
��Q��^�X�`W%�Q�4��t.7=�Ǳ|��cgoC8�<����V&��ޝx�4}���[Լ��~�[�N�:�ɢ����B�V�T7õ�J�$�'q5�>	��L�N�hEQ./
��Uz���8s{G���3YsF�R�w{��'e�+�#��������)$�E ����Pv|��,T��q
[\?���i�J���ۇ1�"7���O�\,�)��:*Zs�#������E���XD�)�]N��dE&_������T�h)�"���N��>x���8�g�3<���c &�}���O�͊dz�����t��� o<�S� +x��� a(����p�����cwp����%C_�k�0�~�˜���!ҊGj�ڠ�O�ī���$mb�^	f��Z��'=��yh
���� <Y�BKQ�uH���dAWD��`ia�Y�t	Ě�:!�(��RI�����2�u��t|u��3J�BG�������K��M$d���4(��/g��]{"�v%}qFhr z/Dt��k�&��zpl��h"�S%^ ���$JGAN&��TE9<}��}1قY-��X���@N�㿝mL<x����>X;�p�]ȵHσ�6ՑZ�><sRK^&��F�N��t��0f�2����XD�*L� ����B�T\�,�Z��.TK�w���?�j��0:�򒉦WdkBz��2b���N܏UN�lt\��>>ٷ�Pc��-�L�����\Bk t��r�g�ȓ�M�K ��\��8�gW�W���)�b�*uB�<�Z��߫��#$N��gK���TH�V��-�I*>�.�ۡ��A���K/�5eUY�ȫd���/'6����:�ܢ*�
��5�����6�;/^��������9ؖo���1�'csysA�7�<�=���tA�\p��O��J��Ro^næ�y�`�p%�T᳗��P�j��/���u2y���U�X�:
Ѹﵠ��a���g��D��}y�����Mu��J>P���6�� =�������ch��=��u橚]�n�Od�o05ŉ�!�EǨA������OF,�%�Wl��"X�Thx�TXv�>�>s�yB4VY>���a�2�0�2�U*�R��h�;���V�;��V�� 4�R��-�$�(ڳiX�0[ ���n��l7�_VcU�����a"�y�W �c���.����z�a�� Ir7<�K��,ls,y��������j`9��W����Ri�X�;����{<��mJ�XZ�?�}�ڸ��)n�P�)��7��A1��8�2�}�V&3��}P�P�{�v�N	)���zO��J<�`u���E	ډ����e����ڪ�b'xE�o�v*Gj���h��/8��R:K!3��V$'�?dz(�`���NY���3_m�i>���Wק�錪܉�[���H�}GR���h�!�]c��W�$A�7h�#OQg�$��Q7/5 ugt�S�}�\�>�8?� �'@iH�U����,���5�,V�+<����ь�������@Arr��/�@����(H�8/���zp1�O�dʼ�]5+�x�mtF����7G�v�X��o��4]@���^�9��n�r�[�]��ȏSI"�/������>r~]h�808�G����=��N�H���T�r�\�LèT��s���� �W稭�E�ZH����j�c��P0���/���_�N��S��yr�H���~s�w���5-��㍭q�Y��V�E��Te�?}jp�!�ۍK <8�w��2zѤǋno��!��L��"�vQof�gjM��T: b��8�<���B��N��z
������]��A3m���q�E?�O��&G`ۋ=ﶠ�xyZ�4�ND����NF�VVd��x`��2���jR�㇙�<�5��A֗��m���2�M�Z�y��ВP O�#�\ @�tL��{���I����2�[kLf�&�Wr��T�^y��?6�����s����}��LgѬ/��@� q� ����/C1��:�oi#�fyG>�ޕ�=Xܨ'p��u0;�0��;}����n�ѶX��Kz���!P�D��Qo?n��3[B�W��I��	\���Lz!2���N���u���
C�r��Ɂ3�u_��ɧ'���r�/�\4����xO7��������?3�|aZ[s����D�[ؠ���h�O�j~^��{C��w��MN���p��e�d�ɬq�y}dm���~f��zd�X�q��Is_���C����� }tg�B7+[�B�� #� ;C�%�Z��	�r��[����v2�(�A9=.����] W�ãH�Uoݹ�XT�o�:BiZ؟x~A"shr�+����q}�~�V�V�K�?Ȑ�m�C�l$l��Y �{VL��~�[Y<Y�K�v<:�Y�s+�Մ߄	�x��.�<�b���tx`CΩ�.�e�nB���Ԋ�䄡/Ȇ��-����p���A�{]���rv�VIj%�V�Ɠ��FKqL@�*-=9���_�ժO�T�i��������;$=$�(G9�"!<�ں�6i�h�V��.a���B= �Qi���j$ن���(�eA��A-ƙۙV9>
�
��q3+ضw,�e����<�`EK����2��k�
��!�շ)�shش��K#�{�#/���1�^p�����t�}�Y\u7�ୁ�	%�y2��k���Dl��uU��� ��1/��9���Y�WL�U��ջm[�'d�n[}��&H�it�o�o
����3?�@���w
�1E���>fu!6�*)y�֟݀qt������ZO���Я3��4�SU���9�
�&�j����*��;0�ma+z�{r��+��:j#�g�,K�*�)�OGfET���Ki������$�ރ�Hc���]���R�J=[	�����^�T4&���f�掍�ژ*�#k1�oH���EN������w�*���-w/�o��n"l��/��i��rU�������-���7�����e��EF�Le�`f�aQO���$��0�B�}�u��c�\$�<3�i���P�*=`tK=;�|a�̡�{�c���w��kl,ki�תS�)?Nz�F!|,�(��m���$$=g|�Y
�ϥ�Ŏ�(I�
��ڀ֚���\�g�������3�d�����o�a�@	L+�9����T�KD�	<�+�ׂn�z����d�*�L�*b9���@���-F��0�@��ˌ�*��P|������?~�a��'���L���)� �W�Ì̋���EG��S&>yu�i o��~{]���n[�Xx�( 5��U��&[U=�qܷe��n�2�����ZF�� ��n��l���jw~�=��ڋ�};�g�?u��m�e�B��HF� [f��o�(<����8.VGCJ
�;פ(���Pޒ�JO�e6@ ��ͨ����DL�Q[�ٵ��z�ai�W �h�� ����e�r9#�44d�@�_;�t�O����v���И�h7���|�2��-W�\y�Qs�]�y�q΃ݲ`5��~��^f�N��Q���꟒kQ �r��Y%�J5lQ\؈J=���b�#���'�I ��`ԅ�O��9Z'��#Fߝ�~��yS��
�kf�`X%�}�X� �B�5=�[3j��<��O�?�`H��{����jS�x{P65CL#3O����}P�8M.��'�R�=+13�k3�}���<���l��~�M�m6z��e.�p�ۃ]�L�ØMؕyn��_�lBH����cTFm���s���s�����$wa��@�l&�u7=V�@����Nfhc�2�!*3:�X�W	���7��B$�Y��M��jh��5J���'J�]�QiAn�镩�<�<��V�@t}��h�&dR�_B�7�3V�B`블�on�?܉;�ҧ��T��%��l�|.7�LrBl�x��}��B@eY���ipo]H-�vkt+Yh�?���sRX ��9��Wg��\#$�Y[Jm���x�7�j��'P׭2�0q"��#��GO_��vH�� ���5ָ'�t�aި_!l}Ͱ�NFN-n��UU��/Ч�pb=	�gW��չS��PT�	��&�Eb���K��o���CR��X�Pp�(ڎ-p�lh����;7��E�M����������uv'���~ewx�a���D]�8PU�9"�~{��g��ԣ5]T2�l!�U �g��*� ���l⏅�2p���4x[~i���@��'��	�ﮬ�@
E�}	��ŉ�)w�F�bEl���ֲa��{��_��"�C�I�M�D�8��ߨG�a*��("?-�CQ��F&��1ǽp�ϨZ�h5멜r  Y�� `�V�"`g�V��}k�C�	�WTv�ո�5/*!�RE�����(͠c��B��0�S�_Vܸ�_4,�W�ApH��-�J��[�R�¾��)gZ���F�z��G؍8d�8ce	�Y���o�%ٽ��)�&n���*�m"X񇡱�ĺ%������x�ފ�*˚��ʢ�	�^��d&�ޙ�Wo1KA9P٧�!�s�x��~hO�<�)c��-ju�'�`�GJ&d�Nu