��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P��v�"<ߞ��&'��k%P碶�R�ӣ�sĞ������FY&� �C��/��!����y��
2/��F�V �D��� �a���������4��9�3������>��CϤ�G2�|�Pw?���B.��9[(f�^߇] ����0s ��uC���6���v(�D@$|��K�p��Sڛ͚6�p��ȕ�#���F9��i��JC��ܴ �w�1����K�Y���*ϲ���ܛ��4�p:�A��Eif�?#��m]�K��S�vԥF\r��C����욠���9��eAI�<�ڣ��\������#�`�T�,	[|TҍH��Q`�2���ч���3lq��ηB��7��k��� b�j�1
��14�����?˗T�<Ɠ[6F/ ��|����1�#�l��,����$F- &=��x��9" �KS��]���]�n������&6�������rz\v^�t.�-�9��8i-�3�O|���MXO�N���wN9(\���r�z���Y����Ơv!�y5�@���$��?׎���ek,���ž�֠� -���X�n>2*F���n��ˣ�����E/M:���Y;7M��пy�y�FW�tp�T��E�����#C��� �*�g�:5�J!�������GsSsΫ�=B)"��	��u����Y;Uԍ��X?�$1�|���㮖��1q�*��sR[o��F%.��Ψ(��bYjy�?D5)2>�љWq�z��z���:�J�_OD j�%CZN*$�i_h��yѩ=����Ubj��.�U�8�Ս���x�mFd�4�Rm�u6��h�N�"���^�1�ۛv�%E��	���L�WͱV^�É�`]�޺�c�0:;�0;�
Va���	��곔Jڨ}��6]�ǣ\�(u��W:"6O
\�dO ���MC�
�֍/V�L2�T
�|>��� CD�mkҘ�A`R&O��� �\\�>�&pM]�{�9]*x��8-���������G���H|H�4d��D�2E��G|�r%��W]���K�Ȉ	g�Ml%��I"��;��毦)�����.��~�����\J�������3���2�qFa���z�_�d�c������`�i����5(�|�2�٘GW�ɿi';(�Q�w+�6�'MهS\�`?A�ف�
���CT�[Mn��|\�B�����
�8f<��d��<1��cx� ����ùb7��l]{u?�v��+��.-X$��h8V>��{ݥ��;��!\�\%4��դgL���B/������,�$.�:��8��h0��3�귓�jH O���S���֕�2)C�w���i�'���JJ�.��:��R�8&	
�e�
�b�)C��7urYϸ�_Љ2�"��c#r�G�إ���U���P����W��T�`#o�~�T}����*��]�-O�0���je%O��hnD��yq�c��o`�~�6��`B�04�i�x�o����=�%�:��J�4����?�$����G�Nȼm�͑����Z�s �#�\��G�t4%6ݡeNtϨ6r*H`��/A�/C�q�Y�b���*W��}ǔ��c)��a�o�5`�1�Z��<8W�c&%�A���cue����r_�}K��5S��LM��������վ0��F�a
�<F���D�xR��z됦1�a�`e�F��~-�w�
�xj���A���zw��3
��Ii l��]u��3�)�����m��O?7&�>�}���w�Y�������L�+O:>�K�^��"P�'��������uK�4Fp8�J-�V�d�����%t����p�/�/ �)�5��8����	
Z�^"��Ȭ�xi�mW)���^��+�{@�7�heқhRlx����������=�Q��t��)��S��x�6𭥭����:�9JEE���M�{��P��0Mk��\�+�Q���6�r5�4?|#q6�u���!�l~�e���\�c����� Eq�+z����z�����籅+l�&m��Y��*�\����K��"D��oE�Ӷ%�d����L�a&�J������T/eNB5{�D�5�T���4�K���.�HF��������RP���)��+~��8��WO���������>.����y�-�ZJ�ޅZ]I�*�c���m��w�q@�{qDS
��,d�p_���Z?,DYMycG8XK�U�:�7���T8�'��1�PL�}P��U�]�}.H����NOw\<�"z����V���}C*a��8��^0r�9��/s*vG)2��E/�k���=ݦ��X���pٰ�oA�I�a ��x5
d�n�t�݉f����'?'_\x�����/�51����B׶EX\�1�$��֤L赱!dǸ�U���}_e9��9rJR��N�O|@�A _T%8���}G[�)���:��QH�.���(H�R#	����;�̰�B񏸝�b��ޟ��Sr&����G�֝p%5�Y�v�E\�l�*xӲS��ai�#�O��?r��j"�����$O$^��/�#����V��zl$�C������xY�<�R����Z�Ρ0^��La��d�PB�~�b_\���?��R4��d q��O,p�7vkl�
:{X�4�u��x���hu/x��Z���#��ii��)w����xp��/�����+;9J��r4��jl�Y��ID��p�e8��cj��(�dy�8Jd�JD��m�����+&� ��m���3���%Q�m����3�g�]����,Ȥ�~�&{LN�7��b���Q�2��3}��-��	P���r��胇梶<��D��գ�)l~�u���ξ=��@U+��)fGˍ�T������8`���I��j���s��^��%�q�W�;6O5�N���\�3th��:%��l!��c�Gh��J5�N>��鲑�\�.�u<���.9k��[[����93֨8�2���z�*C�<d��(q���wYV��&ć�M�[r�BX� ����}q?Jv�8Ꝯ5�&�웕	-]�p��S�0��$b� �*ႆ��|�l�dkC�	�y�S��2��C�ڤ���1�%������ߝTa@�sI�I�
�q��5H���v��X���	l���}_Ÿ��H$�
Pj�;��Q��x��cN�1�����(O�:�Ղ
��e8��+�W'U�;�Śd؊��Z���?��`B�N4�U�a�io����Bʥ�P�ZG*��KkI��b��'�y��`+��N���_�T�%f����!�h% ],ܾY#
P���c9�>x ,�0 
1#]G$%T��+	���	���`�|nz����*�@mx��:�|5	aҘe@��2,9���	@ d�2���o��LlD��#��?��;�m����0�2A�f�Aּ��м��d
�`���x�@��Sm\�Xq.3����{��	��c�ђ�Ե����i�fI�٬,-�F)J
=3���J�������`��`S�g�ֹ�'-Ōl���ɛ�q�H9fjJ���J�Pi,D�Wis�2�%�;,�)q�>��\SI�P_��;,(]i���'%ď�����"/��빡]W�U�����f:�ݔ���� #�w@dX ·jbYu3k_j0�p�S�R�o ^���A}�H��ww�_�>�]ɐ.>�����W��a�\i}Ǐ�̞%�)���!|�mpt����=�� �%/�t�ƫy�4�ݼ�D��b<ڇv�=�#�J���ދ���
l�{Dw[���@"�����������B�@�U$�<�_cAJF�T����$C�{����_�mjZv�U:�tr�����U�VQ�t>C�Y!��f�4�Y����З*�&L�oz���uA
بI�!bÁ�Z�R>!��y��9�K�ex2�юC�9=a+
��h�Cv�b��Jف�����e9�Ӡ����;�/t��V�>�������6k6n���H�1R>I���豬O3��c-���iʬ�x'v;)0�fɨ<��7�����b�#H'/Цd���<�x[@`3-��L���P�5�$>��h@`YҔ��9��C�(��>u��+ӘG��T��H��/���z�k��������2�|=��Z
d����X0sjaD���Μ|�"+��:o�pO�'I�KH�"�P��۸���Q`#��I9�uQa2���a1�o7k��Z��q���[�%���=�@W��2Zu����7"�Gd��$Jܧ�eR�2��������B[����EBk��M��SV��������]��餹LuLt"��&A��׿�ף�Pɱ�Y�z��k;�{4Ш� -�� �e]:T1��5��dX�$������!�t�7�Ph��A���n�Q����ɵ��eI��q?	��vP����ѫN]�jf����z��s������h�Q�Ī�y�����������~��Z�����^M�N#���ږ ;���Tse��[{����� Z�|�l��b�]��(��5��9��~n����=�e���	�����ˬ��/D���P��O?��2���l���c�� "͓��4U�yknmua�C��b�ALs�!7r���i}���[��س�Z12
�c5��~�����o0i�1��z�e|$�%4'K�d'Ŭ�K-�B2������5_�J3�x�iȆ�����+��<���� �(||OT����>Δ"�7mx�"v�	M�������}=���P�����D~v�����b���'%��yǐF0�B8��7�|D�ۑߓ�+���Ç"l�Nh�dV�U���{�!��fe��*��K�����Q7���AwӛJ���W�֒��N���q\o���o:�[�0C$��KW8#3s��y��{B*Ծ	e��e�����W����(�y�<>q`�D��l����5K�Py�����:b��l��ȭCD�
��ț>���A�������*>A�W�O�c�e���}9�_��v}��b���K;=H�ڔ�vԳ�T-^�]x�˖�|���ќ�)�?ą�g$��
�f,�l�Nܫ�kxZ*�1�/X����T��>�%:���o-bp�������#]���gt��"���>i�Vt&J�"��_�͍D`�7���ü�����)�g*=�
w[�S*�+ʼ��:�t�������4���*Q�~Yk���H���U/��硊F�(�z�����$9�o��H{��Qߟ�YP����w۸zCf켎c���j왇 n1>�F��
ҍ�H��Б�	��ꏢ���Ȁ���)�+C��H��Gn95A	��q�)�Б��Э���c�+�� `�[ܕ�h.� ����3�S�����j�'y[�&�*�;�������f҂G��"�\��1�-3j�I��HJI�y��0�G�S��u<[f��6!������z^�֋���w�5�|z9�T�]��e�iK&!�4�i�S힅���w�/T�<��[���:/�lS�<�Зu]��}�7��~M���x�Yf�����s��,�[iv��H���'`o �)��rk��)}��=\��uw$2	]��C�ȷr�M��zW	B=�J:������*hi=��0�a�Q����^ʌ�R�����JV�:��T��س��?����"pA'&��s�	�TUV�n��&��W;�0 �^�k���7B�|�{m�'��(g�J�b���,uq���.��5[��L�M+��`�C]M�T�T���8Tr��2��2�u���0a��y�^�	�G��l+�u2yN0�����=ݹ~�3�;
^+�_���Y�m<L�-<F�[��H޺��7�'���b�-:���l5]8[���7����#�q1�����l�O.u���&�oRD�4	�o�#ebR���0����~I<�#�V PK��Լ�
�z��!�Rۇp�w����2'\վ�z�P��.l���:��+1;�6_E=�;��i��gbj�Q������^�����r�kѽ��i?�!<��B�]Mx��5?R7��R�u���ǣ��Q4��ܞv���aQ����k�f`5��t��4�hV�7�C�	rX��bHa��G;�B�
�6~O-|�g��%~�<?|���Ejdoo:B��<��i?{W�����L�$J���	I���7�|�]ORw��<xj��"���y7Lʠ��`���&���W��T��Y-3��h��QXż+"�4��S}N_����~���M�� �ݯNİ����u,���l�;���i��J}�w�],Y��
+�5����$o�4(Q�w�A�L�(�5�f⚏�4����Ǵw�Ϋ>s!)�LT���_��QS�%�kٟ��;�x�OU���S��2������VV	ԇX�]<'����4l�
�BE�h6x�?���rY>�ؑ�D�m� ��Fg
�2R��)�ܺ00����|�w�����z?Dv�$(c��T]+ړ�Zg٫�i�^��Fp�������k�}@S,<��{��)S�lk���Q~�؉e�c l��䂀�w�ET��.��j�R��)O�#�U��u6���p2���&�:�h��S� �x.����^4ߒ�I��� ���5'����ؔkA���������ըLi1��l��F��v2|@����%K	]�z����T��b���-��0d(N����^��c�f8A����筰�ڇ�KkH��v?�h�X?��U�11p�N�b�R�J�p�Q�E��u�����7�Fn�h��3Ǌ�5�;�%!: $̏*>ߥI��~�ɉ�1�UAqp�6��q��z,|����Ξ��1�̱CV�,v)�sn��8�A��$ak���2w��<�-�q�-�s��t��at�5P��2䦕��g}z��,7	T
�T_6W
�m�����Ԫ�\$A,�)�0��4�Z�^^�Ŗv���<�����8��F����l�qÈl{�
7�a^�kg⃔p)ʓD��߳�\5�ۜ���[z'�������p����|�s(�P=Ȏ�bA����Y�� ��t��C��y�h����rI�]�?q�9p�HY��;jP9����ML>h�8^Cv_�>9��2�1I��ⵓ萬"�y�=�ܫz#�k �C
Ո��p%��.�K�RU"�x� ᜹+[�{��{�Ώpo���A���Og�ܓ3�Oқ�w����|�eW\��*��į�k:چY�·z7p�$݈����n���\��-��? �9�t�d�e�}��� �����,�>!H
��d�>�r��-B(:�ا�~=X+�˅��j\Z����+��ۣY�sS{?x�i%]$�\�|3�7C��ON����58).v.h,W�����Ҧl�����6��	O��'���r�b=|��H���	����U�ͦ�0r���G�Tj'/�����h|:��I��1�l�(�"����2P�wE��²��Y��*�餭����wI�֥RQ����"I��Wˠ�)�YȬ��ɼ���~� .
M�T�H�.>CyV��]$�7_� '��g��ٶ(43Ǒ�$ieGY|UR�f�:����V�
|���G�{���X�EW��K�A��ە$Ul�b�������t9�	�˛��Ff���;%t��L��0��}��'E�����4��*�����֋2F5���[7�y��	���K����Y-s���$g��`�3OGޖ׼I�>�3hMQǓ��G>��\�ʪ������+�����W�'(��_fU����Դ$��WP�YW�6H�/���6�`
U-g5R)�f�\�uO|ּ���S����D�G�&Rt ����\P�JC����ģ艊I�mo�'���G�-7�� N���g��ջS�n�%w�sRl� 9���/iK�«��B��TW���%�Q���|�Phv�*�k`�ꮄ�mU�g�;p�F�~Ȏ��|��Ct���&��ua��_$�?�JVQ�~�֒��w���n��Bǘ#���>pq�H�z�?kaN=ZQj)ڒHC ��A;��.�mXBI�st�iw8�i$>�p)���d�pn�|G��땋N���l��~��������F���d����Ʈ=j
F�8���8|o�H�B�g��H;<2:(�?��XHӎy��OQA�Lx�s��e���۶��������|_*�z��	�iȯ�;L�m��h�b��v�/z<	#pPj�l�ڽ{[����K�q�S�����l�-��O��gb����R�$Gz�mʅ�e`c`[:�GC��C�K�������ʜ�E�L�p��Bg%U�57 �{_v���,�:�W�q����h!�n��j�_�=��V�����M��ՅdQu�w��y�.wF�wV^��YOh��F�<�@��d��1������3u�9f��������0B[�|ip���;����(�X���߳B�һ	�zC����c�MhB��%��rL�N�ثa'��Btf�9yffs9Eӫ��I�>��	�T�����E������HU"��:�/� ��ܢ����	OQ}�:-���6���X��ׅ�2L3v3�a>��Nv⯘�\
h��%4���GAF7q�+�b��(��E�~��@ʕ�˖������)HѻO���y��ܘ�|V�k��M�� !�}����o��Nk���g48c	 �W�p��h;?�K��~��'�����`e����`P�H)T�y�T�Pi*ݶ��{�k�le����a.i�]�^��N�qό���1Qw�����0�y�����@<J�+�pѩ֧�,��P���2���F�z.Ӆ�J���-"X5o���U(�y�=ns6��g3۵��f*�	Y����!����*g�S��&q�����$�-=r���u��f�j;��� qu�ꚷS��tD-X�h v��[&p��-�ur�wЕ%���H;�f�99P�1���#�-JYH�����j�N��g��l��5�G��xX5��7ej��GŲ��	�7�l�#�؀n���ˑ{q	�~�#bx��c)�r���Lr�1q��C�����&;�Cbg�O,�;O
���{��R�L���S�)���,S�IlS�{�O��;r��cKh��/�k/���1ݵ�3�ų�Y�6�l��ie9�+�'Օ�4ȼg/�t��
��1�����*xC���Rf�Ԑq�f,T�L;�N�;���.`7�zI� \��T/8;�pAy(�JV��M���u�j��[�C��o�Ka&��1jz�Jc!㼪���a!��eʳ���RUu��}��ܩ�	SG��ǐ-,�Oc�B��Q�fp��k用({8�4���l��yǩ�j��6�"'�Қ���&<Jd��$.�2���y��C�L{� �.IrT!�w�͎`^��\����[���3���_��'
�(*�s��Y�u�v����3�:��u�A��x68Ó^�%��PhZќm�@e����"�:Ex��f��,�Α7�(�lu���?�`���A�v.6��]�'|��Kį&��W,�yC�陳�{�_x��hZx�r׹=�VA�#��c�6���r�+a��8�
Z7S�"؞�g���S�6���E���@�0>�/�N��{&Z�Dkn������@/�?j���yDo*�CQ	�{�k�n�� h/?u.=u���`���;�L�?.��[���S��c2J �QNʖu�(�s9sp�1)���_�V�wbT��b��6�}�������ɑܯ�������
$G`q�ɷ��i�n���8�e�����mgj�9�����j�f�<�ҋ�IIH�O�呤j~j����`�̩�L|<�ݣ�"�-��{ oc3J�����k_�kG�%�!P�~�"�
u��r����ף3 ��k��ݤL�}�� �T��H黁��`ɋ��~5WT������^���-�É��$.f.d����H��hm�R�{���u��I�H�_ғ
�]y���)���cR�-`e�֜tR�{ֽ�pǪ��C;����H��/I�xR0Rq���#���՝��/8��R�'��c���
-��ڨ�ɐfP��F� [x�v��p�o�nW�P�H&Đ�/�#����p>ߐGm-�O���4��+�	��,�����b�����K�5���B���@r��c0�:fE�P|=�����Eԧ�Z���=�)�cI�`|~n)Y	��-�xW�c�{�,��p>^���&	���B1��\�T�s+��ֹca섥i�A]�ޫh"��F[� m��A��A�&�.Q��\>�b_K����.�!7��\��� >� �럢�.Sz��*G%���N�����~��|�%�1�A��3�=m�Lp�^��|��0���`��I�Z,�����{�'J�+�OĘI]�e�ѐt!pM����AС۝	�P�;�J��V��F�������%���h�q������Q��)��mq>���_E���#���JD��?d��\�f�U��-f[5V�uˮ��R��"�R����Lw[o1����Uu ��Y���ú���{���Cp�/�Ҩ��]ј�Q8-�*F�޹�	|��bX����3�_=M�×�����U�e��i	L���Bp́���B�*�H�s��J�ٸ�pl⚚H�4՜�H�;F��6y�#'�Q�v���g^x�]5Z.�O�F�|X�
�o�vӬ��I)"��:�_oǢ돥�#<ը�)�kI�8J3��Cq/��_��gW������b���B�eQ1n�C����5;�v}�6x�W�Ɋj�hU���*�:L^|w��X<�r�f��+�TƎZg�wP�)�7�������S�v�"�p�q�0���iI�mՎV����.5X3�a��H��$΁�r�U��J'U�g��l|1���rxXA!�s�
ӥ$��֣�A�d'&�A��3a#1���;j�_X7<����a�L��b�#a�BG��U�����T��`�_E(���A�%|��9�i)�y^�C���[~o�����+v���A��>��te����w�a�#3�~�^T��Ŷ�����gb�ٺ�:j����ľ1H"�b��2"	&0��FI"&T�$�}�X������IC%�`�5��g��������R�`}Wa��"#�C��~I���3��K��B&�ӷk��yp*$b�)u�(�+�u,z�ۄ0������ъ_c���]PRP5
���~$�b�;�D����M���\tc�8ik�2O_�s!S�A��U����k�U+`^�W$�q�m!l�R ��Y��F� R�UJ��:%d阯���#�Uʴ{Ŭ�!&H�E8�mao�檗ԯ����paY>X��O29�71��t�-��L���/�U6���P��}'S�A�+�Ơ8�Kg�I�؉1p*�;�� _JȟJ�b��t�q��)��i"�1���J��/'��EZ��^-bC�~ ^n�������n�Z_&�Tn�e����J�3�R�e}sI����P1"�e�Q'��W��/e�2���^+��:ݍg�U� bkҺ`�M��W�4v�6t߫S\��9�^�h�u	���%��K��P��D���]�t�W������G;WR(�̟]w-�8��ޮ0�J��,w��Qj��'�-ҽH=v3����dw�U)�|��&I�����xA>�'�!�h���[V�KjNO�nڈmQY����_
����=��$hp�[�bA`��[�I�Tɡ�R�t�پ�{wӦ�A� O�j$�Qgs
�l2v	��k 0�r�vL���NI!'�����Ô\v�g����;q-j�5�9�ui� �D�t	�[ug~` ÉRI�8�������ѯ�c�k�	�J��:���**�p���Y5�X�W��?^��k�$�M7��^�&��X/�Tw�%�4r��rHPy�c����\�o�s���4z��[~Kܛ]F�	��d迪8�;	+AW}9��?{��Ѫhꠙ����F+=�_4��J���h����?�B܉��f��Ro����@�Y�݇�	���=�, U�?/����ɔ�c�Ժ. Ι�j�۟F�6�L%�/)	g�����٤�M,�v1��Ζ�>H���i�?x��I��K���$�S��mAP罠B��#o"g@�]@�t���c�Xf?�
�h����C�e�Z�f1�Ӭp����������  �����<s?
�y���pɯ�&�|��Q2���)3�U��<�%[s��c(�F�=��'�o)�W��r�v��d8�x�j���ĔLp�&P�hBfJ�لcӦ5��r��ҵ�ҍ�E<��[�c_4�yݚ�?��q��SK!f�-�P$�{iPإ�k`,O��4m��?hv�ϲ��|��TKIp�%�_+hI)�8���.f�F�ȋ��*�Ai�ln��qq��܎3�$�k
��a�h�x�����1mDT�3��7۵�fW�Eb���J�:o�Kՙ(���O��Z����f�t��%|3M!ܖ��\�B��V�)hX���>����}�ceUb<Ҹ7�q&�e��^uLF~�;Cx|���ҁ����� ���%�Q!�I�e� �Lo�
�,+Vv��GB�R��(�ۉ����ܫi7�D
V�7�V�
�o9�|xM��[�������q]*��d�B��\E�������Sd$�vH���q#��w�!wG$����h]+���@��£/�!S�ˑ;��&Ħ y��!�@�WEp�K�(ܽ������+��ޚSC�_�}o�Z��ZM�Z^vB�+Lx�o0�]�SQ�ԩ��r� x2uFe��͗�H�V*����{�Gj$����:�L��Y;\A+L��*b�gN��t��z������6�3��Gw�f-V��;	
���Ə`��*�h>-3 �0��䜔�O���p����%[}���%�4�4��V��R��!�<���_P�O&�;���C&�?�=5��|�tU���a�ۂ8.U�%V�wm�W�|�nN<a`=�l� �؟s���z��y��k)�*�x���d��J��,��>:��,�HA�jf��F��7���� �;{����Q�h�~�w�5�/�4CMwx�ѡ��0�X)� �<G
�+�z�[N��mzyR3���"�t�Qz�
��R�CM��혂d���ۃ{
{���#b�$�l�C*�@���T�*U��zSή���R{�w���^M� ��v��h�r���fc������] Դ���PS�'�SX�,p�֛���� (� ��X�(+�n��qp�����\���ez��W`��쇪A��
8��H<*�h�q���o�>�xY;_�ua�嗞=w1�LVCC�ߴ��f1��/�W���9)���'���ӹe����o}���q��Ub.�n(|�ȗ �5�X�(!:�q�����˾���s��mfD([�����߁NS`��$��)�����Q���oaɔ�j��p��yD��@�s���A@�"������>��'���)���h�+j��ú"n7�t	o���j�c� ����So�=&��w���6�>/B����e?F�7T�]�uD3%1X+Cy��J��=��B�ٕT?J�+����ŵ�S�����.J�с��`�^��9���;�L$T�����ϋ��9�PTْ�oLGV%�jM��S�1�WFɼ�U�"�/C�ɱRo�!x���N�Ɓ纗�E��"�'��n����|[�����d���������QzzŻ�ʹ+Ke*+����n8��p��e��䨫�~������x�����F�ܝ�Ef{t�{�BS��D��T�P87;'Mn���!�t>����|D^\�n�8T|�2�W!�S�����vA�xGZ�=n]�k��3�BC���l!�z\� x���Y*?�e@��a?�����D>y]�r@��<�#_�cq���#�xY�U�
K�n�G�6�F��8ڂ���"ܷ�8��.ٮ���D2�����|F�=��\�p��?/��ˈH2����T���q��k	�&dQ;���h����Ѩ�~����;���Up�o�/ �k�d���e<,\�11�Q�"�a��apb6Ke�N,8�l�]�|���^ݫ�B�>0�!�ӥ��O�"D�;�`����N��( f���v��~=<��5GP��^95��c_�1VU��f�n�X�n!����|��wl+�y��P������i��T������I��2����� �Y�?'!�{mY�M�U&��x�Y�⸬>��6�����z5}y�<��t�����F�wjp��H�s렺���Ĺ��Y�d�j������ׁB�`	���A�Ě��@k)�T_��0z�-�dY���eτ��tm�v�V�>r��n�����-��H��(���!"��/��OVC�Zl��q:H�v9e���S�Y�� ���?���^��I(v�#��_�;��6�cb?]����y����[���.�* �{�<t��HW(�vC�.��k�,j/�u�z�	���MT>���C~.����R[�)��-5�K|%�7c"���rl�h�[���*5�jo^�6��ȱ��7���\����d9�2^�\p�å�Lɓ.M&�u.�?d�։-t���Q>�eh�^A1��r���zy\664�.�T���Qo&��b����ʖ:W��{�2��ޞ���0nl�V��&ه�>�ŀ7#���u\��d��Q֞{��IJa��S��-dI�������0�ó��i��>���m�r{�ԡn��.�7�D@,��tz�4}r\?]�����[၈�p*�^�Amj0K�f�������X~_m,������|�B ʵ��keIq��_�e�v���A�>a�����:嫯͛2Q�(�&+��팿���[�X�d������H~�M��+ڊ�Jq@X�Y�6WN�AROdV�֠�r��A���l{����=��%Py�W��'S�^Ǭqlvm�+O��@/�A��l�
x��ڏ#W��^R��4�?!ʛz�\�j�!�5H��+��wl%�N��zɝ�yĥ�������wS��$�%�aȸj=d5n�XJ��#B}Ujq*�|���-s`&Q��)i���D���s���V
76B7t���G��;
ݦ~�Ud�4�-�Kľ���S�b�kj�G�N��T������R�D2�ђ���p�50���Hpm_�W!X��+z��*Na8�fI��Z�*�������[����d���S󵬟��o)�;U�D�i�|#X�6N6~��/jp�����Y����lZjj�
�u��Iюƪ������oQ�B�1!�Ǘ�Uyj�1�����o�L{8�� �AT1ˤlmEX��������?�.������yL]�k���%�gW���u�S��E�8�/��rp����BޜV>4�[.`���J�O�)���=5�?��T���rlqca�u��5�sj�\�"9)�r�w��/AX`�Ѻ7l%�.�_Ƹv� ��R�<`/j�l���IO��<W����עj#��GƷ�����M�#z^0N	b���rg��	��A���%�-5jm�u�b�5k&�T�� ����+4���$��l�[��ְ
�Q��pӋ�N�Z���ȉy�W"�������ly^,7�{$Ѕ�[Jk?'�ٲҙo?pc�p�4��B�~�����7i��D���=�z��M�� gF��Hf���}!�.���Ɵ6��mJ�T���UrNb�a�1�k!�X��o#�-u�9�f�)��*B۷�`,�,�X�"�����;�HcBV�̹0a�1華o��0r>%�n{�@w�\����Q��ƌ�?2�M��P$�Bba*�B�rS� Ci�C��+�@�)�yKk��w9.���2]ɛMa6��|h�E��x@��g��m ̪Y�����ꢰ�U ʙ+JM�TKM�&pT��뺋Z���;O�d��o�v'�Eʀ`�j)�E/أ1�0�o|�q��u�]Ɨư�����C�\%���~vqc�}*^�KyǶ��kѲ�KW�+J�=�g�H8�7p7�c�A��h@�e�6��m����cun�$��5�w��oj>�����6*��]$t�:���Y��q��Z�K�����79YS�Q�Pʉ����
��l���36㧴���<�2��梲jًҡ��?�b��dȯdf�X'��a��:)󣖨ü"m)(��>UÑ�M�E����I��%�Ĩ�&i�b�RN ��<��
�y"������<Gճ�{�ޞt���8�1mv�v0N/̙��&HT��\lߝR|7pQ}J��~oe���Q��7%S����}�F�kALX�ޜ�����c��e�>���j#���8���Ao�<O�������CW��5�T��J^�\�U��Fa��@�7��JD�(�ʲ����e��"�
P�N��(&懺����L�Fן���l��n9�C�WA������08�Cn�l���ч���F�D�%��;y��.��Z�0��4T�VD��=o`�URFf���Dw��G ���Ej�(s\�Z01�r�v
���2<AV>@��D�)���)�aF4h�3��g$z��ތ����J:҇'��G�d�B��Mt �o�	Ӧ�ZRf��4p|6��n	���C�bY���f�S�(��=�;����iYi�ߕO����f��荆��{$��(�JW{s�#U�q�o)Χ�X��"e�����rMӿ*�ۙ��ٶ7w:�봙L���	L!����/|�p��s%-�{�T`��S�6����e�k5W[K�V�(��_��c=�L�[L�b�A&��p��]�C�FV�	#���qx GLva=>\ +v��9����
���D?�"H�?#���<��'��y0Bvr:���{{��0m�|r������������_�)7�Pf�A�$C���������@V
��1�ΰ��>n�<-\�/���P��?>؅��+�Y���Q�刎~� �;>���'���u��}��?,����fDF�� y�A�5�G���̻ݭQ�(��/����Tv����\�s�~Ђ�Jhz�N�dS�jgh$=��uY�n�9m���}���.f�.�S���k�������}~��P�� @Qo-�p��HP�;�']��H��`Y8�q8D�{Y�Z{�.c'��Rt�rK�ʣ�� +��ǒԞhN�z*��S�X��K!R*����ldO)Z[���ѭ�D��6I��Y�֪���Q]$��}��T��ۅ��S9�� �4�x�_��+�2��s������"�&�X�����{��t%:m��O�~sP ŸL٦��ċ��̰r�I��w�qɤpx;�ͦ��cgl�(�qBX�<&�es Ƶ�����mޭ�[Z_[tI�f0ZƓ��7V����^�_�ٌ��ha�#�[*XK[�~p�?��ct�|��1x���j�K���7�i �gLq]�,ttf/�e��r�]L��n�Y�����C`o���WڤjF�|�	�6L��g������F�� ���m��]4+��K-�H�u(oF���8:��Q�G�{ٝ�1G��
���T�oPb��z��,�YpDQ��5�k�r]%V�՚���i"��F�ŧ�e)�u��d*ڠ�3��B_�Ӱ�9�y>Y����hy��],30�(^�[���H* �Ų�}(�<i�ܷxc��4#����GF���UY[��{d���ƕ�.֢�e���In.q���������w���v.�2*w����0���cP�&X��ȑv�������5���=�:�h�GyS�Wom8��T�ޕX�#ŘI�s1b�2Х�&@Xaַ!H�@l�R��8�s��:s�y�)�j��*�Хr�rRT���̳fsMI��h�:���Dl�.z*��+�nk�lb�l5z�o�Y�P�W7��G�����n3m�3�FN����o������ݠ|��b�L˟���*r�K t����d�����}|*�D�Ie�	`�E<K�_џ�0 ��k��1"K��ƆϏ���,�+�p9�4�g���{u�P̫�p@j��\�c�*�0��)
�{(��Z_�0�n����9ۥ];�=m���\�kn2e��s�*�\o��,l�(f�l�E��%�r~k
���d�)V&�w!aE��VٺƧ�ev$C�A��/�@�0L���.����U�K_� T8=�Hic�N��	ư�^GUO�+w]�TG�.��p0C�q�&�8���hY�}�d}�F|`��U/Q��Hz���'Y�P��[���>\��J:��+���	'!��0�7�D�����ǶsyD��w�L�z�B�Gd���
���,;6����3j��H��8�G���q���ۙ��H=���}�lgHÅ�H}�{ޮ����T9"� �T6d� ��� 	9H��%ǅb������6�ѳps�O-�:0yd�έi
���om��(��v��a�}��(O�}�<�{�\�v����yʹ�DʍEb�Z�?
��ښף�j����Ӟ���-���@�|}"C���E�}�=��35���E�Wi��r��uOPJ_�$����R��xJ��,��n��a�Х��`%k��lz3?���[C��9;�]��1�u�h�d�-;��s&�vK�B�W�cF�K#Ē��5=Z��qX��A~<�l�o/��P�������ءN>s�����<N�q�s�P8i�q��,ø##���d�y{�C��'���@�yGB<w���\�\��Q�
���U�AT�?����g�n�;���5���i���F��*���j����H_��deV��lU�=�NB�:�͐���8��)�G�rѨ�@*7&?,��c��h�Ic�@�G(���y�҆9]�(L�3ӂ3|�P�-ΉlNC�_5������5,_�f������Q��w���m5�,"���+�=�#q������U^]�1B9����Ջ.Fb=%_n]Ƿ	V��*w��a����@����ݎ渙 K{�8�$ˍ,{'Q0j��\�&Gj��]��\Ի�g�����񒮒��Ʉ����3ҟ[�rn�"ntW���y�
�,Y =$(b-�ʽ�@����In#z�u���Mv})�X�g�i�%6�Z�8��wK��]l��Œ)�^f��+:v2���o�K=ݻ���@��V�>�v��x�Y ��C�݄ ��J�?v��! �R#��j�,�U�}�m�@n���z*��L���K��}�Ӟ+���3���֯�#�
k(q�UȦ��Qڃ��Ђz�{O��u�A��B�C���7@��B�\Eża�f8/#�=��^��.|����w��|���a0=�:y�D'�LJ)�a�����!Lp~]B��sUO~���T�Y�l��UZ��|w�z��+�����N�m����y�^��2�w,��7���Yv���CҜ�p:��,Ȭ�4i��0:~�ř��?�S���O�F(�^�w�=�>�԰YL�	QL1Xi����W��®�*��#@�J��� D//���ƫ$;����6��ǖ����g$������`� ��u�DF�c�g�L�������j�%ǷCUb�)˺��ڽ�����vA�rB�'�Z�H�;����h�� �EL� �q)�=ˎ�+�i;�ET쏮����� �J43��!%��Q�S��iJVP	@�<�d�ft/�v��<\�� Vjx׵i���|z�Q������B�kO%���+-��.�s͌�Vs�;+9�$��Pn�&��u�/59�k'�7$���0�j=���|�c`��Jl<;cT��9t�3�W���ՠ<=��� �?�D�k�0h�me��4�_����E���=;.F�&�n��W|��
{b��U���O�qns���]K�����o�`��QϳC{@l[�����*�}ǣ�oc]��E���4_��e�ܮv�e`�/U���G(�"	�X\��n�-_��/:Tu���>������GA���D�.���U�i�[W�z�Gy�������(,�SG^|s��w'<.�C�f�H�}l1%��tj;|�Ca���C��[)�L9!����
���W���>�zh�f�أc�&V�|���{,ޘ4HFd�c��;;\�8,��8��A~��bR6�L0����5I�{��*z�]�:�!+���|Eue�3�i���G}:���GHt�Gd���fF��y��A�Rǡ�-�>�?B.XCQ����&��7�m�'�� Jk@�,:B�H��tj���１w-��վ]u1���Źkg�ݛ�@����]���b�my#�f�/2��iy`��o����������J��>�Db,'>��C�e���[�`}�<�t�@�B5X��Cͺ,Q�y"��H��l���{5��Vrp*�x�Yj�t�L, +�Z�V�G���bPˠC���jKE�tb��Y���3"�p��O��x'\�!T3y��S��#�- F�bG1�7�y��
�b$�rdY]�����/2/ �y�H�Ԏ��>�Rl_�����7Ov����*.�5v�_���:�5�h�)�DADy.�N��b!���x=���[*�_�O������9����MҺ���r��G�F�x88��Ӻɿw�w�_j�f���ž:N�2�X�� 4t�z��!�I��à䆾�FrD�8ƒ�+H��u2pn��/@��6����s���zAf����܃r'}��hs�^�BQ}���e:�.ͣC;��6�Ԡ�'�9�yjV�$S6�	]�E�b�K��77��C��f[u�|)�?,���9�*��%�A�tP�:��)g�hcug�j)R�l&R(~lȳ���;]���Ŵ�յhx�).���ҁ�M�-%g|��$��yz�Ȭ��F򝮪��'�د�]��G��/&���"�s�CF��+6|�����F׃ސ�w� ��
����8��T�)�6�׵�ҥ��RI����yĜ��Ť�/�G�V��YX������3)���ivHm�r�}��u�y�]NU�>Y+P\Dd�(M���:�n9�ݎ��H}��K�@t�/)��ޑ7+�ӠR��F/�GvJm�e���۩B�����P� �U��>�Pǹ3D�9tb�:�#�i+p�@E	
f\�$���O�� X-#X�S~�2�1ʖ+m�2�@��P�I�s6y��b4ׅ�W��@!Ўm"�N��f� �ݚ9`�s��S;���G4Ya<��O��vW�Z���;�~�ȝ�DEB}�U��~s���eʁ�L�:�yo��*�,ی�,���DG�%f��D�`�$�&�ä%24�"���G������l.�7e��y!��/SOЏ���V��U������<���wbC�\����W��GJ߰�"���0���W�)�4!��Z	"�=O�q����S�/oKύm؏-�z�UU��egd}k{��.�(��eǙM�Iz��664�JÐr%�����vb��)[���ńʂ��f�Ú�`f ��J������fl㍿; Uh��jP�^#H�b8�'C ���j��}��#�����/�`I��V��.��vڥj�p^�%NvZe�0�#�pE�N�?Qŋ�����IK]� ԡg:���lm<�f�,��W�!}Pe'�>�	�Z�fw��Е�JMr���K��85������8m�p�>��S$速��2C�p�S�.�uT�<Rv�6� �->��9,�'�q��GoEQ����E��S���(�gh��:�����ˋ"eN�ڡ)�z�X��{��"w�HQ#,#�\nD l��\X�r�)��[`�rQ��hG���q�m�5�D�iW���>m�NB+M8Gd�@�]�q�N\�`���wS5�� �k� $d?-�����QK|<ra:�_�&�s�'��4������Ue��H�����u�x�Jt�!�㍋����u9@�����J�7�]���tb��~@��ӵ�^y��x�
ժT�\�;�ͅj�U�帝��p}QK�y��ړf�F9��&�W,Me�aP���kM��֪�z�<�V��&*	�to�C���m�����[���	�C��,'��Oo���X]!�.�»�������/�/�w��@�U���!���%/�����dh`D|A���M�醺�t1j�ep������ �Z�O���6:NN	~H�~��Ћ)� xD��dćC;{��H�������d�!I��=�F�!D*&�-����Cn���I9p�1,��o��{$��Ĵq���gtz���
�8*������n>0�E�vؐ_���a�K��y5��i�W� t�+Tށ�+7&\�K؉]p�n�@+�E#��Ŭ���Kڔ�zy�ڻ��h�>�BT����W�IQf����IO��;�n�w�q�n���:ńR3X���0�{�������6��9�cޙ�� ���b8<�������u��(��ؒw&�r*����<����
9j�/�ٲ���\�)��RGͶ%�7�tp$6�J��-K���j7���U��ȱ��������PT��� �zZw)�@_���ZR��]����b�r�,�+`�4�r�E��܊��ۑ�?� GNc|�\J��xM^��PB��ϥ\@��@ ��E�r��-W^7W����4�z�V����QI�ڂݨ������mìdKi��囼���+u�#�G���O�եRg�G��=ɭإ#HjY�x��T�r���+��杳�m�s���d/����;j\�6~M��n�R��T���?U_� ԏfM���Z!g��ee(,K���z�� � ��;�Ƞ�(�3T��ȡ�猸nbi�*����\�k��C�yP���,z���2�h,�7��Mj�I�Y(A��ܾ2i����u�%�9+��$��I\Q���ֆ	7�'��)�F�H���5A+�zZ��"��*��F�3�`�Wrhn)N�N߲�@��s�0T��7ǡ���G�6�
}"����x����a�&\A5�M�9��qd��8W�r���ej�T�غl�.d,+ZbP7KW� ������G^��7c)��Ƅy�"����&^3jo��1�,�MQ�Ѻ~�V��bq�KwF.$O���r��K�:l��$���<��g}֒K=�+.� �޴����Ji;>���f�<�2d�Ib�y�6�3�{���^1��m�*L�n�s����h��a&�F��9�27*�lC�R����]!�`
-�7���"�T�{�!�N|K�0C�aY)��!@x����&��Kk�e��A��A��-}��]�a��/7�"����0�*�44�V'x<8m���7������Y������-f���G+�j��B2؝|B9�I�5h4��3I��}��K�Rv�ic��a<.b_�yt�0k�0t�=8��8aVv| ܼ�0d���ZvFS�-&�|��.��q��MH˪!G���GGi��#W]ra�Zy�>���>��C�Q�
�����g�2w�9vۨ�Kk�L��P
��4�P�i����h� �a��D����p�d�_�ޒd*�Q�!�ѹ&�������$��ҼaH�h�$�cG�ҟ�V�&�n7VJ��:�α3M�5�wB&|q�N9ر/�� ��
W�|*�nw놠�m̅��:ԃ�Zox��b*kU��*6�F�v�r�e'�ܼ�tm���M��>�V���`H��K��_���)x���_����N��P���^�������3܎����^���q�竲LpD�.{�q��$#6��Nq* �#׋���[��a郶�q�!S�EϙR��h��E�cuq$h]�2d��6�\a^_|m���V��ߐε�pb�ZE��������Ό���-��D:#��\��n?P*~��᧨��N�C�[G�4�Ƒl7�(n:�=�����RL�F5T�Z��m�v!r�(���"������baI^����pT!V��lM�x�!.�C7k�|��x��ڶ:6� R���˼�)_.ϯ�t*0G'���3,��̸�Y\|c|,�!�A!����,e�����VCM�S�_��,�v8䇜35޻j3!K�r�p?_ ��B/�����q^��y�����Idu�e (�v����xH-��K7\�1��
���N%e�?�o��#��j�9��ҳ�?��PJ�8y��m��N���{��b<&��N�����\�~��9 H���ǰ��Y����y;���ʳ��~'i�y�w��Z�)�9����,�Q8<o�A�xډ�_8�w�����_���J��U�˜�Iy���)��aT3�F���0�,��p#�ƟHZg��߸���|���l$��ó�����.Mw9�X����i%�����kȐ���x�'r���L���M3�M���U���a�`��+����2�[0'�G��B��|�JW���Gi�WrK�<1M��S<��8G@� de4���<�Y$�P�t�h�\}�Z��8Ti�ڊ�4�����ͪ�Yw�Ih(��`���xc�Ls���]*M?5�g{W��U}mY"����ƅJA��v�Q�X�I:2���0��=�2T��د�J�@�΃He[�x�0֜�&L�{1��=9����&�i�͞,Fŉgd"P�^qk��z�a53o;��-)m� ���4,�- �3 V�2�:I��Z�PX1�Q�G� xwb��A��~:�����MJwP�2~n�d�� ��;q!@���?C��iP��F�Dt��O���K*���3B��G��"��5[���$o!��vt���Ei]����/�0+ϫp{�XNf-,u	���O|�|[7���
[��"a�����hN��uɤ12װZ!D3���uOM&���L/�x�r�(`%'�W*�&�U}ݟ�j�������Z$#lD��|��P�4	\6p�Z�洓���j�$�Orv���#v�!�yUQٳ��"zS*�������{�+�6�Fi���FY�a�V�y?�y�s�[����#����e�z�&�T��1�Uߪa+�x���6��r�@qN\�ġ1ňC�`��@T��נ8�cn�?o��7�6���
�)���MZ�V�|ϥUap~o�x���%c�5��yR5�DB���&�H�/Rh��Y�kO~Љtr������Q�W�e�"J-��� ���W.�Ϗe��ӁA�)���/R�_
��8�F+��J/�*�	�]j��ao��)�M+/p��6eX�15ң���LM벗�-������]κ%��HpF@h'�XK.�eF�`B(?��w�}����K+c�"�Z~ʚa� ��^`U�g.\�!������>� \�<���̙�@у���d��B&�+j�YBw��\�>9TQ��.]M/m}��%5�J��`��=��%�`���լNhU�|2
s����4��W�'A@��?c{<_��F/�?�A:���\u`S&񾩹� ��\��J���ʒY�+�uD�@v�UT6e��^��Ӻ��}�@m��mPC%z/v��~
Uv�u�7�`$���8��pȝ��V��s_���9}�9�h+��]_�|'V�>���#ݔ7�5�����d'o@L�_|~]&U���k+�y��#�_�B>'�q�nn�L��P�����E>�ʮ�G��wP�H\�����j��¬U��Im�*j@C~ʮ`)�*��O�N}�V�D��?X"��C$ƃs�GAa\7*l�޸��W>�ĩ�z#Q�j�ڒ�yi�&�Il|��1��ij��EN�pVS�n��_�����j59fŦuSbI6������il3қ
�Rb˹]sYKpR�S[� :1s<�Z,L�z�,Ȭ�Ǉ�/e0�6Č�W|". 5��g��f���o:�Nm�ze��Z��̃MDp��[�y�4�G��Ku<�">z6���� �O��s�][�v
�Nza��u!����q� ��tl��F'��,�7Jq^�Ax�f9���xQ����ݭӺ��	�+��}�s�54zX5�'�	��@!8P���x�ٴ
��M	'V��@������ZDe�/s��7�y	N�N5�'��gě�6h�R�,H|̯��?����VDKw���?��ǩ����$�E�ƶ,���ә�[�D��[�[��%*�-���.R���7��u�W���Ɵ���g"a��"�,�U��,�5dUvR6Fgj���@����,x0�ά�3�V'p��AO�l9��$���'_��'oVLm7��)�<����h$�O[V��*c|�z��? ��3% j�����q�tm>_.��_?��`z�d�+4�0h�c�Ȇ�>ֺ8�n�U��J��4��x�]�1�"�l8�٨�X�©�2ؿ��y�ɒ�	H����S�'b��F�-��83������!o���d�T�c���_R�}~��b�5_��¥��0:��]�1� zg.�=�cޤvݾj�i��Ĭf�{ʼ��k��WN�U��8\�X7�AT%b������r:�N�5��R�� ��` �fA���W�cF���P�����ƪpIʬ��Ǉ5�x#�c{�+T?��{��$���Hg���5TF��F3<����e���d!���E�}!K�T� �.)�^y�h
��=#T�L��i�(wen�wxݛ�"A�k���-���і��egj2��^�����Q��b?�?WD��gM۪���R�C/n��<o_�H���?^��SD�#K�mxo�
�E�^�,=%Y��,T��&~�>>D��yjp-3%e޴׏'�?��������̈7��e�{Xa��I哘<t�¢9.��$1%����٭IŬ2��X �Ȟ��h~�q�0�'/�(`ƅn��h���0�36,=5!��.��1l�,����#(&W"�fu�SA��A��Ӏ=>��f�����b���@崡�{�7�Ӏ����.��Cr��9�cfC.�< a�[:b��3��8p�L��Vp�%=�F���n�a&����2C���Ua	R�����j\^q�a��Q,�}J�پ��Q�5��� ��j��A���*˔�HP8��f��h��`=h���l��ϱ�|�[� *_�-)8�0W�����Sj�2BbRJy���.Hkb{�i����s?n'�%?�%��A�6����T�\~B�� �p��� f-�e_ �K���/h���L]{?����0v[�A�޶����?v��`C��-���o�$��n�ُw�l;j@D��nʣ~�j�-��J_���cߣO��� T/v��+l	2zH>Vņ��rNt�
X7!M�N@U�g�'#�d�)6h��MX�;�'U�j`��$_��Fi�� b�p�Tc*������fK9��(������_��������B�u&�V����U�M��-�#O�sG��]r�2J+Y}Kx���Rn��.�����e./�K_���m;�ڲ�}�~�t�#W�0��<�C���Hgj���,��/�C����'��+@V�t��#�ϟ����^�	�{���3rݍ�>���_*��u �vZ�4SDo5jN�J�����!e�o��7�*��'=�b�]O5�Q��<Y���D�C@�wi�R/�����ȵ B*!��r�2�B��g�L�ϩZ���l��­�8Z=#���('����4=����P~x΄���K*�2q�EO��b򮑰$[]u�!wd��;�l�]�%:]û�q�zc���4FI8P�c2F k|�6�9�Hv�X��?[|�k�� �T�wV?��Ë'�$z��A$M�F�9�܍�Ũ��D+�������w�"�R;a�>�G�}�`\r��B\���ZG��E�U��K�! ���T~�R�XkX}��w&��
��6Xo���F&)���FS�������Eߡ?]��u��������_��aT&oh�",��K�ɉ��C:�
�� m�]�*���5
s!KM9�&IG��T���C��(,�=�_b��a���><����Tsb���J���z��H�A��;�\��p4��Q�W����{�S^�i�;L�b񆋁?�ц#H��@
���Z�:��{������a�h�e�N���3�f�����_B�E�A��HD�1v8���9�M>7��y��Dw�>_j��:��N�L����nݵ\��|&D�u��V�9�P=0��ZA!1c��AD#T�a*���.WdUkӠ��M�t= ���A�>���Eq_������`df*��|xR��i-8K��	'G���-��{|�v�����ޗ'�̱ �-�?�F(��x�9�J{"�o_�|�kw5�1p��~ʯ78!ʁ.S bTc��y-<�ܔ���!�����B��^�M[#�|��MbR��&�~,���^`Ti��iaHه�d����#s$/;�z��m���t�OH����ɍ}�]��i�;ܹ~m�(7+%	?�/�h�s6��O� \y��R^ygt�����J]���c�@<2��2FZ]����?�lS���3`w��pS�T�(�JrC2M�rɼ�N/#�e�|+W�3T�����|�}�Kz�=�0��缇]��8<'xFW��]�Ѝ���?u��wA��:�D��|����@޿��\�nHm����"��$��+)b���N�<�%V�mj�Oy%.�l�6��F	mPCm��U�eJ�f4�<XD-R�h�D�{�s�if_VLD�ԙ/Y��Ҿ7j��C���_�gC�yXF�}t��!�ۣ��9�����7ژao���#Z܅kUi[��1�nߩ���1������C�{�bN�[�~
�=�D��^a�'����Ր?�#S�ԁ7��RF��!������\y���������9؉ �w�����s{?�"M���������MG���M�I�k���ǅ����\�^d�����B��4����&]�N����.6���������0�M�p*�I���MoY�{jD�G���}����q�	n�F�9bgd���ؠ�P��������N�e�1T�A 9l��x�A��l0ܒO�n(�\�oLwݺn�Bx�ޏw��/K���j7��9��X��s~B���d},��٦�6��'���3����b!��2N���� M�Xv��C}8���(i�a;��YF���=���V���ob`��HN�U$c2�ttU�Z��0϶jp�`���Y�?����\8�9dp��'~%lY��%cк���<<�
�4��
_��5�Z�����#sY毷�9���ν��SFA2���<�4�1k��7�v��rzb�u�`v�ކ�c��q��@�D�I�џ�t�
�{{:焄����'^/���tn�U,+B�Y�6�	@��ov��������:��(8-����/j͕^� �Z@��Mz��zw�G��An�-�Y������ϙ8�!-׻�:�Bf�W�X�ѩ|nrO(,$��{^��}�M����f���]c]e� ��%��0:!(�J2#]����=Wm��d�/�$4(ЫR�ɺ��ȍ��k�d����/
IU���l�3����B�qr@��G�KV,0yg;\�<���=Q/8Yr3��������F�����/����Ƚ��/8/j"\��L�u�ż�S������!5�Ah�?e�y̍�����T��x��x��p�J�`��R����>�{������\���w�{��*d������4l�ס�r��f����M'��-.l/˒�2?j*ۮ	�Z��"�DD�M�I��W��S�s$��������
�r�'��r��N�y��^'����x��0����m|$I��-�����'�?�����'rIF���6�׼R�����
�T��]�썔�A쓫:+�w�F�p��i���W4���(���7;으f��A��Hr���CJ �9ND)�Y�ytڐ]s �I4v�ґ�����`��Q���n<��31O�˽~8[�˫1��Rۧ u�(_��M���q�}�U�}���+NQ� �B�����dټ|=��@�����>	~�h�K�0�{�\��|��[M�˫���]�{��͍�	��=��\�~�б>��5:��8�w���b�K�tk2-��YS#a�������)�"|��;1F$����o���l�G.��؆d���p����`�VڸfEu7��cfS�}�fU �H�b0��[U-R�_w+W�J�/����������ƭ���uS�'��Dx����+�o�6%Iw�>B�ԑ�m?��	[�����پ�,�DÉ��Q�xd;ٓ	2�䁶0%��d��?�nioJ�t��������"T4D�l�ˋ�9���Ԅ��
sEꩋ����ذ-��K�h���S�f���yUuE��Y��Zs�S9�ؙ~�}8��fs9�VL&	~��e4�p^��}�I8�+'^@�eFi̸�[��-��+��xH�b�b)�R�_�	��kãy�0�|�".��������:�P����WI}_U�h�	ǧ���Jσ�!�V@�����6�-HJ)wU�ʹ�-y��8��� @HcmC{ ��%���u4K��{�.�5�B���G��>��D��ׇC7�dŚ��ܚ����6�fZ���R��)�dʲ�@~�|��J�n+��/5v�N(7Hĕ���q��C���,d�;�*�!�&zb(3^�v	����s��OR�|���=�)yƆ/e�I���˩�\���t���],��-z���GF9���ўKl���������o�0�5�k[��ު��uuH�'�b���)�4|c>�W	�F�zk[=��l�{F:}�ɵ���x�A�]ݨ�#jr����~�{/�zn������l�.w��g���0):���4��m]r���j0�Y@w	��@��R�Ky2H���)z�f��j��k��K�<�2[�y�p����oԩ�U��@�����B�~�_����*���3 ��İ�-G���y����i:���܅"�����-^ͺG�;ykb��ǅ�
A7u�u������v���2�Sx���5hDt:;ɰ��\�w�]��F�bv�M�=.)1��`x��w9���K4.�|������\�Hb.�:�4o[=e�x�qB�'�Πf5�r"�2����Ky�X!�ȝ���~?ty�;��-�z^=4�vCՌ�A�D�~�yz)>��/ź��)7�Iw�fd�<P�&�!5 �zחʙ<���53VR�
R��1�y��6g؃��K�u��V�3ڕ��uh�&F�E�_-J[��L�aM+������S�Xa놶@C_p��;�?��.�u�a�a���k�䵹w���^o��~�Y}F$��\2��R[Ǝw8�E�}��P�["d�JV=���s���cփGFb�2mG����T�ף�T��K�Al��'�)k+� )Ъ@s��8`��N��T��SL��9���9��/�}R<�`��p���x1�i��aN�s���J���j<�0$�VT�w&�	d
2�y+xh����(���?Oz�&[�H�Ř��2��k^�P���/��2���m�&\�I�x^U�[�!�Mc.+Y
���1�?��h?�������8�d�!��TC|Ay�x��F}QF�v*O��I�3��1噎��ΙS��`Tt	!z��E��7���CM^OIɯY�w�&��)�Z�U�+��i�ݚuL]��gf��u��@���%�H^��X�Խ�p��V}��!���੍q�:�PQ���t����j��[�\����nq��O��M���|�ӿ��N6�!�2�IF1��� ��/_d�Ti��o"�G&9��Q����[������1�\�n���҃=>=d���т߮��#U�[R���!��)� �����!S�TRlGf	@��oM���;??����n 1��&�N�h>n��.�rc>�%ɮ�-�H���?�� ���4��q w�%��~!�fJQzE��6�'J��2�铗}��4?��I�"��C��
R;�,F�������C�HY.s��]B�[��)u	�U�jt���	Q����Ū�O��1"� �Ә��U�ʅ��^f��$Θ����7��L��� �jz��S��B�l��P�q��4e��$߾6��Ѣ.�5[�s����1)�=w�OU��8,7%�>�,������%�X�4<��?w[��NG8ZdZd8	�_DnQW�T��g���yN��l�oDХ�#�y���5NYQrFȸ��T�Pպ�8J�lW��1yR{n8b�J����6/� t �xB2�U��<�ĕs���1i{��cDV�}H^?(Xo
�k t1W�9�=﷕��W��+�5�*��{����ghsV�L1���:+򲞋�z܉��_�@;7ԍל\������`B��ҕ1�y����8�� ��KL	��'�����	N�pzM]��J�Y�+���ۙ�M�^B�إ�&(	���YkYed���1J�h��i�[~�6�l�%�O���d�ΟW����$�S-��6ce�M+(���]%�,H�H�D}Q?�j^c�Iɻ!�r�j9S\�IX?.r�1��}�g�Z�,uq���W������B��+�"`�i2TĀ��
fr�~����AD�YU&mٴ�vsd�a����q�B�A����[��s^0=8ch#;�v�x|�,kE��~�|��U�&Z#pC�2���>��F}Ȋ�U��Aak�ݏ
 ��s$6y�q֮�_(�cytߪ��z���2�X� ��`�r�a��]�On<,#�3���7���E��+;�\��̪��� �at��z�i��������jHP|��n�ߴ\�(!?���Fvdzx�y�&LMcK~6[� #	��/��Ƽ>Nw�Q%�g+}����;ۛ�&r
v��U-��er76�Z�����Jl�WЬgF���	�b;x��x�7髩�|���yw��k	�B�1v4�*�oH�*�q-N��4�����^�� ��Z�!
f�

�F4�u6��sͥS�K��c$H`?}��e/���V<\Q2�j�6��V�����]R���a4.��*�y�L�����Q���V���J�h6շ4_v/�	�'VxB�:�oul�-u�>Ȟ�]bm�_�u!�kZ߸�p��,�Fv����u8�b:��'e~&���rB�����^K��G���}�r�t�^���)�9b8�.>�5�)s�>���dZM��E��U�Q^��FO�
�q`�L�$~�+��-BЬxo�C��?�����v~���,�O|������q���<�E��з��=A��� �Y~#7���ׁ�VG�����>�w�5�:�����t���n]�����d�1|"x����=p�_��5 J?&�x��S�T���?�Z��������Z��cs\��(��3����xb���.���rC���֨�b��%����p�4��=��e��?�; �z�����2�k�m)�Ty	�/f�5�br�J<$����bӱ����z����ATv��P�.��Q�<�:�u�r�b�cX,�{pf��
}�Ų������5�j{�Ý6&�j�(�=�@������T��ھlb���9g\���Z�~7��5��=�x��L6��G��Wm��W�"���t��"fS��n���wK�Dp�2տ�X�"eAlp�HlUVP��9�<͎�7��`S�ګX��F�϶�T���`�\��� �xI�ᑘ,7s����wl�$ά�yM߷p�~��M����|���'�RDyV�� ���s!��ɵ(U���t高BT�p;5�k6iU�Q�N����TKל�=$k��`^�y��A��^��I�J:��k���*���DU��?Sz+Y��
�ˉ`�	|A�q�,-s�ON��"<xA��rm��h���N�m��ˌ��.�Խ2����^��q�L>2&����Uϴ�(��
=&������}��$C�L��d�0fR,�҅=3T��X���l�Io?h���>������=���6�ra<� "�;r�Q�摸\2vs�wꢕ�	�&j=�Z9c�m�H�0/�6������j2���j�z"�[UY:b��\uEl���S!�Ԛ��P�a@i���%H/�F[���\�0Q��+�s�h.�#ϏjC�ݣ��0T��z���=�V��Xӧ~��J��9y�؄���`.8��N�o�ϩ��3�E*�/Y�ζ'Ʃ��q�=���&%<��]]'��o��IB���:�tE�xH�/�W��T7���ƄZe�X�r�A�Ep��댈�d]�	-i\qۦ>80 �bMB����O��7�d��uŎ�dujC�� 1�r��%b�|�'��}y��EU�f�����Fc��] (x�=���D�.Hf����B���8�|���U ���E�?��yύ��u�g|(���D�����n�e|I��|��1�S��޸Ø�x"�����mR�9v�aAWH�r>7-R\A��c�1?M0eSo���C5���,%�K���*�٦���L����տ��"��m8_"�c0�!���$������DҎ�1=M��<�HV9���n�E��5*A��T��?�Ų�v���L���X�iO@�R�~������8R����u��k�f�)�(�Ip� ��-H�f�?u�\D�XѸ�eG�)�	��� �2[���z��ag�?r�6�e���-Fu�5�5�/�(���#`�!+H�@%4x6!��w�t�ʦª�����N��)�PO�ue��EԐ�S`kr��"х�-�.S<�.�-��V^�|Z�fY`v�~{�x�܄$�n����M�.�����ZX"[j��P�k�w�Am�VO��@�x�E��<k��
LGja/���Si�J� ����)b/��5t0�R@�2�X��>u���U����H�e\���L�X$�{�ՂCkYZ�C��{�o���x�y�\}C-�>Ж������Ծ����ԷQ�D�m(��R�a���π��w�R�r�$�-���}y�������$�R�x�
`'b)�i_�w:���V����-1�4Z'r�%H	��,R��dK#�v��[��-7�����/SSv-+LJ�G^���扻ּo��.���%c����ʞT&)��M7q	>�L�U*NPA���Ƭ�ɜ���m�NÁm��kCYN'�6瓓n�@�F�*]�dɏ��l��lk&�NјlY���-k �����y[��g�
��+O��Q�������OO�V�t���֨��_��n/��}�+�D{����muXli8����"�'ɡs|47�Q�H�B��P���׭��/(^�G�3�V�*��J��i%'�mD��ޭyP���\����Z�lm�:���t��֝�TH��)W�^ћ_wJ�����)��>�ќ+_��zѴW`u.w2M���x&�c�MvΌ�0��K��rթ��xW������ 0y�6Z��0��#�f��l��\�	ũm��GL%�^�}�z�׷��9�/`�34���RӉ��阇�� V*���fgQ�L �-��M �fB(d��$����ȫ��{�{&:	�����r�96��N4�Yp\h5͏�+��������o�Lق
#yvRZ|���Og�� �
�e����B9�T�?�=��g�<'�A�	gB�
w�#���h����dԒ�w���~(�k�s�t�4J�!ĵ9y�h�඘A��B�,��)&�:Q��'�/�dSpHnIZ��MW���˕>q�
�Zg�RZ����i��ۧiȀAl�@�C��Mh�Z�������o��7�S�V�1�@��V^N�T�k�4dŷP�&֠��/>,Y')ج$]i��5x����%�@��W'���ɨ�?صLH+�W$)��WaT�q�(d�(��$����|��y6�t�bֿh*8-&���US�ԴⳂ�4N��LFc9Ʈ���k��I��N۽Xg�FP���� �ejr�L��F��w�e2�i/m@�.$����P�.��t��X��ld� >�@8c�6۳38Ԝ�ؽ��6 ��	�;��;�0M}$�ܭX�~��*9�W�g�e��8F���p��}K+Nq�ַ�8���Y��V�ZPn��b��P��<]2-��H&�,�L����0��ܖLi���固���o2�m���o;G�}���K<dO��,�\3��COH�C!��i��+����T�Q ��T��*�:�)��~҈?cݕ�]~��2����!V��b5�ًPu�e���5��"G"j��8xW�5:����zI�ْ׻���:�	vwT�Ԛ���|p/����.�8gU�b���O��솃�	ez�vq��r9q0R��h��ɮy�"����֋��h=s|�	йQ%]5������&^�n�d+ճ�T���.s�t�d��Iǜ�Z�!�Lf��ΘH�a9�ZA4�e�ڂ������9�
z�Z����t;���tM�O�\T������O���<�}�k!a0֔�D?���d5�/B�����ra=.��5�.�A��L7���W � �:5`�^��mjGX�������
f��;�;1NS,��D�A�&����ať��%f�v�x�+`D�XdE��D�_��8<F�o}k����X�B����Ǔ��M>�6��V�+xy�Ͼv���@e����"Fa�U=�*L"�����|а�=�1-�[�E��ց���wzQ[�|���j����vN�: 84X��*%�/�k7J8��~�3�b/��GD����3��.����>ʨPF�	���8������s-+�`Ìi��á���&h`"�������ȴ0;��،Fl�P7n* ��o��g���]c�//)
7�Ҵd��R��A�����j�P��g]BB�m�5�A�_?�U�Ł�7v��k[}e�l�/q�QD:�QPK�W$�\t�u��F	LX�K�_��S����e;U���!)������Hf���q����g��z?X��Q\ҙ!��a7+����z����4�?�u�������]��X�<J����J������CϏ�!��LU�RS�l���~3����iFZ	*k!&� �ˉ�Y� �M*K���X4/�jf˘�T/wN�7ʆ�ny�Vl�	e�*J���:�M�Gd?)��l��3r-�MK0��u.X�uh����;�z�'$`�X��w� z?�&~G٫� =�i�^�I�X2{c�	�~�����c@"�+����
|I�x6�����hʚwG�u�5��g#��C4����`�t���}���o��	�?�� �$򩆔̦�����R��`��c�s)��P����F#R��SSC�Ґh�a��>*~۳��*E����	��6")!�%�P�Λ�q�#A��w:oa���[���)M���c�es��!����q���t$�c�,\�U���Y*_p�KP�92�A���Ų�P��W��	�w��TBa�y�,Z�_�5����n]��}�m�ˑu�٬8�?��&5����TF�l�$���h$��sc�b�?��'���?�	��Ᏽ�6��P쉥�C��h�pnY�B� �q$`|m%i�O�؟�`��G���$1\�a~Ĥk>��m�or��z+?�������������cy�EIW7r���?P��s�3�p�ꈕ���x/�����Vo7w�7����i�������Ñ�ӛ�FD�Xpޙ&,���k����.�V�0�Q�j��:w�-F�Y ٦Ab,�$f�(1mw�mqe:���!|[
-D'�9�.�B�0�vCΙal� r�v���A�zq�y6Ή*��p��g7��k��-b���(�+FZ�M�o�%�n!F�
_��8Kd���u�M��4O��{Xdg(5}�*��2'S�Vl�M����\�p�:�	$��^�[��bK��n~���X?o\�u>��!8a����o\0�����1��H�B/�pg�W8�����*Uc��d��o$="�פ�6�S�����/G���#)(���r��Fy}2
��Zb�X�;���S����a�m/��C�?���XA6�����n�Q�:(-d�p:Y^��U��vv�Ͽ��pw�ӻ򿃻d��Y7���V�π�Y�1��Z�N�0]a���D;%�v�ȟ\�?�=]H�h'E @���@" PK�bw-��y�(T��И���Mh���k8-�.��g@H#�X'c�&����8�)����[��OY�?{�{�V���V}U��PKgM]*eæ�ck�J�Z�zA�ԓ�^����[>�ǘ��<�� ��`$g��5*���\#��5�R������`�
�����kA6ZE�j�����ʪ^DQ^�i%O���<���PH�L?�L�r�����/��<��1�L�r���ܾ�g{u���RL���mk(�F�n�S>���;��"�gs��h���큔�J�;Gz�;�f�Jw~�cST�8ߟ����9�͠]&��g��q+h)��p�`��3��҅���(f���<�cpB������tU��%I�D�!�q@;-yՠWOYb������uaS3���
kZX���ێ���Ƨ��n�l���[�D�])��� f�z*K��ja͵�N��E�t���k'h�y�wfva}AךB��DՌ{�f)�`(�C/�¯K��~��C@s��r�"c��ޕƗ8���=G����~�?����N�h������`�HJ!��7�"}��0��OWW��U�����N�Ԩq�/r���Ԑ�L �y�⁲$��g��i�� $7����� v�R�ׂ��,���n��3ǲ!{G
�Wb��Yy�M%ם�H���\��m�_�6���:���>��i�oj�w�$v���aؔA�.��+�DX�����L��K��t	��x�2�8�Ŵ-I�F�4x��m�z�"���Z:�m�K�D��v��.���P�z�d�a�zVb7�h�d�KU���{�w'�á.������aϹ�+{�r�OA!�8?K��,�6;`�'���p��`S"����y��S^�4�*�{@�ug�c�y O�; �Q�3��t{7�FH�B�75L���!\�*a��mKQ��myy�����V
�Jh鲖�
m~!J�㼍5�DBN���AE3��KrA��8��.<T����"�9�qbQuP7�>�j���^o_�|<����1g���W�<��a����3���(w�x�Д�<�]E׸Efe�8�MN.ܟ\�1g�bi��kE_Xuϓ�����T���e|��D��O}�n	���t(��"=�06��[�D�J��lz�V���v��UA��jr��p/����Λ�Վbƃv`�U��r��
�E%��YG�X9��S�7��<)�"�����̈́��{Ir��ϠƋ5�GF��MV5��};ah��fW慄#��zH1=���y�y�R��� g"<h����l��{A����OM�|��0��mpG�y;��HM����K�a�s�������>�-_:z�?2�!��C�~�,��24ry!�Y���D���uw'��Շ�:N��A�@�n��Zp�3�޵ �l㯹���zC8�O�d&(Sn�_�1�� �������F�m�,Y�g����Yǖr��bתR&�WO��<rB��m��g���� ��X�g�S�%�̱���,p���zo�R~����A�)�Ru{4�����e�x|���-��g>�ǒ0��f�T�%��G��oHIԝ�<iQ�U���#ɧ/0G�ӅS`v��$~,O[x5�r�D�bfw�%.vf_����CWOI��*�]��#��]l�ڰxit�&�q��/�d�%��a��]AT>�i^��4������OM�W���ĳ(sy���������J��5��	t1`��mF�2J������n�����F[�Z���Xdj����^z�*ƀȅ.���L�el��@�d7�%N(U���OV�:l�qi���ع��e���
3v��Y���k!���ܐ%s�z��{���7��G�T���iCO��a��'c����/�wXG�3�H� �Iyx������fy�	�$RO�1��s�>Zܤ�5k*�5�Dև���z)��]kV��q�e<k�n�e��2��3��>�'h\dX��r&Y���QqD:��������� 	��y��\��M�;F��L�S�ۈe�kG"���
�$�1F�h��}B�������C�>׋���]��9h��Kӳ�1(�G����K�qy��K�|׺J�\��-���Ύ�k�9p]697�����^1�2�6�hZ��Bś_�L|�~1T��GW(2.�T� ���̝Y����C�7�LW8��`��x6�d�/trn���k�Z/�j��W�4$3��{��^���"s]?"lқ` C�Z�ؒ�3����>�f�u�,p��CT	ѵ��ʺ�(��D��`>��%���`��2ћ�� �ѬzBU��>���uw�&.Y�]�<ߊ�����8Ҥv=W T�إ��D�:J�PO*�U�3Ipv���0^�Tʫ��N���9�0a�pXY�©0�����a;�:.A�O�CB8���M{�]�bX$��>:܁@9|V�*~�b�~��w�SRwa�n���'��),��!Ԑf����8�e 2�ˮG��
�	�x͙cBp��q߉����	��S�r,ku?�VOeH��v�uo���r�|���)$q0S9�H�s�@6	��b��f�En`ww��uo�J)��v��R�`'3�Iｩ�.f	��Ԗ:J�[�?S2f~��w�U~��t�w5t��i�o�����PJ�_
g ��n�L��ơy��Еq��M����48���"��q4юgT�b"���Q�&NO*���GfX�4��8�b��͝o_�9$��Q�6���n�by?��(g&�^/��U�[p�.�����/i�����0���>�#�X(jɱWǍFf�~�G���f��P�g]�.���)�SL�!�j5�ET1k���i���']:'�T����=eZanz��Wk��&�,�	C����I�5Ø_�z�� 	�د��<�`ǤB���bɲ��N~�"���Х"~�~+�b��zw;}YZ'��`��y���R�X�=��et�U����!�N˄�8��A��4�#��[3[ݓ-�1��c���a1*�j_���k%	&L��YS�i�-s�-�`�Ў#\�l�	��U��G���EZ�;�TK� ����7á���u�E%�&͜UNTD��3�\kM��$�v��f�K�
���?�թ��}��A�:�^uj|��Hct���J֧W-�ӗ��w(6Mq�Z�F��v��(#Z�ejhlڑk�(�2
�痕����$�a���!�r��߈�uO��K/��D)�T%��Z�wq�m��^�t))���R�I&Q邨t�j�ǭ5�>�@�������|mY�t�MqK��L]
$sə��MF�ଂG��i�ig��.7��. �X%�*��J+;Yqk�+{G$�2�G��w�Vqza���������|1$��zϜ��橐�%gD= \dK�{o|��u�)?� �ͨ��������g��/�7Pk�E��H�Y��g���U-�)�8I��QS��pǓ��RE'����	y�<.�@����(��,��"Y�kW�'
��-�ԫˤI��~��,��ѿ��Ky(�vY��� t�~t��H�`7�cJ����P1����߁�ޙ���n�TƘΓD@� Z:�݃W;W>�?�&8G&�������Ej|T"��Y��gے�'��5��7I��_���Cq�OO�"�3a�p�8@&>�<�������,��0C߽ƞar�6��`藧�1xP�|��ܕ�x$Cb���ݗ���b����&%������<���8nmi<�q�T��m������bQ>G��B �-5=x]=�����	��[ �y�&�(<ץ�+Ρ:j��0���XC�$���
��6��.~_'8�Ad��z뛮�҃�/��B�8�6���o��W��sZ6RSǀ1�5��V�|'�<�k؃&������g
�W�%� 2�R���=��������y1�W]�_��d��E@�C��
NN�=�>+$�6c��$��N�=w���/ܰ�1��a��Ȉ���Z+h�Na+o��"��e�ef��Y���2�0-�g
z=߁�Q@�p�%���D�
�R7+�㕄j�����Yʜ���Z#�at3�\3���֍�)]�[�e�+�a@��k�!莆���?�?����t��t�Nx�"�.t�Z�P�R��yE��%���O/�f�Qa��/��H5���V�7� �����+W�M7=��u� �����u��#��B��#i| ���15�ѧ�����WN����1?P��o9K�N��<���P��I��w�� ���qy)˦���]��Q*+w���{#�"�C�fS�8���d����T��2m�	@,�h�)9,H_9�^vw����Xk"���l���b)ƫ�NMb��A�P(�]VIf �6T#��Ԯ��Qʖ� �D�nu.�Ȫ��"x5>��	7(�ʎ[�(Y����ml��rz��J%�LW��T���\4bE�g���-�|���:�46�S[q��w���4���?KC�0��3�]�M���~489���M��ف$��tmӛ�/��ε�n���mRЊ�b�|1#�;dU���Z9E�:2{�ɔi.�ۡh�4�ݷH#=&0i�,e]xH���ˣ�4����%��:�:>9��e�n�xY��NQ}�9�
}�y�&��4�b�	�J�(�9=�-^�+D'܍�
~��E�v]���)��8�8��o�7֕���ы�n�([�م�v6
t���2�;Xt��#��=j�Ij9^���pzX2E_TU�<�&�֞�U��Ą\�d���"��K�����)BS�����pK��d��(��F;ޣ������	Q8Y�!r��6!u���F�P��`��k��p�)G�)G��g֮7��R~�[;$8�z�
��F_I�P��Z*�)<�4B`?.�:6!�I���Kضˡ��s�iԞ��9N ������D��w�KI,�I$w�
y��6�C6�"n�av�*���P6�da� (n3�hfτ�f��y4㷳ֵ(��y.��ǯ�1��g�I��Z��-w�W�u�@�W���Nw�j=I@'���V���;;�0�Z��Ѥ�J�H�)ϓ1���f�P"?&7o4�<��+�̯�K���P�t#�d}���r���!���#1V[����?�Dd���俹��u8@�EJ������W[9��ɱd^���M��q�s�P�)6����,v��P�:X9�+��.�SNNd"8��L;�������&����(��M���ģ����7؉"_5��� @�2@����v�0A�҇�A���#�C��WC�60H�i��0���%��B�Zˉ����W��r]�
��؂1�¢s3��"c5�b��8"Jp���S54���ͅ��~5�		�~��&�:���w���D )����u��Oy���m�U�F��F}~"��z�kН^V����z�5F���w����vp��d��V�GYyV!T�Յh�Q���5Iow�R�-�+���|�r�N���k=ݏ�2��F~'���蚞c�NTQ���ݩ�JV,d��ҕ|'�uY�ۻ`����x��B(M�0�t�l�6���F!��?w���d������=�4bΟ��$���sg�b]�.Î���wr�\�~���/�hS+xu\�L��,��ZS��'���lڟPf�5�}ݛ\���}�u���HӼ�AR4�%��S�8����'��������!G�ƪ00����U�ڳ�ŷ�r�j�CEp'<T�nHVz���G�`(r����߼��!�Vn�&���Q�"�o&Y�H�_�0�fME%.&y���>\P?���֘XI�dEk�y!G�����\�����[�q�rk�F�+�<r|��[��t�[5�
z��;#��.�T����a#j1�����ː����~�߹���HC�L���(�k�(�!�Qmz����G�l��Dx'�u�ٔU�jHƈg�/3S6g�i��0Sk�p����K�и���Kכ�a@ �}~�hf��J���j;#�Ō���l�e]�O��5F�b��)�/6md�l�y�?���U��;b���E~�rV�h���4u��f�QG�H#�Kz�(١���@.�`���F�J�	�c?UV|�K�U ��-�?�zʶ��C�Fk6��'��@�)��<�!�ӋA���,����g	����G�2_�t��C�1��H������1K����0C�⻫�=�v2;`�^�+��Ц��:I�NC ��z��n�쩦��| �"x��m Ct�:���ʕ��h��d�ʧ2�B�����$��:�����&UD���0w��R$e�o�6Rnʍ�]|(��kv��Dql3Q���/����FCNc��rH����T�O�R�K�(�T�M�i���-wl�H��e�����/�����؎�i:p~�'M�'-�^\K�TR���*���N�#�H�ݠ5N�`����#��~�.�)8�,A5t^[N~�"A&#��3A�|}׾�m�(��Ґ�!2FXQ��oOn���˩ܚ��6ٺ�!e*�7���9t-M_��$��h�"��2>�W!�c�����&9�XxFw�yߞ�qB)�M��1����u�^T���s��!.�w�Nd�\�~����4Dâ���ӹ�XE� ��L�X՜� 	lȈ}Ǥ����f�*
ָ>2y�jx��L��<b��]Ʃ�>�_iՄ��hHI�|W�ͽ���zZ��3#n�f�Ɋ2\��C\��醟�h�/c��r��N��m�Nh-2�)��j:j��x���ᔂ9���R���d���_p�&hz��Y�0��=P�׶\�
�'�ߧ����O���Ȫ�ԏ7|�V�X���"l����b|׀��5ϧ�u�]�w�b����.�a�Blԙ�J���Vc�5���B>@���_�|7�w�2��,1|�4A��8���w�P�7���8��(��[S��3�y� Uw�mϙ$`P
K0 �ɚҗ�|O`��-V*��jK�l�&�y�i܂�jȈ�Pvr9���Y�Zf$�� �]�f�uC����$��R��z�� ���g���������/b��c[RpL�D�����P�%����p��=C�|�F7�-���^s�d�>�S*⹊
I�lEr�J��ͭNƅ���*ٺ�*����L�%j��b�H�U�yN��5c)/�qL&bq@y���v�.v�������!l"GK�I^�>�
�@/���nu7�i+�&�S!�u5Ŭ��J�[�`�F�j�j܏acڊz6<{�U����\�-���}KM��6�-��昸"��l�A>լ��DC�����t?�T�&�l�.��g��d�@D*S����T�����gvJɿw$�ɕ�.mw	֋���a�)6+aLPٸv�W�d���O�^A�G������҂gž����,�랶��,u������O�N=�1�+k���dj�l�'�F{"lD�q vcJ{|���@�_�?���Bf�aPL�Ŷ�4��!���]�)�K��o�*).8^���A.a9h�gUM���<Pn��F3ݽZ�c�]�iCU}qW�.��� +ӭ�	��(���xć��-�qh �Ѣ� .(�rry��C�4 ��t��6��6��m�-ʱ����vr���s�[��/��n��F�0�e �`ɓ��P���L��']�&x���[G��@���[�X�������GY)M�{�r�p7��(��\��n��r��Rv���I�7���8M�+h7˝�u�ys��z�����Zp���`wb�5��!������Tw�VB c���jh�{��c�c�6���VyV����6�/�`2�l�2(��T���M�|�e)��z�D��%���R x�Z=�:�	�p���}���>F�_�B�aO�"��0���ܰ&M���/��#�
�!DY��.xג�W~VL�SV?�o=�����&H�Ȩ����P���\(k�se�i���r�i8��Q�S� ����O�Uan�d���S�*��\�_�w�;L�w�;{�]��6��G� ;ɪ(2�O�-�hye��<��5o�
ǩ�?�BG����E��]4�l�Z�!Ou�PX��v�;���j]wm0xi����%О^R�>y��q ��4LuR��j5��A	��~:�Aj�$T���:v'A��dm̿�z�t{zT�C�MH�y:����M7;��>�o?�G��˳h:�1�	��\9��zݞ3j)D�n�D���?���8�6� ���`w���iz���%�Si���	���^��j �xyQ��2Y��*E� �g v��΢�x<�7�1Rт4�@4�g}�𰏴���Zw	�
|��
S�����`P�xSŪ �lM��;�f�"�ݚ�"�{�_��fZ^	�����jg1��^���iWSF��v�3�&gu���-�ƺ�.p���BT�]�p�&U�kF��u�9��w)��a�Q�h�(���D���{'F0���H�i�5	g��c:}�=B��V�4���a���#UQ�n-�����'E��'���#�T`�w{v�a������{����omy��:ePdP��N���E�I�W��$�h&�h��`�"	��=O �{P�� �A0�[Kih����:`O��TN��+w���se?d��~���n��6�U�h-O�����+������w+��ϯ��dp- j�E��i`�D���gx>�BF���]����L���5�����մ8�N�SKD�kAM�6Mͤ?AL�o������y%^�@������p׽psq��	#���~]�j����d�L�$�%f���hll�>NA�^�� 깚��}6�F��j���qp��G�z�hMx�!�;o�Ͳ�P�tb�pf��l�Yj���I`�OQ�o��_���Lv,Q�Ɲ7�,r�e�K	޹A�O	��<m5�m�By�1�Am�C�5Og�z�d��%U�	�]�"���G�T��m��F*{�ns�8d)&~��e���Hf��duVh�{
�g�)��`�j�w9�>����u����	��,��xQ����3�N@j���a��`�8��N����җ�x������!��h�)�v�q_4���F{�,��C�F.Ɉ�����0Z�$ꯈI��Ö���ؓ����nw?��j�S�ʀ�~����hS��@�,P5��+{�����*��*ܕ��e��P�W%ߛ��T)I��6����|�
p�leg���U��<ߍ�����1Cd�t�8�zrH��h�˯r~����9y��o?OZ��p�@p���T�@gBY�'�
�= �r*<��l!t�G~�ef��t�u��,�KB�Ln������R����^.�cū���'�s�7���lY����n�oet�ݯL����IH�M�����w󗜋�X��\����۬(��!/6AÏ/���_�8�Z�B�j��ō@ȭ�P�:�=��|,��?ŕ���E�q�\�$��M���D(Ek��Oƚ��Ъ6��g�~l��v���n�7ŤX��&%�1*��1�/,)�/��	��`a}�%%���}�_n�"/��jbt|N]��[���~7K�E�
>K�I�`�[<�[��� ;���<��P�LG��%��V{�/r��>�9O���6λJ����ۄ�v�r��~)�p��L����%[�(�&��dӚW��meSu��*��c[R�fo�1��j���po��5��Y3:�����w�l���ב�p"Z�"38�q��N d·i_p�7�u��dw���K�J���˱�V8
C�a~;)�S�r�0���m���nJ�/ jD�[��*
��I[a|F�N��V�~$���z�B����f�yb�]�%p�DЖ�$9�oA�8SQk ��䌘$�+\���]�3�}��@gt4R,�F��um��cl?�����ɸ�{^�H3���o�i:H;�Z���ƾ��2 �)�~z!E�
�T��y�������؊�
E$���{jF�5��;��KK�.�I&�%���3WmƊ�� ��GI|�j~���,��4�Wfi�O�/��^�=�ޙ�BÒ�|����a,�p�5�8�U���WD�E�
�0�cO��{D�w��^n��$w7!Q�o��bM~��"�/�:����)��a9pc�w�sʭ��m��EL!�k�3�TkJ0e�'�8B(�"��ON���H�6^n���ȍ�5��ѩ~��^Z��o@&���Z��0pQ�mI���,�q~�o#P��ʩZip������~��Wg��6�͸N�Ԃ⪏2�^��a�B�ğ�5a���r�L�0o�4����C�d(�9��^�	������oj���YJ�#����^�N�������eo���_��Ol	�	��xe�P~*��'y��n e2R��L��T���"p	!�U��7Dk6�Mc[�i'o��)�q}��;��Ҝ-�V�'���M=GQ�$�ue<�N�.Tھ�
}��=�ȧ�
�N�pã�H�NkLfE��c-NzZf��pػ�e�*�2P4�M�6]���p�TL֩"k^����*�&ۇ�LH�x�	�OӬ���"r�[�����i�Ɗn� �'�?�!雩	��
,i$������^T���9
*ɚ5�=���X{d?NL�1�i��څy���EL�@U��wʱ&Ua)�ƃ��Ýhl}=3"��x��ݼGH��0�"�KN��lV������&_���}v�c��9����Z�]禀��H\H�dF�uu=x�3H�W4�@�\�Xĕ�ɹ�)�"2pM��4ڹ9��=��5��O���Э�1��r�W�̣��	˿hl�Ì����=�O�!��M���hŷ�Φ�t����� k��<^r#{��@���@� �[O�<J�3=ۂV��J��+�5�uyW���?�/?�3b������a��1oX}*p�6�@� �-mp6��>��l�î�������8"�������T~�)�Z�y�%�6�oNBH�Z7,�Ǐ@�ԍ�DФ@��s0w��V��N��7��}1v�� ǀ
yk+%�~I��S��J����	f�hW��݇� :Q/�R������V��L<���N&Ċ�kT%Sƴ�|����[�_Ng�ȚZaܲbF�P�/Ε�1c��z��C>8�P~C"�z�{,��Ig2��V'���:�$�i�m!O�b��f���l�l�n�����
Tɾz�č�JcSi���?���MY�3��$lƴ����bt�Գ��J�V��(qO�M��?bBaD���y֕9����6����"H�R��Ñ�l��0pEx��1�5C�=�|ۯ���;WA$ Z�*v?r��ӯeo�3�FVM�5�$��� l�'�����������^�3� h憅��%��̂R�e�#c�a8�w�	tk[�@$�����i�r<qG:y�?n<<f�܅���w�}���
'�t�%x�Sќ��u-��q���OTw�vڿ�76��5x��ٰ��Ѯd���:�V��
�%
/�O�M:�W�x<ѻd5���Ou�����G;9�ww�l�Ӗ^N2m��p'"
mG`"P�y�W��f!�{�����U%��"�ߨ�4�Ouj��&�?K�>��5ٰq���c���jޠ�3|��o

�L�'���U�	9K�|���'��K����[������0�mjW,Gn�̀�v{b�|��^z���:@�}��� �[d	/hφ*����+E�ְ���-P�Uf/��	�Q�&���e�gC�������s�$�/�zV��[}�n����c��Nʼ�{>�~B��Yˆ�u�|�G3K�c���y����D'��䲍-��xSB���x�#��<$�� ,�l֤U�����:�w5黿�$6(���6�/«�_ʌ�ϻ�u�:�9���ٌ�	U�[�e�����mL�}�bu���M�`�aN�8��_ fϣ|)��������䯾�#K]p4D���J�9r����Ӷ�k�V��c�!U��8�v��R2G2O�Z��h���i8���}��!Q���b�-O���"�ӊ
�3�酡�w������gZ�vњc�b'my��[�L������D��!�����j�g%/v[r*������ȃ�L�	mT���^�3fI9 �Ο�d���:La�!Rv25�'�w��[��O�0D��鮗����:8�@��_�Ï�'����mw�Qi�J��'�u6o�޽hB!sRH.�6e��Oi��%�c�^#�ǜ\���k�I�>�F�,��:����cF}�����aڝ��S�^^ ؤۏ���� �
����k��:�I؎��ῧ�N��z�� 6W�$1�B����k�%X�9p�nS�ybD�"کiYm���&YF��ms���EpءH:���I*����u���c�a�\s��y��w4�e��e�P+�@��6�=Tڐ!�6�w-� �ŋ�rs5^�W�>D|-�z ��G�g0�/���^�.�H��"����P��zg(���_+����x��è�Qؿ��,0ު
E��ğK�졲�}~�;gL:�z�Ol\r�V�񰋶U�� H3�NjȆ�bEt�j3W'�3Jy�\��ˏ����`��k1r��x��9l���X�[�3�CIxU�At!�*��N1XK�d@�e�2_:k~5�+�@k����3-��N=z*���ƚ,T�j�,�Q,��:'�Ꮶ{ˀfN3��ʒ�c>o�,{<}��]�q�,?��n8��+�f�wF�D��ls��[K;����k���b�<*Ȭ��'	��g��q�*Wܷ*N@��PIr=��V�����ۊH�^L�s\]��[��<��/��nវe����i�����
P����d捼�&�\�46V�D?Γ-*�ÝW`��أ�c���!q/�w��Cz��ދ��%��;N����U���2s��gA���#���^m+C[�녯S�W:����8�3�g*���#9��:	�¬��Z�6�|�@��������'o�GR��H�6��J]U�-�w}7<k��yo�(������(��"H�<d׈����{�^�ڽ�bOK�1�C#ҫ�I���w��>��["�� A�`.��{{IO����Ty�/��9,[�d�}�S�G��#by���A��&g�$�Z�rV��U�i<r��h��;+J#��[ �d-�R�Ί��ڹ�l��M�H��ԕ�Y�����k��L�����y�ܭ������@�̂��^j�F�����Uɷ��1�,�b�pН�.s�6voq=� ���W'��g6�z�l[p�h s��� .DT��mxY/Z�͆��MM�Oo�{2J���E�}���Ҝ+Bo�����^� �Hك��˖��q�]�������S�:��-<u�&:uI!g>��6alk�����4��DL5�Y�?���VF���R]	cR���8#Un���fV���̿�Q��E:/���2ŕ�!0����W�b�QI���;��4:�WH�}טr�l���QlVN��F����@�we�ޘb�qй�C�mjN9U�~�vSF*��@����([;������_;b���<`��AU�@ѕ������p>bi'�YN���8�`�۪6$�ڵT�,�V�ݘ�̥��;$�s��vQ޵��/��j9�M<z�c�O~\�*wI  ��4r�c�9� ~8���յ�t.�UT��/��ev&I̩����P�L�vF�%3�������Sn.����@��b��ٝz�+9��s��<�;;
�@L�'���M�ZKO��a�R� ��o}y�O�̞`gK~#�sk`��bOg��Be�-������XB�/߽~���D5��hlJ.�T����h��E֢ͣ&w��T��h@7=�r7�f-�G�VP��Fb�J�y�9��E����C\��&r�R���O�����p����dI�(���Ⱥ���*��+%|�����Rl��0�Ĵ[���������	����^��[��+�|/b���jחs����2��u�x��NN�+��\ڄ����_����`a#�T��i���C�,��~���Bխ���Y����F����L�4�#�v@�y��$ 
��_.2v���6��&�Taf�g^�̶^�wʋ� ���������p�*�|Y��:'ˡ��h��/uǺ�aT�eY��!��C� f�Uܻ�مI�0O�(/���Y؃����������j3����tb����Ƭ�J��M��
�ǋ��G��;�d�ln捏�%�z��hU��?������|d��(�j�Sa<ɺ�'!,��kaM�<�9&�{��}%K?�m�>��,.0kqx�<㍬L9�pc�P���u�/��nvȟ��.�>�e�g|s�;V�&浠�#�Ӛ/4w���:��K�ȏ�%0nm������I�����?ӿg���*ip�6�=U|T����!�uD��;�	 =i�j��Zo��I,�K�k�������#f)A�c����(��Hu�N$��t��fWך������(T��W3�-?h���A�,z��66'������l!6hoI�n0�R�P�r-:sr[�b�
8[�#��H?#d�=W���Rc��5�>��z�)���{	�CZiV!�j������1�G����<)��͸����R�qȌCܖ�Gcʾ�����8�<���X�7kꅕ�+xA�9M=������M@t�*"0'�A�^�Ei�kcRo��:d]ax��P�
���F�����Q����ymq�_}H"�V֞A�q��T
���=�,ڠUj��t�۰/��':�ф!��a�ї�{t3�u�5&'�jp^�Y���f���~J��w�*�[����8��o�k��=���p`-������C�%IL21�fB �|��T,�������"�if��,d�#y�[�<�f�˷Xꃌ���m�2��c���ӳ�jk���f��+�o�R�i�c�` �ƞy�Q�hSXs�9ܨ�K�^z�1�'�vT�)R��ʯ��Vf��P��<��Ȥ��2)	lՆ�p�����`�633�6_9�T��i}����%�R�����?9 ���0��ZQ��\�r�y#2iO1�?�1��H�T@����vs�ę%in7
�B�:���;PK�����[v[�8$��)�t��F�3<��+o��D���|`��j�G$�	�-�>�����݌���b�bE�%F�Z�|��)�w`�<EX�'�g�?�v���[�
����#����	�Bgv
:B�8Y7��$��U��׷\,t���}S���J��~H�*I,ߤ���6���W�&&O��l(o�c�O��,W]�4~0;;�YDToh�hd^p��.p�Y�҆���J�y%����W��P�a�cW!
{�Z��g��[�J��y�]Yu����_wsꈿ���Q[��1�E�1�*<��ԌH��ƀ+��h�#d蟲ܼ�I+D*�ݤص:�8�̭��ﱿ����"��BL�|W{&� vT:���m��HT�v^����PhcԎ�9�p���q<-�I���u�� "+}���m�gXw���V���lkW��'*X�X �zW+D��7�Ӎݒ��xO6XT��qT������i��"ge7�Q��}���(�u*�8��K������]�2�bh�9���B�]
�m����)�Ö1ϭ�	�.z��cʏ� .e�fPo� R�|���=GkP�I�r&�7Ư�",2:�d��bϙr�9��;�v,Ŧ.�R{��
Aӽ�Y9�g(Mh�o��ߌ����N�+��t�H�z��.A%tS됥��*t�������A`�+?P�F
�PskzG�i����z�y����y:����;#T���s1���7tKm$��g�~��MPxy�j��U�{����t�R��H������8toO��i�='7& ��C�BJ��T��m�+�� �AG]m�=���ȥ�*�<.6q���rE��W鎨
H�1���3���(�Ԫ���[W+�~��c<�u��Ѧ2@ڷ)S
۷Q�ZZ�>
���AJ/���:��O�Jw[X-3�wx���JZ�`s􆺜A2XK��{�2�f_�b,�LӉ%i��nʀk\����dM6��+z���ŨF�V׳�^߄�FR[4Q�Ƙ�N1��2}SZd�����C���o�Q� 1�]�$d�;" ֐Ի�+�8_| }��:'���Ms���?������J� GP���4�=H�p~���3���`pK�U,�1�i�m�9� �M�.!��Ap�-I�mA�?���J�B�1L�,��lnᖃ��8��S�������V�G����az�I���bs.�c/�uޜ	Q���9ʪ�3���2�1:�<8��6j��Ũy'��?�[��Z��O���У���KU�2_��KG
�'6��h5X��9|���\Eu�E��E�^Tu���X�䩟��<�1��~I̟yh0"H�x(����(��.��,?�X��lx̪Z	�(��o�(	ka�j��:c��K��K�Sn�#�^�$�������qDJl�t��9���P���Z)�EËV�Am��ZK(azG�E�E&���'NC���D[���:��<��Y&��K��d�������o�sԢ$I�/�>��|:������ys���XD����{��t`J��:��#	�Tj�^t��@n��͒Q3D��y�i����Iʸ�fdP1*�Pn+.�A� ~��������v�V�������n������4p��L��*Ø�RP�
D^���*��)k,µ����<8��B �m�$.��Z�/��c��:�}���\m�d\����J%��*�����i���1�͋i�h�B���R��Z�[�tej���v��T��@ۛ�{���;�ߗ5t�e̹�\�T=i�t�E �����li�&��l�z�֓!���p�=���`l1��m*�[�?��͐Żװ1C�f�=�oJS@�|�E�������HzNK;ɤ�x������Z���E�J�b��_��7�����Z�������o�%���F�_r�)w[��-��
�`||Q$��9ʶ�iH�V���������.�`!$G�W:|��B�Æ�/Ѣ�i0�Y!��K�T#Fi�#@RǨ)�B�����Ф� V�9��$:
\Ge[-�a�S#^,X��`z�%�kX?����]q�S"Z�^ �[^#�1�I����~VJ�SK���`��iTh����/��/�?ߖ������$��rj�"PU6߹$voYӧ�h�Y|@��
���K�0�w�'>��5�a��d#@�v������Q�ä~2�L�(�<"Ǥ���7W��g��]�rf�V�I���:�I R�!�3�+�o�'�#b���O"/�+�X����9��b�d7,�:W�6�"=��'��l0��Z5������Z�����F����p��tb�	������]ţ�7� $c�5�̌���0`\Z}�cP�Hv�%1��T�w>=�G�v�˕���{�������z�vs���A#���~K/6��K�;@�y���㻍������V�P�r�˖��7v��]h.�#�`�|V?��l�5/5ߒm��!P�u�͆�9�Y�W�]P�P1���4b+8����J��^kK�DKo�5El�_k02C�K��%��oyE�
�{(�0o���\�7"Q*D'���v��� �^,�w3p�16
;��SAɧȻ�ʶf���
�`A,�']MǠJ��V
7���Z�r��<�.~vՍ������(��;�����|#*'?}���V����Z�9�
AXO{/���u�f�[�I/wB���,Ze)"3Ə]���-� 3HN�����y���ZNy���8\Y̏,Q�0۳�`�^��|Ih���ܳ�Q"��C�i�������" -�JT�K]�͈�@�QveRn�F��>�pĐC��mf�ȅ9!ͽ/ڍt;v�Sܝ�񼾢��H��>#��:䆏�n8�sYjY�a��[w/*���>�y	;$cm|0^mO@AHt��z"���<��+�%U�T�?�O'���jiO�vk9�g��94��~nU)1�6����-R��)�m%��D��{�H��g�3pc v����ȁ̑&o[q�t���Q�z�E��+դ '���`	���A�KL]snʳ��}�;a!�(��S�ë�i#B��yn�l�n1��/����?,2o���Ѽc�">x:�o�tsS�\�P�,�h��,���x�֠�&Ye�=�N��2Al�N���DN�h�f#�^�H9�09a���:�oÈ p�n/��u1Z�q�� �W�ȠbTw-�]s���#ȓ/@��!Q\�0#����x�3q�����y����+.��Ã��Qu�j�>9e�K����M���as�u`�C�2�'�N�ՐC*�9�\���D����|���nY;*�qK���e��I�\��`�ީ���¡~;�A�j.�h��z��Ϧ��9n���W�����Db���0)��+������aŒ���\�I�B�h��[s��l�G)�F��2�T�0C�c7𻜷ّ�Q�U[$�¼TS2o�o��b�J�v+�~�$��#!`c4EfK0�;��(w��������}�ӎI�lLT�>��X�%�o��4_���dNyl�|� ���j �YCc���	Փ���ŝ$�q�uklî]`�F/�չN�cF����))�A�˳�wq�:5A[�d��?�z����Y�xW��P�{�gM�~r���K��2�[���#]��Z(�I����G(-sN%g���"	K�2�įv���uԀ
y��a�pI�s���,a�M�gx�O���ӏFd�=G�����+_�4mȰ��l���T,]h���&��_.?˨vU�����Ќ�O��J^"��ր�����!b� ʱS���+�&�&�y̏a���Ft1R/��)�=���1��i�)�pd�@�7a@�z���>3�w�H���ԃ,�*~�P~~�6�F��`�mq���G{���6&J5193�4O��d������wz�-45��zQ�&�����a5��V����1l�qN�X���`�0@d� �g�-P�E|
�K�OE�A�5xuTXx�ܥ��ç�����dD�^L��.��矃�B*�;#`���u�{�$�<B�
�z������fRC�u	��̐���J��fvN����5�j�������n+����Q@G8i)uK��:��=8,oj���۳��c,qp�!��U�����O�.��%s3'�C�xHҦ�~,PN���:-��M�b!1��`b�L�b��m�|3I��˷x _��F��)�ɓ��$fF����Ws�#��"[��ք4��fK>��x��~3����� h�R��	�f���qZy�BIB/rF�.�xdmY���5�Buo����Kǲ)#ꂎ�#�}�6˨x~��_�w�Ey]�AE�r��!�_�A���ԗrr��%���aA��u�Qv���(��X�B�-�h`�5��=^D��S���k8`CQl����n��c�\��V�]��P����x���U�Q	�&���n*u�T�vd��Ҟ�g����I3���wL"��D=<%���d�?���oU[L��j��ʳ&��ŋ.�$_��iR��������Y�۹)���%k�F�81�xoZa�������0��E��"'�4\J��x��3��LB���r��`�s`�D��n�U\Y�T��~���?�J1O�|�˘о;ർ�V�Aw����h�O�Nd���K�����[�8ՄV����!��0㠲����n�rk�3rf�V^I�]?0~�˕y���č��C�^;Ob���.���M�2�\y�����Q,�����2�OF��)����j�*��M��;�c�&&M�˅���k�"��PK<7�O�~��j�'Á����?"GZ�[s�.�X��'�D��/��!ϖ�٩�ç
����9U��4=��h17���PkVH���� 7���\�2-s98&�}�q>��]�eD��|dd�"��A���6V����sAX���\X=�EH���+"U���*GVoZ�;nCv&ieW'�b�q��A�f���DmoJrE�7WN�][a��/�ڴ�w ���wi�1. ƚ��l?dK�P}�W�e�Z�	������?((� ����� � ʖV�o[�)��U�4g���p��m`�M�7�C��EHL=*fd#��"�FD03'&�T��X�p���W��[�|�Ċ$f�K���H�����
gg9㢗F���V��60���T����1��Y����$�&�L��Yۢ"Y�?\��ϙd�s^Ff�Y�$�I+[1�Z�[UN� �� �Bm�LediD��#��S2�u�u�f��Ip<Ük�,h��W.<�M��������� �D���%�_�;����_�����R�c;́q�����#8�Hr��E�PO�ӱ�M���&�%�k]h?/���zLx��>��W��e���=࿝˪	z���:x�l�rߡF`��Nf���'O8,������nt ����c l��翳��,��O����������?����u����N�PT�!@������]�iF�i��c��'�m�gf�ZIzfډ[8K�K;�����p�Г�"�R��'���,߃Q�&9���:tH�	{s#yX�8�ٵ�#�㠙�fV��̓D�V~�����mc���<؏}1�*�!��BY`�-[A�\pQ���:��$-p�>�$U�\u��S�Vv�opdȯ٬Q�=4�G���d-�M���a��Ί�E�D9�w�	$ݯ�Q�]%�h�2!0�p��#`1 ��!���(�b�<�4h�8��uנc�j�Tj���@�c��H*����t�$U�z��L��n v���	e�� b��r���)}��&5k1�E5��T�J����ӈk��x�=�ɍ>��ْ�q�۟�I�bT$���Ro��,��R��_�嵵dPhvv��08��7�@��k15�����{Y�sǻ�F�d�>�<>�HxԫMjXY��y�\����\D4px�=��>p-D%��^IU��ɪ��L.r��C���(���/0.#J�*�wr4���/�щ%�<�"mw,�M�����G�S�7Q�O�RL�E����u��ރvX�����N�\���a冸���1�r=(X\Q0�XH�r�瓯�H����MŤ�+V}���ѣ��KJ�]Z�[]��L��G3�e�����r�Kv���Q0*��V�����}k��@a,���o/m��=%��v��$Rw<�N�l44�@!�}��[6������%���$��(t*��*�p$�O45=h�;������l�v���v��U��Exu{B�jT8^�o��=�tO]>����
&��l 	Խ��A
R�y��M����,�d� ��G�#����+{�_��E�&�p�v|jJ��L�����#�Ч�ǒ�A���6�����P`uT� QêJ+�x�߮��{����Fa>S/��a�$w1����'W@JhF)L�w����I��C��F��7h�}tbJ�h��/�(sW�>	!
)V�j�dV8�q�O+�+�D��9�.��p��-@�?V�����@T/��{Pjݻ����^��0H�,�|���=WL25k������q��r���Z���ID����)���Q��N�ey�ǭFi��yD�f�0{�4�^I[��Fz���.���G�_�����\�$���ʔ3֖��B�#gl�ǿ�~o���@p��t���o� ����s{P�}9�{��� (�6������>���qb�����}���]Q	@7Q�k���¨�ѳr�o�*"g)��g���H)�!��ShU��SoK �����,����t$ݭ3j��ãM�����{:�yŏD��ϼQm�V6�5@r�-����ID�~`!�P�R���ߞ�_�`[�W�h��[�Ԁ�Y2�=%d�/��%�Fs��i�T,�B�9oV*\f���B�E���F���7|��Ȝ��a�0���\��92��<��{7S���<Tj�8�R�h0�z��^\��Z�hLW.K^a���]��j��[�0������������Ș�TL)�����\'�eó��ゆT�C?�@�V�� >��6�w	�gI��r�NT��(�>;�Xfeo�Tx�/VB;���	��u�K)m����X��h�����x�4�cW���5N��Xnm��ZG=ti�|�$������Y����	Ke��u�_ӈx><$_��8/
�n�Y$��M���)π�esՕt��P���'ma��/Z���	Y��0��ޫ��:�h_��#Q�B��o^r�o�C��ϯ߅�t�@�����>+̩2���j!�f�����X��-7�r�'�AZk:Orq*��b�T2U���Ы�.��hjƞ���U�;$�6���GN1��t���v��R<���;y׃j7錘���q8���x�v3^��0� ΰ]���.>��5���o@$+���<&�5A��m=߭��o���Tv$�eL2k��C7z�B}k�����1?cno�[�_{�������$αŤ�n���tc� i�[��$����`!is�b�����]̇�j�;��(�����g�j��=��S�^5ƪ]A*�6'l�:��RxH��z��6�s͔�%�isi
�Z)1^���;�M;��Q�et|H]/m��Ɓ�Ova"+������r����x���C_o�z�e`�	}HO���]��ɋ�g�$T��[�h��H:W�ˣ]��͙��ie��d�]��6�4V�����.���i�[�Et_ǽ��.���k�$~|n���������	��L�v1��'o�h�n�?q���,hy^ɨ/d:�v�l4iHp󣼥捘_�xT�X� י�\6`Ӝ�W�%�AN�'���ʓ�>c,.(.���V���Z�����UO�Rσ��L���MP�q�z��D���c�+S�v���o��	�:F�����������a��Ǩ5����~n���0^��ML�mS���4��,O������pf����!j�,p�7ӄ� -������-Oh �a5��|�E��K�t���{�W���e�JZ\�+��m� �N���x��Gȩ��]����g\���CXǩQ����H�6�7�%H*����"�������϶�mZy�>I��|1Y6+6��8�T����`Ŕ�fr@����<�q���Ы��5
�n��1ũJ��I}PȺ�~nl
k�1l,�6�/�-�;��i��2<�����	��l���>�_W߫�S#�,��K�q�i���gkP�	�mMo	�*F��$�	9Ï[���������8l�L�Ci�il�&)�i�	�b4��M���ŷN��}p�6������$	��_.����"�s%�ƪ�Q���@Gm��A=�װQ�A䚧����&�y��;��&uq�s���*�������5����*�k-�s�����4s�,�SV)����X���l8Z?Σ�ݖ9h�N��*�f-��:��� XL�=��I�dk�Nx�ê����0ӑFos��p�i���MF��H�_*�<����n3W�v�T�	���D���{���� ��@��p3'aF�XoE��#��4 )���Œ[*Y�ğC{����������7N[ �
;W�򇵌2!�r��_��K��Q<���p�th�ʨ��s���c2�[	q���������G�L�Q}�a� ���.<�O�Sw����^W��4u� Y����A-�Wc��6^�\A�d'r��E�,�%zJ;��rPH|=ȀB3��W��׹�t� �ʕɭ#�ȧR����@��H�ۈ�EAQ���}g6~~��[	���;V�f�q��^ �,S9̷�ʍ	�Oy���{���S!	�v��NL�r&�tS}����)�Z���@����SK��L>��;�L?���+A�["��''�p,�},����lu'�FBj��
�z���6[�s{��t.hC7WZWiWԂ)3�\#���o�J�}/-cz�3����!x>��7�';�FsV�`Ds��ا�;����:K���ೠn9��΋,�rm��j���5����ET�Q=q/NM���<�b �:ߧ�g�k��%�v w��gaNZ�h�e�Q�~�y��_PZ�O��Db6��*���K,��	^�Q���cz�)��kӊh����>�}���2'4>1P6��񨳎T����> �6���W�-ݭ�,�I�'��a�$���i2τm�l�77�̨̼�w0Ѵ	s�3��j�l*� p����Y�*�D6��<�?l3=I�r�l���qHU0���	���ݜ�]<���຀Pٹ�ه(�~���r��Ǉ��Z��̀����y������dS�p*�uj�Y����jd�ۚ�w��{v�{�g�fp� 7s��\����Q�*Z|0�\ҧ�1��Y�u|�o���i��[�o�@�4E�u��q|��r)~�m���!yt�e5j.=gG	\w̹�ሾ�!����JVp�y��U�H���и�����{�o,��[yŻ�F�:��,ġq�)�v=�%q���|��5�P��M/�| �ޜ���G�Q~N=p�Cϋ�q��I�
��,�s�{m_A&��e��@���.DJ��g� P�:&������F��/<V�䝸�x���K�:�m�|��]�Ÿs^l·�S`㇝��ݶ3�T������@n��簾�Z���TF%������L��Srƹ�;Vu����1<�ö�NE�!#�?~'eF<��q� ����_�V^�N������=�t����̺גе;�+�9Qț���j ( ���U���/8;Z�
��zU�$R��?A���:���A����$?1�e�З���6�N�ΟÔE$�5k�^>�zt:k�U�O���$�ܮ�uU��S����
9��_56)%�H��>�KǆU(-
���Or��`��hXL2�Lr��c�{_�PL-��K�@��/Ulҝy���Etl��q��u�t�W��h�X�K><�^]%�ý��ۢj{^�������1�7�jŭ��[zzv�o�S⤌�c����J�f�}�O����b$B�Qn�̂GQ������h�bJ����y��#*�����+	 z@�T=��7� ��������$C�aN�}k���h�.VD(���X���ޕ;;��rE֔�Q�0x�&~�Z�M}J$�7��?Fƻ #�Be�X��M�q7r[$M��E 
�|�FϿ.�i��̥�����f	�t� ��Ox��@_�n0;��Tr����eV��<����{5��Ț�ݲ =(������h6LR�WK�W#����q��l��ތ�#��+�D7��`I��9�R��/ �������H[(rx}]��I��,T��J��+����2��WD�̈\�7FX�^d��p)f����I�l�g\ă�����SQc�N'K����μ���yY~7�1���5���w�i*pC1[�A��C1���a�K���B��iq��S�ߖ<��+<�:hqՙ��J\҅��I�ʶ����z�C�q�����0H|�_ze�c�l�F�ؐ ��6�ִ�;��*��㗅�c)������E1�Y�\�����%>ؚ�30�J���(�It�8���ȴ�@�O�f�ǳ�ܕrz��g�"�F�2"���g�q��fL�z�b��\|�-�I���]r�<��P�n�p���Pk��B(�vO& ���,_Vݷ⅜����[���)CF�������3�|ލa��V�����8_gjQJ=E��9e�4u/]H�	ف�����b��0Qyx��N���l=�U*Bܸ����A����3�@�*K�pǌ��5�9�/��u�e���������nA�砵c��
�C?���t��[���#�(Ý��+��\���H2>	\��@6�%t��� ͓m�x�\�C�_�lϤ���=%�Ψt�ZV�y`?�ld�\��S]B7;Plj><w�p�a��ָ�(�5n�{��p��KG;mS��ʒ��˒0�t����5,�͘gx�E`�rF���E�@�=���ᢗ�H�X ժ�h TB��:/��
D^`�n�V1+�������E�P��WAܛ2�ׯ�V%aJ��x}��G@+fr��F��uO�Z��o��ďvi�|Ƴ����=��F]�1���,W�@^g�4�1���bD����h;j���Z���V�R;�
5�M��&�6E���a���|�<#�eC\��6�@m?������93�&f��W���f��Q�>�.���IL��3���w��.V��R�CDa��H�0����VN �[�5'������GW$���a����k��]�'�	h}r�.��ޫ�3m^�a�z�Ԙ�����3i�dx����9M���*2#pS\b���~�mBn �a<��ڜ�&�!�
��t7=� �'�2��}	`9L�G�ɓmp�Z�$n�D��!|�!x��d����VCi�Tz�y�&�v��"�
A�&�Vsn!ؙ>��{�E( 4�!� ���%IK�>k����V��
�UӕE�������P$��N��8d�`�:�6�!�+ወO,{��Hð��~!�\�7�Iv}b���;����٭ˬ}��ͽ��u�9�7�E�2F:�NmJ�!YΤ/�����K���^yyþ�A�6�;�
>�Cn�|�Յֶ��xWl^e�ߧW(A�Y��& �[��#49v�7���:��5��wc �(0i����<��_��M���
i��_^w�S�My:��@*��}p#]ɮN+V��yx\v���� U��'@S���k5I('$yVٛ���G�NO��q�8#'��]u!��dp�F��$�p7E�^w?����KN/b��x��N��1�g������{^1�O)�0��9��d
���!<�R@Y�x��U5Y�2nkgPL4�S�Ҧ�Z"��E���),�W�)3Y'Ҿ���t�fG��$K�(��+qH���I�C�?����f:<�#e�Ĵ��O��K��]��z�Nh:�6D0�=T�i���b�CƦu��XGo؅����(���Xr�#���z�fo�ƫ��2����-�[J� �ۘ���鹎�X����\}�?����]pl&2��� ��%�<Ds0�d�W���!���,}����`}�k41�Ln��/��I��T�)c�;ǝ{� ����ɘb�Q��t������a�s��@�	ρr{��zX]e�?��4K������F�p��N=D���1���~8'�	��i�8�([�0#�#�%��L�TQ;����m�rwԂ��ƛ�ʇ^뮖+����C��6����&'!�E��h�'�l;�@-�)u����[�QE����)���uW��`�z[�c*��Y)�%Eڻbn��BHI��j5�������lf�)~�_p�S�s�mAW��R��z��ߟ��i��K"0�#gE@�����7v`��>�meҏ���5=H�^Ҡq�
n����	I碭��%U�X����+��[�����h��{��v� V�,%!���x\���/�?���x����˚a=�=b��L<i��.�Mm��|�dg���u���?؅6.�7�ΐg��(��O�-�O��i&��ﵰ�0��y�!���l��� �P�_@��\�;:�|��/����dR�fԣ=������$Y
(���re��x`��S��!f���O%��7��5��H\}��P�M��S`L�X�dX:!k�n�(s�tmӽQ;0Ix#Z��P�T�v�܅ �Ǯz�GQ�[��f���ٺ���e8t	U����Nq9�VR�n)/��������-Pl0g#��wI<����c��c�W#^):� ��A��o�)�jݦnE���s�pЕ��3Q�3X,v�
U��l����ȴ݇Z��~4K���=Â�t�;;�[�UFr1n�(�|���Um�b`S���j=�`!2�����:Y�`IM��kW#_����'1���=�ko>��PƦ�`�dS���|�+�9-7j�M&����� 1�?���m�e�Œ3��=BŔ�ޔ�3���".Q]!ƭ�)؝Hi3��{��=�CxRG_$�iL��MCɱ,dH�`��c��ͬ2r���t�&����&I��ˈG�2��l��'/i�2��rr�l;T<Y��~���~��WX%Xq"�x�W�+��Y���G�`���˚L�]����\��օ��Au�;�IU�69N������O�:M0��Ȟ�9�)��o�A0�� �՜S��� ��lߊ �	aR"�4m&�M�˝jtH�;���΅u���xd�ⷺo��\-z���Y8w{�E�6���9��ⷚ�<sNį���i���P(��O���y�݂��$�]-�fخ�����cO��x��ي�"���m&0b�;WFy�P��~����fg�)��h��=Vb�BJ?��<�� ���ZXܹ�
��ǻ�cY���_��K���tM�:V/*H��^�V�o��cL�xX��}!�jM�!��缛
��3�pT�
W7N�)/wh��еt
w�i�3����泯G�e����P�q>zޑ��e��;$�{Ec��^q���Y�8�N���s�{LfɵO)���q{�d�(b�r(�ϜK��Tj8Dy�SRJQ9x�@�\����)Xe��E�<�oH�R���va�[C�g�Pu�y.=]f�f����j�-�UI��
��2\��@��<ͻB��.#���F�;���)��y{�k[~X'-`2vg�u�k
��`h���ՓJ��c�Zr����Ug�l"{�a!'b
Ӧ���:<p-�yau��I��^�%�Z�Sc�	ym�B�6��a�B��T�\F|k���\�o�xs��|