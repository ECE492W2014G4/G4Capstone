��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|��&���i} Ĳ?����D	m\;���k��o���W�c�$'�sĒ&�� ��Kt)��A9z=!� ͵r�hQ|�{�9G0�&��o����ų5�غ��6H�T��~��QOI����b�� ���k1�|^�fD yέ�L+�U
�����>�D@��?�<W�
$�1넙����"�U�I���<���s�;���E���WW�	�o@J�a�.�\v��j��vY� ��54���6d?7ַ���YH���atZwo��y�/>�E����uQ�f�}smD�N3��?�N�A�x�Q:BP�3�&����ս�"��Oi�K������.X,i̥]�>K�����V�P{��-S�E9a
�B�N7�ۇeT�rt�.�u�8��D�[6�.�9�����3,|�MUJe�D^��H�w�N뫝q{��bh�t�9`Fu�S4� O� ��ab:j�u�^�.l8���� ӗ�s0[B-��I�J��mV�����5+����n-"��������p�I���~�ܠZ8�A/�'�uy��S�,}�En��<�*{g�!�04�v��A����M����t��ye�g�b>�w4�����;��<~:@ ֢�8[)�8z�t�Z��j�oz̈�6�Y6�*s9Z��ٜk������������7*��W�n�հ�X;W3mon�E]^[�����Tz�@P��S| ��7z��*�2 ���`½�|���QD�أkܲ`N�wVb��C��W����CLTg�X�w�$�vL������g�I�v��&4�}�2?�;��L�50X?�8��_���p��O��x�%̕��:�`[�"A����$l��c��0���COz�ީ�C�R5�s
St{YmZ.4C�t$�����T�i�;h��<���2�U�rИ���G%	׹���&AĶ?̌��V�N�S;f*T8�k�0��x�u��,V���^`K^$��O4��`.
������qt"zB��/v7n� Ј6n�ջ[��B�V7�񷇨�m�k\Ky`���y73'_��LWk�%ss����_��,J�;�"�4ɀ��[D?7� E��U��O��m��80#���(���_hw��u��rs�Jc%��F��Md���j��WX�F.�I$�q����N�����h�8�(Q"�fɅ4�^�Z��w�+2r���Ѹ���]���L�S��~�Q�@Os���8u��OV'V��H�r�@�͎��?� ��7g09�Br&s1ZO��кb�,�Rw��vTVT�Jwi§�p��d�Q)�㠐J �Ь�d̿2¿6�����&8�u
��ykRz�~2�&�6�������h<�[Y?�<M�,�|�5��g��V(ʑ�c$�X�����0Bm ��|6N��� 3�̒	�ni9��S��ev�~;?�,�Y��ab"hq+�ܒ���%1���Y=0��e�]����l֑}��7	-���[�ĩ4��\�z�Pv�M(pD�	����x0���g�?��IV0�A�STt_�#�H85�[僟�$�_OwU�y�W�3_�b��/�� �q�0�U{����{��A*��r����aD��zX�KKe��A���84"q�2��1 �9)D�ٞ�.N�:6��1��f�g⮬��.�Xw�}j�:y�8��B�C���lZhkbS�[��!����鼧�R�Ty�.�gm�p*B�{������Y�����C9�'D�!����Яԗ���v���9?&��J�W����X��}��r	�=�n=��w�o�N��J^�E�`�[��p6���I,/B�Fb��?j%{���C�@S��Z©���4�>�V{�	F|t�����ʱ�� h�z�U���׾��쾸�d�s�]b?S�xp��K�A�3��!�YO/F�`�Y�Tz��@E%�J�g,�Cmn�|ӧ6褖���;/�H�	�9�a��
���>�g8��O���ܳA}t���M�ǎ\�v�ʜ�s������<���Jm��/�5ט2��:#�� �^�t��R�"�,�fĳ����7
���E��3���¥���z6�Yj�-�W�������<�(�4W�e��6s�u���m�J�S�HY��uPB{F�'Í��������U�g�C���V2T�tK#G�q�z�h���,l<�Q(Q��)��!��𞞹���\��F��,HpKg]fҡP���}�8J�@�S�ߵ���m-�<\����J�0�ڸӒf����%=�
���OD�{j��i�E��L�i� ��1=�zO���h�]{a�ǌ��H��2��B?���%�%�wr�f�S�u�%��2[qP���=�n�к�����Ż�u�2��b�![a���Jɧ�]�����5K;u.o�(<(�P��J=���]J���hү�����c�ɂ�y��J蓦m�զ���a��Rxwoq���f�'׬�Db*�٠:�Dmk����Rp���x�)����[A�u��"Ozb �$�O7�m/�&k�iHԛ�aȇ�s	�h*�"d�$�@?����LCYQ�<�;~W?qt�Ʒ�>��C�1b4K�n�f�Y������I�s�t_���a�� �Z�8Q�$��<�UvP4�?88�����^��qf����U���q*Kc$Z���I����þ����w�cʲ� \=vC�E3�Ѩ��!C� 7�%QNՌ�n����%��v*�� ��BR%ze�bP\��d԰�O���8�Ni��s���;�<P�nt��^�L���㎊�C�~x�46Ѭ�}���K�7̘y;�<��0��!�0Ѡ%;eJ�c�~Ĝ�	��[I�ϼ�Q���Ğ6�!��X�oC�;n`*Q��( O�YU"��8���,N�ؚ�T�p�J�.��I�C`���#�P/L��0�3�Tl�:��iN?��������Pز�Ix>r�\z�l@,ތ��?:Qi���Ge]��D�^5W�纥�y��HC=B~�6����zQ�'��l�@���s:|��9�rh������5�����L%⛲�s�R�bN���׆&ld$�b�C[��u'Ў#�LB�D�_��Wњ>�a����r���+
�Q驓f��<��̀͡��,�4�����Q'���-ޠ��iU�(oV1��u���i��LѮ���=|�
��}^FЧ����)8��`������/75@VxU�
��3@�D��o~���C�<f�[<2�ƙK���1�c��F����>�t�x&�!���y_�b"4	v���Z��߾�E[��/�[�}��_�ߙ9��b9(I>pAׯ��C�v2����t0QC
�9��a_�9f�_j�!L���ԬȞ"㠂� �2c����(�l�H��E���K�A�$*D���?�l�oX����d��¤V9�A`�U����:c��r���pQD� ���n�b������>	�M6(4�k}��	)p�[<I��Ptr����y,"(��h��<�w�S�T��{��
�i�-*@��b��%���cr�q�o(n�+��p�j%�Ƚ���y. #�,ߵ��H�F�N��Z�\[��}uյ�b;��(XW�v�~�Ȼ�\5n/5� �y�C��3o!��A��fW�z�@��]���������ms�9���'1-��Z�7��y^l-46c5"�A�L`�WMx��v폣Z6%����:�U+;�m�16��ħ����ǳ�)����H_^�
��·3���O�=D\�[t��}*�gf7a�z#�NA����
�x�+d���{_�=�r����F��ʱ�2�d�fN��m{N��BS��A�&�7GVJ+w��G��H��G3Ɖ��w9��t�KHyC������I1�H���(p�(�3�c޺�7F
8���/y��"�E��1��T*"���r�Dr�cc@Иh$uB2��U֌D�}��7�	ƃ_���ö��Xw�������Oo4+.Ļodp%Qc�x���'���(hH�ɚ�iDy
�P�6.F�̥�R� '��Ӛ���lh��d��7�L�qoo���������L��||[�>hEW�o*�������������h�I)�'�)�O�O ����xT�qn܍[|�9�E��y5C��Zյ��!������@���i4�m�x��h�94@�9�>�B��)}�>
��I�{�%�ύFn7W�t�)2du��$FMH'�G�.�e��jA������N��P��1�r����	_����x��f�A�f�ě��� ,_E��h�f�]a~�h_�xX�����LK;F+�L�>.<�,]EL�eVe5M����.�W��[;���8����F�K_v, 	ٝ�Ÿ,J�����:�r<ǹnC1T3��x�Ј��e_�(߲[Y9�5?:� 쪲Gkq��������7̢!R�|�L�/��.1�ɖ��g�鳃��H��|6�.��M22(�1x�df
���o��$�M8z�$�=��U��Hή��rk.j��8��K� ӂ
T] 1����S �RD���p��U �s8_L��DƑ
,<���|�]h��8�p�ǂѡ�"��ݯ	b�2�����c.h���b��]�ت��u)O��+��R����LbN���n��h=1�3)�JU����fm�l!�w;9�D�bV��}��-�%�@;�0t��R��c����DY�:��?Ըkʗ�(���1�e��H|���s�I�/!L���?�_d���6R`����ͮ$����� �v�۰:D��f���B6�s� )���q"�O-ZT�DOT����q�<��˂G�-��Y鱂�G$[.K�����-�)Ա��t��y:��\��:x����>�)�G�K��	����HcV(��S��R��M
&h��5��s�Z��х#����>Q��(�_��	<;��Q�~�� d5��R�Gn�G�x1�#I�9w�G(TZ�G����Z�� �
��Ul^5�70���~`�Q���zH=Z�w~v����j�2Rb��� Qݮ�x��Y	 �>�@yJ�e�E�j���|�N.�$��T�#f�u�E�Kg�+bRW�����4�^3Ơ�{��D9��숌�%�Q�����ƋvV�Ҏx��U��d���:kT5 5>?��b�nb���.�pv��"��U�h���+Dt텧s��B��)>K��ι�R�7���m���5������"|'4�O @��  i�^\`����@� ������s���E\�'6�F�{ ;dqI���o�ߙ�����^fp����˿���U=�����6;�/�����%>�fދ= ש_���8^L-�(�1�����U�E��s�)��	��%0y��%���u�nK��nupx�Ԟ��������jrX�9P"���}ߓ A�"q�wY�~�>ΰ_�1�;:޺;5]��@T#�n�ʷ�T`�*1��/$�M�]�����\�i;Al���;��-�$G�qJ���m�϶h@W�u�g�<
���{P�U
��[�P�Bb��NB�np��O�;�QL#'�_IA1�xx2�:�.H��ϗ,���>0�PL�N�]:�}�}��W`�@� �t}�[����z�ۀ��Y��)�W�!;���;斮�D��(��Ҏ�g� B��*s���@O8�"���BR�/M�dZGJ�X�݃�K�FD������}��b�2�d)=,���=����P�war�e���� �. �|4�-c�'f=aq5C�4|X��`9b$j�Y�VSdJy3��F��!�E 0mN����u���k����䓙B`Us��z8�ܠ-�J7�3�U�Z����+�_Z��A��Mi�����`��Ko!�B�WF��̚��7W��K����;�	�|/p>��򔛷���Lx�����~<�m6����P����DeL��[!�4正���C�S�%��R�d!�t�+k�zs�b���*,�a�P�n}���Z��3:�08#*3����\R��
j��8�Y�*k֪�jN;bą�o��[P��V�𓞸�_�S.�b����D~Ȗ���9"q5-���vi�On��B�d��Ɋ4��<	����.�5/b�pa�J�@^<?	(��$<��	e'uS�L~F�a��1'@0Ov�37*=C$�ig���~�q�(��uo~<�el��QEX���+?,�ͭ����;6�ưP���P~���� ��w�c���TJ	Rv�?ٓ�>tQ*J��$�@T[*BI�;�_�j��<�ۺz��1h<�W��c���_�W��Q�s�ln��kL��8��x8ŌH�3AS6��QbW	^ş�%�`�{�Ǿ'�}\��r�s��f��������,�Ɉ�$g�eUn�?_��?|i�P�NqI�׸� heڣ���RN{�
�v��G}0&<����=�Xp�VG��v���#Oz�#N�?�0������+k��@��ޡ5Ӑ�hx�Ι!�L)m}nu.�y�B�H����ѐ6Σ�D�|���:�x��(�j��wMh>��� n4���f���֗��{�����R �$��Y��cz��jH��|Fsn�Yij��j�r(tQ�����b:l0^*zJ.��^m[+���|�����C�/�e���4
�Y�ۡ	^ :�l"nm�AGW��.�a��l�7�1��#�eF�|Ii��yΊ&@��p�`���t��]��oj-%L��c|���*C�m���"�"��5S1��6w�ݒ�����yF"6z.��A*��t���Kg��2��$0Y]�9�G|�H��:�y�yL�����H�>�(<#�+�j��D��}�&֚^�òpB3�6�Q�D�a�p�����U���Wt�);�Q���M"9���L�'֜�I�H�r��O�k�j*��)��>�=w�y���"ߏ��u�3R~�;e��j�� u��
����T?�������\25 .+�"g���w{��4�F��zUC�Ѱ�E�3<�-2r�~D�j6>q����tGU�����r;a����:F7	�#�������"����'ܮ�HA�x��������\�tӴD�2���-lNF�d#i�P�,V�cCLA�ʴ~Ҝ��rB')B�H����Za�� �{45h�}�`m"!���1��޺#���H� �����{8�C~]���Ề�ZΑ6G�c&a�d�hT��o]��Ž���F�r��� ^���
O_)'T�҈�z�¹~�@Ē)��Q�f���&e�wk���B � �ݖ�7�q��/�V���O*/r��S|�wWG�~>1���?վ�H+��#��D�f�������
F�m�7���8�~�<Y":[�nv�yJgԖ*��5��CJ���v���vV���#z�cR���LW�QG �-E�{�M-�~;� ����l�f��H�R�6� 3���'a��+p�?�݌�.&�1q�"�KZ����~>z�:����⭥>x����.tU�������\R�)�^9�3����Nh���<�'7�<������aLH|���](���H3�W~ _�Z�la����k[aC����G�U��P'�D|v���/R�q>��I\��PQ��jJ�Q�8%?�]�r�aS�Ɠ�.I�҇q!��q���i�)����@�;�,�@?f{m�<ˌ�~�j�?O�窳k���T^�upܓ_�;ŵ�l.݄&������|��%�j;���Yg����%�{���t���/2�rJ�r����>�Sh���xm�+-�0�=�9�:�����
���̎��/���-j��B�cb\��n�ZsGf�`Z�p��C��b�\�\mk�D���72#H��p�O�r�� q�6ڿ}
U�TH�ī���k.�N��!�J�oְ�R^u��[m��ޱU�4-�Z��FN�x���{ni�{���8K=���� ���ot��+R�r�}.��|�}�a_j��jT8w�-�C
M���V�F�A��h�}0�c�^M�<	*����s�(�4�S��1�E:����S��zZ�&�X�ye&�� ��t�>���$(�te�y��mN��:g��ͅ���A�ѳ��G$��v}u��]"��v�GϚ��~:Z�{��W;pg������:ۯ-K�d�7��1R��R� �%������p
��jlL�}9������s�!�v���Mꎩ.N��'�8ƻca�m���(������_hkb�r����4LFZ�����X��<��s�)z%h)�]�*��u��;�HB�u3���t^�AZ�ֽp�7��-:�x��#���]Ќ�(�����B��!��U)��v�"�0�u`��Q�/9���&<���7gb?��yS�gf�V����9q���ɦ��n܄���
!=b��F�@�R��\�a�;���X�XW(��c���154��¾!o���h���НE��{$]�����D��&�d�aO��#�d0���U�WUܙ_/���c�.���D'{n���"��.a��؀�uJU�o�'.R�/et�Q1�j#�n�ߺ�D�kDw|�Uޮ���֨�<Vp�6"sv_��������^�a�UЬ����E��e�w_DQ:Dcob��<FP#��s�r���zE��D�H}c�7. �)�ώ1��7V����QA�A�����#2��/	<9鹍*�}��y�vTG9ߋ���WD�1
_�f��+A�N���4�#WvB�KA� ��!���Q{$Eu���ml�y�O�� ��TЧ��cJ���5lMH!p�oi�"K	:�?-�N�9D�W����S��uiz��T�>�!xB_��"�q	M0pkJz	=u�8���dE�Y�R!��F�]r�n 	Dx7B��G
c�3 Cj-�$��ʳ����gI��|��%Ԩ��'> �_Lߨڽ���ξ0bs��L��@�=`C��9�O)'nU|�1~�[B�B3��#�,�E�C���%��qg]��p'��9K�U�߂�؊t��ת?׀t�w��N���`�3ѫ����<aa:
27SE�0��h��81gSw[sϢ��U���O�3�C���ىdV�0�q��^h��@*�9�޷����B9Ma�Y�.:�'�8������Z�'"w^�r�*��t�`1rִ6�9pj�����5�Ec�o���C�6Lj_��b���d�Sѯ^*r_�7'��u� �����5L2�����V�\��1@ؾ�-���K9�MJ��Z���B�`Q���J�/�d�������͌���Ӄ��w�{��V�1{1P�?��f�
I2��t
����w0���K)��ŚNv$�ˣ�6� ��p���A��>`�8(`0�5#4��ž^�r)E����e�݊V%������aD�Rr�nۨ`z"*(R��*ӭ�垺��X�s/��,�UW�"��5|Zt嵶0�J`��f���Pm�����a��h�Mq��3�;���x>}̙?X7�x��r�Cg7�=8�+=Ѥ�`L���0�Ŏ}�К�`�qu%�_&���7{í��D5��8��Q�J6��M{x;&~j�$UO�������-�� FE�������F�$i������a���O������n��;����i3`�(\���M�}��I7t�vT��\�T)V��k��$�`m�q}ݕ m$��}0ZcD0q�e��3}�.�jz��h��24�/%Vx��ᳰ!*�r�����T))����4���
�B�ˇ����Y�Y>��������6���Kǳ����ú�J"��hվ�_|_SҫGF+!�8o�d��=Z������ۤu�Ɉn}��=nʲ���~_�$���M�r�G[�C/�s��\���lk(���CH���+���xud����.�\��js�l7�q�g��G��x-0ۉ�ǟl#�M4
����/^�h��*,/���@pw�Z����Gw#��v\ⴚ��x2ʩ~Q� ���uAO8$f��e�4wǓX%EA*�|�D1!��H0[Uԛ;M��p���xW�g��� �+�o�^�S�-g賞� �Jj����͖a}���{��!~�7�X�=6�Ў�K�0�Z�
2qk��G(����L�]Nb�	����р�=`�f��y˪��-!hqs8J�iH}5�|Ƞ��� 2.��q#��B=��Y��0~�B2T��/�7�(4~{���lK���c(������/�i��>���yBII���0�����R���/)4��&#U6�!�=Z�X4�����+}NQ�i k 4�x=\F{��%D.d������_��z��l��P��G�i�"}S�|5`�����(��Ѭk#�Ţ�Y�^��X��A�lS�ߐmmK��>^)���,��y�� ���u�坣��8��zX��Ji�>=8�C�$ŋtG���d=zC��Fu��i���֔�9z�O��L+R(����c��%CFX�b�٨=cW�p7�ٟ��b��y�-��.o������C��qB�a�1�Q�,�uV�dym�9���x�:�}`�N�怈��fXZ�F+"zt)n����p+OG�����	r���P��z�5�	z�ދ�8��!�Kj�x�<#�u�@��,C&nl�v�r�`1�y�L�5�C��?���:�S����w�F�9Lߣ�L�=C"MDݎI�G�(ߴ�����w�ů`�i*d���Q;�g�[}J��Oy|�o���Dufz&�k�Y&SvX��\%[��C����L����1��� I�� (�_]��W?�3_IXn�>�\���<�5lN���Զ4�wƧ����.o�MU`q�$Q�̡�}6cT��C}����]G���A��LA���w�N�S��5�1�H�ES��w���>�ubyaIx����$_��jJ���(�2��v�SCG�6��a���[���������Uܞ@���5�:%���L  ���"�M�_	.g�Ku���1y�Q�,�/����~�*��O۬�CI��q��-!oZQv��U�i U�`�RTy����.���}ϒα��Y�{�_����pz�I��^���/�4�n!�m��`]��DFӳ��B�����9�Dk��'65��8��yq��O���y�_�����	D����M3���	���{2#�K�#��m���u���6�%+݅����uǿ�ޔ�6sn�-�~���$sA�j�?�CR�e�m����Dϗ���t-�#�ٿ۩���Z���_�(�y��j���������q���GE�#�\�#��9����Π�$]�_����
A?
 x�k/m�e�;�s���.�>Te^�� �/l{�q%�_
M�3ϓH�Xv'4��6����X�E�03`�y�Q�ں�Fp�x"+;�Է��?�2h������&	� ��Aw~y�,����0� �t+r�4��TS\���#�M��ڒ�K�}�Zq����c!ž�=O�;m$7^��L6�J�=!֍��׍�D�^���Ś&8��0FcϷ�� Nb],�ko�l[k4歱�f�t���S%��Si�WC?�jȶ1�����>�vn���S��5��k�������9��C�����6�!�����*A�f�R�q�VxW)i��U:V��v���Q��]��SM��2��G_�/�ov�q�IF�X���7�9q�g+m�NN{g��v[n�Ȉ�U<�n��a�q/��t�J��>���4��1Pz���
���W�wz����.�e�)��q�� ��op'!U��6nQm/n>���U>OD�@��lաq���n��̀P�:%�2ԡ	����x����X.�y�*��Ӄ��r\����ܻ�k��j<�ĸ�ͬt}Fw���i���AD��c{�p�.�V�k���O�3빦Fz��U1��yܰ��e]�M�����|ي�T)0U�poBk�M��&_,���R�y8YǦ�p�;�s��@���Y`����˽V ,��}7�B2?
��+��#�oS��������������ҷ{H ������ĩ9���=%��м^ܚ!���k��܅|Aj��vv�f��"WG���P��o��t�$%��C�<y����8P������������V�ĚJ�)۱�/Y������ Z��kT�jT$���D'�3Kmn������J��l��?P� �i $͑I�F�j;��;��5%�GC�q(��a#G��_�	w���F�� mK{&FPǎ�ԭ�Rp�k��jՍ9[�a���3����:�R�_��~�=����5(k��M*>(Q�k�R��n4|�T���/:�٠��Z\���[�e���z���Y�u֙Γ���{ 2lw����ue1l!�����a� ����6C�osQ���[G��_V�Y^~�9�X�x��܀;u��H,���"k�W0��ڡ'�r��7�%ť��Q�Y�:�5<�F:0�r�h��)땆dCE�ߨ=��k2)���xs��HV%/��h��-*�crР���q��_�M�1|��+CL�?IM�RqV�Ba��U�1�.��֫|S�$�d�5���_T�iP�<������[�E�S��^7��>`��G����FS�FH$��>��u��7 诋z��K���93$��(�HE%a;k�4���q�~6��� �Y	�ye�f	��[M��`1��&(O���25�v=���GG�:�a�Z��|�5[���54��C̫d���+���1�6�~�\U���&9��uck�+{ۦ��&*j��5�p��<=U|���I�k��
a�k
q�͈�k>N׋����� �ڻ��C����;�	h���*��L���CP��ep@qȨW�&��'����l*K\ ±�J��X ���j�p�#�4	�I��&���k�c�i+��OP�֥7ֿ`<��V*�@f�+��)��A��{���e��cd&DD���TT��k�|�!z˂����%�j�+_�۽"���m6�vM��+�`f�F��Y�Tkܪv_�7~Δ��*�9@ة������[!��wf�ZS�A]�Jۜ���������u�4�5a��ջ8���(s��?�e(ֈ�����+�{����F��i��2tD���M��}lR��&��zޟ�E�۴��*s�t��˘V�����o����!�=[��9kx����T:��*��o^iu�^k�;�x,|��:X��ocId�9�|ն9���`H�*�pe������h�ϽO��%(����d��a�cs�t���O�Җ�#��Q���T�����x�MD}�J�<O���{Ob���Vx$\�Ċ�����5�[���*���L�N���%��dě���`H��!�iz:cH"���m�w��e#ɕ��~d�^/��������>�Ζ��l_��N�W����1x��ϗ"\-��&��Ӣ���1F��</����K7*|��!uĶF����gX��h���Ɠ��i�I*7a��]^��p��JV����h�1�&�
l�������5Hu�r���c$�y	xre�MF7u�8���YN�FE�UDD}pƌ_po)���3��)#�U��\PSd;�̧7Tt�͵�
��h�U)�5��"�}�Dh��q]�O7��/z�_�x\R&δ�����K��y�%d�r�e�E`*ݖ��8��c�z�Yt�G��>�|���v�Ʈ�Y���z
�ͳZï�fpŸD���
�G��D?RV	 ��B<��:<	֘���`��F�Dζ����<��ڈ=�^��
[��=qB޶��D!���t�f,�E�VW.�b��U]Y�eu��1������M�p0�!�� �{�7ǅ�<�`N��0fƁDPo'3.��Wb�X�G�f�r���-�����|�mB�U���B!x���F,���e�70�T쎻���n������1n_Y��d�~9W���t;#I��)�cF�8�X?�lq��1LZP��X�!������!����`�Ŧ�������'\�=3�+T,��;�Y��B�:~��F�6�B8�?y�&y%�ޗwz�b�tu��f`�I�ㅲ����M�e-�@��]e�����c,Ɲ~��5��5��w�����""1�ع�bb�Y1G��x|%́�+�F�hG��	@�sf�?���'v� x�n'9��8�	�H���M�z��!
])�L7%���Z��5]����y���1
*[�䇜17u4���2�̶�@����FB�U ���2��;�m|�bLQ��� ���u�s�?�,ا�9S�����+pw+G<ֻ5 ��UC��QeM������M�6�vz�ybN��(V6UC��}��}+l_�
�F�����g��/Z�-����l��Z�1�7I�_���4�� 
�����ղ*�u���e���{��#��7�NÐz����&�6�vo&��F!	��]\��\-�I�d�7�43�i��t\��<���γ�GY�3U��*J�������u���qvWl�qy�}[+�.�@���Y�-=�%w⪩�S}��*L��y��9��a���o��L�]	S[���B]ϳW�s�S�q2v����|�x+%\��iD�H��n�'�@ͥ}�M �業�[��9���v?��2P HzB�����D�I���f#�f����T�e�] A��i_ɐ��[�׈��^�0����!Wp��w�u��$��s��DO�\]
.n��O@Ԫ�J�'�=���#�E-Q�Px��SC���Vw��=�/��@c�;��q�����\�	;���f�a����v�5��sL���1���ck4��}r�����!��a��6[�G�Su�1�[ॏHZ��u�[jy��zl�|�������3j�T�q�ʳ��]���|k.~�`��b-�-Xg׳���J��5j�y�h4�Z�2��:ts����� "d��u�7�GG��	�W�1$�X���R����ٔ|�ѹ2�7�� �x��xH̬�k�ym�y����h�9�*��uN}jiFͿ 5/�)�+�׊;eQ��
�P��8�ŝ�~H9��d��\�ʵ2��q�
w�-�����?g�W!�]Q��Twj�� �l�<>�d��m�)��HL�GoY5��!�Uǔ�W����?}�����.��t/�x�	D+�k��6͒f!�f���TN*'G�]|
���О�!��BG�C�����e2+�d�J�������Ez����}!����(� V���ȹ�Y��A��|\���~^���#��:J ��q�:�5�ɰ5m;q�gb�&�p�0�oU��wSޛ�)��^ @�CxY�ߩ���j����h"�0��r�.���L�[Aw<�n��]���cj%:�'���<ݙ���+I���{X�u8�g����X�s��⃋v�$T�W(� �w0 �C�e{��HA��$!w.�w��@�<��JL�RI� *�/��ξO��K����(�C�0�ѡ�B��Q<��/<�G���g�r6�.�v����kF8=$�/P,m�.��*8���� ��W��4MV���iW1i�Eo�D�,ζ㯊�b)��</����[����opX����N5�OC��,�3`�9JFj��1�=�ɗ���r$��mm��$)�Of�d������	Ό��R�w"w	R<���qq�q�)��9��<�m�B����䟆E,J�~_�Z�G��{_�{ot�ڲ[��UΊϙ��}�L�T���I>f!���>��i�lW�d�2�^w����Ah:�Sft���A�]�?�cg��hex��v�������Zz���[X�ZXN-H�#R����;d����I�HZ�F&+s�E�15mӴ�y0�I�55bh�W#(D��l{t�������ջ��p��%���s�d���f��XǱC��G����l�IX��2�!Y۫;,�bp��2�?�R�i�fVv3-F?���H:Yu��Y��/��Ž�������(�`�λ��գ��ˍ�j��r�ʛ��v�`�m�=$$� ���ִ�1E�44gB��' �֭��)�!aw�w�K�\6��h&<�L����v�!X7��mC�r��dpw�`�������[�.�&�t��nW_�]�.4���pԩ������W�y��T�㓥�C٢Xq��q�c_R���`.�w�r�
�gu��ȲA~2w�aa�\��/��d�=r:�ۂ�?b ܛ��.���F�bCG9�j�g/�c��r �f��;���7���i�⷗2"{/։$�?�+t�oE*'s=�P�^q�p�V-?{w��9�a���z��a��V��=K.�4~��^���וկ�f?�r����H���K����I;L����[Q����8��S<���IS��-�!��-��t�?�Ne�|Opx(�'�.�Ԏܓð�K#�xq{�,抙.?Ȳi\�S��?<�Xhj�X9(�ǂ�����=- 9�����W��rѝ1D�W��w=���'
lUka�M2޸�-�ɢ!�mgZXb�_;���8��{�7H�mڸl3>5���.j��|};��B�&s[L~�,rznd"�{���/̃��Ab;�%U`wJ$V_���M��|p�U��ZR>�CI|[��3�<��/�ekP��:0h%LJ�J�o�ҳ%��z�cqоck�=��9g����e�9*�	8If�u��̩�u�	;{�m��U;�Yq��ݷs�Q|B[�m�n�@Ə|YW��� �ڪ�Vٛ���A�1h�p Y�o�q��o�B����e)���T����ˎ⠠���2�y%T21c���!��@շD�R,�E�:9)�qħ ���<��tx\�!�o���+Z������b-�a�0=*�oI�?0��w/ZrI�t+���,��z�^�$���=���J�~���������4
Ts��H+T`�Y}�py��J�MS�^���aҝ����B�d�~��U6�R[3�ƫ��ؖ���n���	����x�<'5qEȝ)��7��j@S��%��zᑍYw|��4�Z>������1g�DQjXF:��uDb�7�@����l��7��ӭ���"�\����m]���{9����o�����u�*�@�?��N���xH���3��
��IU1o�_w�T�a+�B�2�x�����νJ�K����u�� �,���Y�U2���5߼b�bƛ���BkuX ��[!1l����~d� ��U�$��ȯ�E�o7��י0���|�hb��?	!E�9�ɯ.9��{ZF�^���a���:��ٹ'���	��5���S��d���U�ڒ��ޡyG�t����I�X� ��p8g��ުD�F?-�����w���iP��i8 �|����v�����/����J9N�,�G���a&��]=�.F����"�n������{\^n�=D��
BRu��2�t��CP�2�C�6^N��Bf�ח�a�wo�u�/�g���>��2�p28��a�,ˬ^�M�tD%�[���[���W���Eh���~�7������^UO][v�+�-���9ڈc�h�I�K�y0ޒS"kk<�"}мV���C6�q��P��^�(m�F��7���ዽ�"�	F�Iu#��cS".Y}Ј(�f棺:����L���_e����U�7�v �S*v#�)Cz�$.l���X���5��n�{�i랒l��dH`nŰS�|fL�3��'S:�su���z���w;�>���E�K^����3���^�d�m�X�5��֛QiF�Cc����wx+�	du�B�ߑ�Z�v�����E��"DP�e��;Aq��gs����O���u��~�r�T6��$}C�� e�}�xb�WEN$��x��u�����A&�Q��S.B��}@�[9�k�T��&��Z�*穸�_~`�1�Zwd�p8���F�T֜xh�XĽ�1�n�ܰY��\��h��	�0p?��`���Og��Wd��wjQ2��I1�v�W�!%���(�/��;����u�;-M6@)�#8ݮ᪴��\e���������+,WRĘ.EZL�v:^ �5�J�s�_�D���!����� ^JH��}�������M<�Υ/��7��
���$c�$ۭ\�i��=g!>�%� $>p�`�FQ�h�@ĥSl+ƕ���M�D������ٜ��l����&�a�Q��~��%�D��ͮ���[�)���ȉ��>����"4햱��l�)�7*��Gc%�5�=���j���\��4S��+�x7;�TbEU�T�� ���$V���u��@G�P��PG�?�ԕ�$Cg,������)OnF�<�_:���dM	���aA��3Kb�WL�7t�K�Sm�̌`^�w�����1�^`�Ꭳ-ARv��ay�ﺃ@NA�.�rQ�
w��:�{�N�*G�nG�L�\�$�j�y(�<۩����H%J�~7)^���º8]�K���r]���1ʛ<���7vU���>Z���=}v��N2�a����^��Q�`�@�,��+ω����u8���6A6 �0׬���
�OG酳#y��͒��Q�/q5�FdX4�ѵ��{?� @�w1��_�ZYl�8��,���e��t���i�幱r[V��9Q�셞1%X����y #�	�X�h�Z���u.����}E4}$c����Dt9����������{O|�k�5n�{�����sL�-���̫~ �	)2>��nfp7�$�O{Ұ�������c�:e+�:��p�S�U�˼uv�Ћ		;6k �b}��e`�ͽ�o�M4D�
�$�!�9%�U���O�U�Lu5���O�]��9��D8�L먳�[�C_��
9�X��ƴ�=���E�:,(i#ג|�'@i�)RM%N�w�����,�2������5�KO�C ��s�/���uz佝�y����kq!:LGя�D���C��H�2�Z�li<��į��u��͂K��N���: r;�k���Y�z�!4U������R�]�G8n����e������A�Ӡ�_ω��t����ԣ4��q��B>WpƟ��^C�\$$2ķq��ᆢ�ZwߚK1�-KzS�? ;2�,��!|u�Ů��lB�_�Z�������Z7�x�Z�ޥG �ջ9������\>�Cg��&J�=�֍��~��}��pݹ�&�|��o�%-b����t}_�D�@��t���]2:*�5p��?HRM�]C��n/-��M����~��0��������l�w��C���x�RsC?^6��!��1�S��~�`!	�M+`�t�Nj��k��O�*Gi�x�)=-���;̡�t�m��∄.ĭ\\�+kaS��NS��]L5�����,�1�q�K�9�眥6�ǹF�9�ap��D@�����bY�0q�`t"�c�+�к���ka�A�"ۡ����D�G
��gy�0������U�D�̭
��1�Q�~�:�X�Xo��%��Y�@�8n2�,�̶-�ÇQ94bBN˲8F��r��"gqтV|�*��:��x�⏅�B����dQ����>�h�!}�]U�P^?Ā`cLZ�o�ju5��8� ,�V91�P�'�C�!�H
3mb���ھ4��v�I"tؘ&f�I����g�.}��|fE?V-���<>a�miSW9|��]c�	z'3qK\7���Wl�8�Usn�<CYF~:�(�e�1�vlx�R��':#wa'�i��[l*x����q�CӨV���X�r�,�1CO��c��՛ ��t-� ���� �SQ����»��_�|9ç���u�S/�|���\��w����iB�!�(���4	|U��5W0���jY�W������VUnޯ��P�����%���E -������`��'�,.���N�̩��P= )d�j)���]E/q6o�3^k�S�v��'��wϣlѹ�TLr�1�� L�gB��{Ld�����d��kMs(!�h�u!V�G��M~��)4��BCy�^J����S�T��q�E]Ui�zh��)��%�|1�d�D$�w�^'���k�"�V'�>b�^s�y�2Jh�[>$�]Վb��%饮�L�
�Ƞ�dZ}��hMB���-3�3O�c!ӏ�����i�����fr�ԋ-Y���ࢵ��u\�>�+��m�\�G�~7������9���e�|��A�V�Ľ:����l2R��"/���l��U��s��Z�&��\F�`n�mS#���������0�z��11������]�1�e}$\ <3g��Lg�?����.�R:�Uī�q��8�y|��n� _^�nlEi��ւ�W��@�h�hN��ua�M�a��A�mRr��{
���?���W�X����i�G�o�8���������f�e�^���ndƘyP	�@#�'g����8�BD�DS��d��^-r��}�JP9�8�'?���:8%�YӪ����)��tn_BJ�(Xp2�T�
ϹcL
/��̅�D���`��<t>�9`-gZ&�O�G^�ͩ{܉m#_UB�3��0�<1@��|���E]ͷ�Iy�/o�=d��dC#Rdm�ّ)�
O%F�o�`�3�ߜ���6�����<BJ��cN\�cW���1�w_I��2\��?Pr1��FC�Q�V�:1�y	�����d�S�֖έs�bc��)�/�)�}MyP=�b�Tx/����(�6�����eRaB�4�O��,�r�[�a(����E ��|o]�f�H2�i�6t$� v��_U��7�	K%�_�x-n�@��:Q�w'l�����_�dr^��(��:�/��K!_W<��Tk|�\���x8b�α��?�W��M�~����Voˡ�F��[�b��4��ln?U���Pv��o5�vmB�%+4�a�U�K�s
�`�� �_��V��+I?j�LP�d�R;ٚfF�r&Q�C��]���`Bx����n�s-m�E%u��KqH��9��͔bK�Ļ��T����W��;��m���"��kP��-H�7mj��$E0�i� ,���-1�n��MqG�X�zT�b���Z�'�����.���靭��z��XAB$2M��&�w`���<����z�]���p��r�íP�6b����N���тW����%[�m�V�س���#K� ^�+n����e>Ӵ�^� C�u�B`���aө[�?��	p!u�<������������=�#U����P���8MݞF�݃l�ô[�o!n�pE	I]U���V�� ��{��v/�*{�^z[O�vkg$(:~ۤ��1�y=�=ݔf��7̀4�s��t>����쐄LA��:�Q`�e

��Df�u]��;DP�x��X
"/Y[�g7��]Zd�%�|}o�Io�S����$u���%��z�.��!�=�P���i���r� ,�XY*�	!�옐wBx�(��c�MVד�,����;����Š,L2��zi��_{��^k���ߠf�7X�˯t��YL�A�m|E5�\v�
��U�DA�����	#�	q�~M�9�F>�>A��(�#���&#S�S�9p�{�����M}sZ�~�
��hOɀ�×Sʊ��u�vFj����Z889����]�y �u��b����=��By��D�!<� �Pn?c�`6t���	��S���V>D���|�K��Dm�l�z)*O�����A��BJ�}dv~��-��/ټ#����`3������Y���ٰ��l�����p�<�J��g�o��"�˩&(�����l0�F����mɴ��I�g�3���3��)����uY�I'�5��i�`���cϐV9�3�}௿�1Ï����Gg{48 ���@u�w*�����H� �,3i�L�FeH\��[�4g�z�x��~so���튛�lQ��:��H�\�6ӄ��!�h+��'ڹ��`�F�#�����r�˻��m�t�2)����P�T�9���J��{4)o}CF�T;���R7�+D�	��T6x;�@�A���:V����Lb��o�/tcR/r�$	�����oN9��&�f�!��G�q;�*���{gr�-m�D*��6� �TP�w�d!���w��	|�I�s������F�Jˮpt��Gc�N��'�@�����^�7��/Xv���X��Ɯ���>;�tG��ۅ`wF�}�؇�P���[�:�A3T�hj��C�7��e�	^/���X��y[̅T�E��Zy$	�E�mv���]��\�J��ɑ[�{�,0?5��/9T��ω|���N�7�d��aT����ɨ��5!̘ܿ|�����m�(k:ŁC�u/��.��_	4����z���]���f��]���ڊ��1��f�n)D�UwZ�o@ܶ�mc��d_��%��Hb�����y��g�  �r��1�n�$��Ve�p��\
G���[6NU�Z�<���RÛ��%:�].��8V4�o��c��s�2ݰb����i}ʟ��rx^Q�7fSn�b1�3%��H�-�iҧ�oF��LH[5i2Q��g�5��ؔ��5x9�wfW�����5��8��@5kʙo��kjI����[�
-�S��1(���"����_C���`�XL���Eĕr�=�}ab�i�O���G�a��0��	|��U���qg�eZ�/,��W���-39�-)�8(�qv��.����r�[���@b��X�,�x�ou�|k�H���4�v?]G�:���I�_���Qj؆�u�V�B���za]Mk���㺑
����G�0��ɟ���Ho.��/�	��}�؃�Kˣ��6�����ؾ
���/��m��R�ݲ5��95t����i�-��v�x�!9$��2Ť��-��f3*JHܔmVdz�����i�ܢ��/�{��G���$'"�B����%��<�$�7�J����m��&�bY<=_�@0Lc��u�r@�^3��K�c@Bu�U��V�E���Ae��.if���h0-K�����e Q?�i�~|�ٳ�3�Xj2!�6?���'�]��.�����,�\e�A��"�ʲRƽ�ۡU��h�I�PU�s���7���a\��;�G\?kg�6��^��[��Jr� ��b��3��L�vdI�f��K����
5t)~����܃&�B������� Y�o�}��?�^r�#�Ftr�Ճl��ck9///n�C��>���˦�u�����wLsA#OW+�-Z/����e"�&D�)<PBtU���lu�[�k0�$���.�o*�
��	
$�nk�W��5�Q?7a����녈O��}S �t���Jp�2�ؗ��џ0�^�3{.˲����,;p�꾜�"�$�N�>){�=@Fpw��q>u���Ut0�(���� 1@�����Ձ� �$�$kqꭖ/�ݨ
�LiC�>��fb�8���S.f==(�NdϠ�T�'��`��[#��Y�-t}�;���@ٲ��rB�K���k�l#CBƟ��P�UTif��������sF���`�g��j��嬊����gUm*�v��c�0�]�� ��%�M]���Y=F6E5��4�i&꫑0m��o{�O
����l0�W0v�em��#<��a�ku)�(�=���n!�S2Q�N7����D�q��