��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�"��F9s�`&���a�oq���F�g�O�]�<ݲ����eCL��D���{�5��8̝DFI��Zp\m|Q��
�}�6C���UnF:<�jΈ�2�����<����sf�k��,jڙ�����2��X��Ss�HL��	�������+g?���N�Ż�����|�v7�{M��VNB
��Rs�゙�Ld\��X�'��R :�J���^�����kMkx�Q���3!P}�e���Z�Y?.�U{�RP	�)��lI{tI(S
7ZF`�ͪ��% -�� �o�☀Z�V���?�����? �8��.P�_s����_���1W�s�ߴ9o��'Z���j��
��G�I����=e�q]m��wJj�3j*�1�jgϮ��rn4�\�TRaZ��|1p�C����t�o�F'�.`1˥�tQ��$�X$3����o�K�Xi��2ˋ�~w)@8,�Gk���'"��c��4�By���=�c��gg�,2�6qa|��!W��f �=�B�2T�I!�a4�� ��yG������S��=+�L�:�d��_�d��Flጿ���Mr�X�f����W�����1<�ﵢ�v�Ԏ�O�GPd���j�0��,�c�FДg7���C�bc����RU������"�d��� :)/���� O���&�Ƞ��_�n���Y�}�s�eS4:3��%s���s����E�U��̟uڼI֤��}=�\�1|��;3t������l���j��_I:�����\�o,�n�V�in�=3vM�!cK��=))�XԊI7X�_4
�����q��swv]��jM��DS�a<�P���o/��5X�/|Y2���J޿�ϕ�,�y����(��91��g�&nB硟���
�S&RU>���6 ��Tiʈ�	m2�ݿIڏtdCk�3v<W�[��lF|��E;%�ԫ�(��5�5B1G�! $ߔSgyڌgj��T�ҷ�ß%Bq��b�j������G�$��G1�+�5$�2=�=A�N��B 14��>�۔g|��6rD�O��C���Ɋ���i�7OY8�"��ɺ��|H_�)=Y<4����B� 	���i�򰡳�"�4��~>SDKE�	9�ʠs�R���-c^s�2�e�H*��F�뉤9I�~��q���'N�w�fk+ �5R��}��r��.��? �Sc=[s\m[p�`u���D��gX+-y�j��CW�.JԄ��"M[� �D;�c;=T,ᰘ�b��h������4'��\�+ �J�P�,�šjƫo�{�495&^S��N�H0�C5�����v 6��<a�OɎWC�;!tzE��u��t7�+p��a�~-�#on�1�5���qNѽqDl|o*�`���.��ٔqح�sx�"�_T�)��,Иˌ��ّ���*D���Ԇ�f]��m�O�-j=�c3����u�F��H�������5]�A�	�-ߕOi�Dw��gS�N���	�L���R 1o#��Ř-x xw��6�o����Ȇ��ݵ/{0��K��(1<�Y��i��E
�>�_�	�m��#US�P�����-�2"i ���f�� �	�C2��{������ˍsb}`R���@���ѣ;�z�����}�������Q��L�Ö�'�P�p^ٗj��у�T����jAB ;G�������6��+�7�Q��[�rܠm��,z�x�qaUk��2a���i�P��ų�фQ�B�I�������l��s=4�����i8j<E�}��r�v�	b�ڱ���.��X�m�P*3�6�f�sU4�$�l��k ���s�;��|�:��#�g��N��i
����ҋ:�9��
�D�%Y�d���1�z���8�m�������ѕ�H������|)��$����P_<�V�!9�h�F1.bC:�r����-�o<�� ����"�O�{%��z�#�$��b�)�� ��'|����㒫J��P�0�\���>@�w^�+�\R�0,\��-��,���}e�S�/Q�&{����#XX�2���9�|"T�}��_��H6��L}����-�x��Mò��������>=k�B����֞iV�ۯ�Ai�cA�Z�4v& ���B�5���ę��o���lp���	ǖ��@e/Kӿ���-T�z$�f�ɖ-<$��NQ���Z0�Cm�u�9v�1�#[� J<%���t.@3��O{t�A!� ���t�}���3��+�Qi�)����t9�.@�V��lA��qZ�=��r���wX>��'���h�E�2�'����%?�!�q������	0Q$�T�J�����{��Qs��φ�]�~��Q3[p�셦3��+mp�~W"��9��'�������Vj��6�'�.4ik?��ֲ��uWFZ����bhh�q��^�CχP�����f&mX�@�	n�S�4�Ӯ�%��R�&G�;�MB?�^���*�n����C��Q�*�:�A�_ �!Q�V>���@��T=IL�_HoJ�v���f~���h�Z��nV>�O��rx�Z���r���;���U�'���C�S��P�D�}��r�ִ:�.�R�� .����. "�ᓚ��tß$��p��WS8b���1���g�kS/4e��}f��5V�_ A�$&>!#jͺkWOc�N����A��b�&Ń`�P*��N���w��*����Kd^�v�S��
F+��b"�Z�C���bj�@��2IǱ�v�
,�ɍ���z��T���%� |�{�b�C/���*�sq��@S�ِ���k� pF#�2ag�I
��=;}a�ܽ��ɦ��Q!��,U\�Z:���5<�>C㘥R�0P�m���
���8�0z'�%��\êa�Iy�7%�I�\�k9�@D�\�6*(����@���J�s�Y�px��R��p�k+�QA�R�ȃK��RYk}�d�p���}+�'��Ֆ�k�_*#�$����4�s��H%���b�"3K�C��k�0���Tp�7�q]>�cc�^�"gt_�踍�����"l�g_k��a��a��[*P�Z�8�W�^�R�����%��܇7��63�K���RԘm�P��}�=��(���y 5��w�N'T}E��ߺ�̱�xBXwir��ʛ���5�dY��1Eyu�t`�ɿU�L�qDj-�� x��?�8U�Ŏ����X��^o~���]DE��7�'��ߦZ�&U�pt�D�(N�X���-Y�ʫ�#�6��D��Sț�/=e��	���ICXg�-X�p�d{��e;�}l�;�oHXn�V������M<H�a�R�XS�!�]���D(�6����(ɂ&@���ǇuF������#Yl~/����FJ�r�G��u޹E��*e}��&S�ꆶCک�F�b�Ş��l���B�Y�g�Vѫ�����J@kp-(�*���
�*���\+�V	���~�>��Caؽ�c9�MGڽ&�{�RTu�Vܙc9s��0p�D ��k�� l�	U9pfN)<�5�D<_���g�ɂ�~���~�,�L��;��1V�=����s�S��a�O�#:&k���\U�������' `���� Y���5%�"+�� t������c� ����6��w�R��P�����^��8�j1�M�2UЖŬ��=�l3#��P����D7Ț�f0������L����GzZ�/�����|dO��л}�Qoio
�����C3�#�%Ga܋�-yTz@�-,��2����$Δi�>�O���d	�ײ�4�Bc&�pf����#.7��8���G#���4<���; ��Z��n�;���y��sK��n1�[�²��U���*)ݷ%��ܓ���U�5Q��4_+��yKh�!R�>Yw,������,����tܥ|f�Пo� &����d�{�^B������{	A��Vf�����_�JS��D�?�)�^���ٗ����,D��;J �p��q���t���p{�Z�n
83���_>lճ[%)���4RE����xrS��w�w��s�d�6x�ݪIA]��շ���V�գ~bD���#q�O\���}r�3�V��5V=�Z�PmX�<Um�岭�@Ix6A�!k=qU��ʻ�<Ӄ�}���ޝ�)���V��HWT�"o}^�į�2���V��Q���˛���x&�Z��t�eJ�=8�`�_��9R)H{j�w ���8YZ��{��Z�Ս A&���W-��������;inr�P���S�_� s7'hNO�v�!g�KBP`㺟�+����#��ܚ����[��	�L�q����v>s�ɶ�ߍ`CdG'7���y̾uw	��턦I�ƨ�.�P��x�p�ӂ�&װ�
yI�Om�ʳ��/�W,��9���v�U�P@5}v�΅��7uzCs9����w��w���`��c�р�#2�x毪��g��DW0ڛ�j��y��d#���)\o��s���FJ"^}�h���4��s���e|�SHpB��n����0r�'�����v��s�?��T��P�
��]>�](��@+�|#���C��$p�眆?�z�����rf7�D���L�n���A>v[/�n:���_.6�%���p�hj�⋠`��My3�#�i���Q5S���Z-0�F砥8he�v��(H3���0]���P*ײ�~qS�I��-��<v�TF�.&�e��XS�e����e\�<��U=.��QKM[kM0�5v�]@���N�q����`��%Rl
uH#�٧��@]�z�N��>7Q�g�`E�����0��WdHs�X[�Xۈ��(gh�Q�3��T-)����=7['Ww�B�j�d5ǻV#�޶|8���(X�uS��O=3���V��t�!��@O���[A���I����
rE)U.į�a].�_��v�`���I���n���!�+�*�Գ�b(ke$Z����%�0,15<���|7��m@0 qS�l  o��9S��qL�M��_�ۻ��2WO=�$�#��e��>'�q,��=&����+CT��q;����� ��V�s��C\�����6vYu��V�Z�3�����$����Y��F��*��ԻJs�]0Q��-�{.�����僅ى;[&)��z��A$����'˧INTU��� ��,���®%Ƽ�i���/ o�";o���!18`N��V�Pܣ������-��ڄ>�����i�����6�[<S�&,aˈ��߁�>�h]����ؽ�K�&LjaÆ>Ti�W�۵߻�+7��ų;�����)��g�N�U���� ��N���>	k���$��C�����Mhį(U�$"W$3X�4�3��,��;>$Ni�S�'��j�+��j�w�H�����7v8V��W�"]穼T
泶Mi�FW�ˢ���E�R3��z3�.�i��BLL\��G�eK���Fƺ���<��dئ�&�Ο^Dݫ-ifX;䅩o�r:�o�]]\����y䷰$ĥ����ws��j�Oc�q�-�qk�>�-�������[�A����w[&[	B9�͕O�΄��_۶�Sw���#�E��ھk���!:KC{�����P�J_�	U7�)}�!��I`ѱ�����?�-9G���Z�K5�D܏�O�8��?���#E�ws�ا��
(ExY�Κ.���oz$��)GQts��o+Y�J_xr���F�]���3\������z� /����0bb�XC-zc΄����0�\�lA_�H5t��M��塔��|��+.iZ�\���O֑�.�q�@>d��̩9[4�'��U�ub����5��5�����=��+ӤA��K͏O�H��P�27c='^5�7�l�����6�.g���91�w-چ1�4���hѪ�ۧ+p���H���a� ���]po���L|�,Sg�.�^����/Ȗ�V��m�<]�0@\�:eg��o�a�#��M?��H�ݻ{�
�`:����RL1�Qͥ�Y������~�T��ae�!D�RiSew����Ȏ�
|�:,���HH�M��a(�syFi��hM!��Ι���l!"�ȴ���7�5�$�h�+��(\!�$&[Iq��.|^�2�)HQ���I�ՁUKf��;8���y�
Y��mÕ����ؙ6��%v~�mB��d�
9�q�͘
���O��A�C��F1�ZYU���#�[�%�D����p�W�̍�?��ș$��r��O8OQfrU�Z�N%຿�'�&'��ʛ@�S&��ɾ����|GHH�?#�G�Y"��y���$ 8S@���*D-mLJo�	�a���K4�>�KG�4q��x��'���9P��5Ȟh9`�sQjE�zy��Z/I���&z�J�E���Q&����,�rsd��l��L&�&�C���JB��\0
I�w_r�wڒ�����S���Z�t���h���­D ���4:L��I����$/���� n����fB�!�||jp.�.��Q�V��6z�c0���/��g��:.���m��?c�W�L"&��1��)*��&��#d���3ѲlR�V��7�s�vE�[��/|�J���Ӻ>ӳc_�&�t�l����r���{��Ar'��y��Dh���Uoæ@�&GZ���o[o�7h7�1�B�C�x�x��/�4���O��R��E���n�H��b�%�L
��gՆn�n��6���lRE#�BFlV�o����⮅�P�����J����'m3 �ߺ9�3�1��!�t�C�R!�Z�>bB�k�ҭ�����^���#/����P zZE�LW2��:�H��0��Hۛ��>��p�����։h�șH˦�he.�� ��qZA7��l6�t����"#r	^��=�x�#R��3bBo5mI�z�6����ek�.C>w?������ɫ�6����>Zf�qJ$�e���<���� �u"����*�|���il����ǜ/����mN-=5yP�����H�hέM����T\g9�xT�N�_E6D*u{��s�A$ ��֥�|�y��}�Rc�D�'@2�5�M{ͯ�&Y�c����K�#$�>�@�$� �V?	���N���S\�y�yD�=���d��M���owd-+�p������$0Ľ��mi-�s�K3�ħ�� ��l^�����V��$.�S'.4���M�ŷ�.l�M��T$%��g4_H|��+I��/�������GI�L�gZ��L�hZ�ϊ��V�k�l�������M��U�U"�/V��XE���_mU �p�ze���P��P�'%��X�V��(�9G���{ޑ;�n�6)(�M�R��O+�����r����pz8�v����ݐ8�tԒ7�1,zm�X͎�����4���V]z��n�Eմky�?'��!K��e�Z�N�u�k�_TC/��?��J$�,}�nT`��/ۙN� �,�<=�������_��N�ȭO�u�@��睁S���n7���_���#,�7�������]P������V3�Σ}LW��t`��M���\1�&ZI�B,�<��̋f�*JG���\"�҅,5��:J�sۯ'ʩ�gP�>������l��x9��Tb�Qٱ��諶1��g����=*����X?%���
^�"O��n�X�I�<t$8U�=A�uuEv2�8X�y�(�������5I���@~���83�Xo)(R�qq�����F�s�[S��#�ŨU�P�'4�n����G��jI��Hﶡc3F�����}��YQ���XyФc|���Ue�3��T��@�{�HՍ��%���H�=�*N779Y��2�7��ko�1�l�Z0�����oT&1��ݳ��[���z&xT��ostd;��i�n$5��j['�2Y ~48�-�Zq`xL-��6�q�
�T����b��ԙ��E��vZ.W�����#���a�v��%���ƾ�R9@�5W��S�d|��"�k�r�@}���qĽ)��0Zj�F-�mD뮊yuǯՎ�+�}�qk�h>cw�U�����09����g��I��y�}�[�W[<
��:?Nm��_r��E63�_���� Yձ�z�V��L��jߔ�sh��~NB��4e�r�������t@{!cJ+��h�m�g7�zY]��������ua��B-Y����3�d�1R���coSYglSv
�X�Y�B�Ϡp���to��tA�{�� �&l�����n���;��}	���f>V�@ViOv�1_.@2�ؾ����5�|�~�:�2Q���4d[��r;K�*�b�S��e��+cM�AB{_'6���K3�]������ �0��-��rw%��ͣ@�b�y.#s��t��8��Y�eM;��-J���ǻ`�l'�SY��tB�th~��5��$Dx�FꩆX�,�C�L��u!V!���!�p
ʈ�'��7��<N�_���;c���+  ,Jy���(צw"tǦ�e��{�}�hn|p���B�P��|Ax򋹨%�m�d5^� {���J<�h�ζOA�+FbN�'�c�:=Ϳ9�]�QgK�@�a8�r8��)�W,s����`���Uu�8���-m�m�\ 9E�/N��m�3Ml�~�Y\�s�#s�lL�I�A̚/n�d���ݬ�38jk�
]�����AN���е���I1L����s�@����*��а�X���J�c��}�X�t�����BߕQ|[�_"�d=HBr���Ќ��;T]]'��x��"��uZ������]�Çu�u�=��T|O^�"Zf`y{�ߩ\|c��&�w�8�=���Nb��X{5�s�����zC8B-)�u�j\�7˨%jb���z��+��翑A������3�����&C��!M�A��}:�ն
5&k�8���	�4����6^%M��$Of9��~���������6��5���"�ڙc0�l�;� ,���t�.|����B��߭��f�p���l��r1[���E1 �u�#	���O�~N��D��Y�L���7ނ���f-P��DsfUJ�F{��LY�[���o�o�z��:���J"=�������vH��\������˵r2�V�	�zL��s��Ĵ�OV���^�-5��f���ty?�ּW"�9�q�������0A��{���r{�Pp8ķOQU�=�$~�q�jDyy,��#]���d
D�5&���s@6ԽG��"i�H��L��h�Lj��d�~4|�F������{�P;nMG��`�3��:��vV�J�a����w��P��f�1�ϧ���aD6O�!_ѵ���j��b%��̇ ��B�J���y� ;�,{��G�s9+B�Uq�G��[G"`�;m��w����+e�É��E�?���^��'��!�{��Wzv����B̋:����ڶQ��@9��%�x�EU�7�C�շ�<A����q?��f���7~T�>ʨ0��jbz>�R��� v|�"Z����?G��l�#�/{��?�#d"����o�,���Q������ 1��(��!���O{`�˕S����i^R~��5�ED�{x����h�>�������ZZ��R���@�ӭQ��� �-O�h7����}�9ͩ'�hhLd��|�Jb�P��zc��8�j����լ��;Z<����Dk����o�B�K��C�ho��c�OR�-�=��8�så��P�a9�{a���QȊP<�X�;�Qu�
>�j�����D�I�{w���Wѽ-4k�t�o�W����6Q��j�cёׄ>��u����p�v�A׋���;��Ȕ�F�S]1Uz�8У��*s=L��5���%x�Ҽ��7"���]J�C��"���zT%��� U�2�?D��I��>��t�qY�Zq��`\��pjޟ7D%����8��D�NC�
�#��o�91& R�JA��"�s� �RS�� �N�kpޣa�@}}F�d%w�,
�n�{���\;�6��?�E���@,EE�ȍf�2r[)}���y(P������'�NzN@�5�#�_��M��i�^��]Eu�EƩ��7�����褜�g����p>f���e&\����b<ZG�6���С�6	�9�G��}�D��4�*��8
6@[���7�Vk��<����<�R�!o�5�`c�̟T�	
 ���|��L?y�����~4�Xe*� {���*�����s�6���1G6��xW�D�-�T�/��V�@���k)���%*��
VC��� P1�Y~��`�:�����X�����3;�A'�I6�Y_��SR��W�6G���yHׯ$>b-�ɵ�ߴ�� G���|��"(;I�ͦ���=�����jJ8n�d����lbU�y���%8w�mŽ~\�Ygn�8���R��
8}l�"m����l�� 
�̅�p-��H>�����mxo�� ���D2��S�t�KMV��c�A�\�B���\������O���}���|�H��-���<
��u*���Ji\���Ҍ�#1*�r�'�0i����Z���!ʮe����EM�;����hO�I[A�BQ}m��=W�^��E��}�fU���e�!��Gqkﴐ~𖽶h.����F���]�c�j@"t���w��H!��/�;����ū�&R�6�E<�ٚق�xaU����m
r��`�LY�i�):�_h�
X�x B�����%vQ�����e�T�j�lh��kva)�ȼ&)�����_�{l�~�,��B��"�1���(q�x�oM�=K=� �~p�x�yn�m����tG�i���}krA���w.�gq.ٞi���+]�.�� �B�Fi���J�&�p���|�{U����>�����X%
��)�t�B̂㵅��S��l�y&���V?��E&J�m?Q)���6]��DsÄ;�AqO�N��`AD	��Q"��H������{�ͮ��Y�U���9Y���G��tz{1�ۋ!V )�_�ӆ^!���z�����t���Z}d�G�uҔ%}aE�����a:�hP~3ca �!cWl�E�©⌶���mV�����'�w��̫TrpVk<�5���o��=�:a��R�lil����`��_�}s���W0il���A��?)Ub��	����< �2�b[7,@�nDL<Q#'���������9��{��R�)(*�a���1C%�bzzۼj����;��s�4V>Ҍg�D�e��񽃎�����2���z�{^7T�Tu��:�r��kIhY��P��i0��3^'=�#�&�~Di>�+'��r������P(��{���&�*�=�G�bͥ�&y�����ހL��] :�x"�8竺�}�&��C��A�,3��T��{�J�ܠi��P���ƨ�z�Hаo������2Q�n���g
�"�5B����mg���䵗���n�`�5��0��#]�P�iX�AMS��p������3iC!F��N�q�2琥�ch@�ș�@��[&�1����è�J(3i��e��"�&^M��̝9A��C{d��ґ�$q�w�-���O?ִ��Y�9�t.���/:5��y+]���������* h־:�HThG�6}��*B=�C�j]���� �ɏ�݉�S�$�9�瘙�ܔ�`��ګ-cU�6f��{�	�u:�泧�������LR�-���t�X�5�p����y�Ց�Z�h��j����T*�l07�|�A�ML�ԃ���`Ȱ+�)��:�o\E���.�XVC#!�GD�%��F�YN�j4nҌ�%F8DNu��9g�@m�|z��:%TN���(-������o��~l�4�ɑD�Hf���(�ě7�#�[>�fs�%\B�!��xZP��]¦d-Y��oW�1$]ŎC�F�dK<�]�3]9urF�}�'�������7@���Ld��J���X�yN����i�:���:�q4q/�y�OI�� R�j�w�)���	���Ȧ����5��A�c��)&E˃�UHe���Eq��
C��õS0�;��
��P����ä2`�:s�O�A�[���+�H��.g�*f"m��v���+i�H�*��y-BF���a��`N}mg�v"	rJ������w8PT�/21vG��ꯏn���Ʃ�~M�ǸS�7B���c�t�7O�l5�n��i�Fx���H���ҧTޏO[1b�� U�2�;{�^"�J�;��m��A�8�u���k�FMC�v����M`
|��{)��)F4�
�]�:!�0�y��xcު��d́Vy,�b<���h;���p��>.	�f�u�qW�]��φ޼�q�du/_�x�_�"{�Y���� ����V)��M�E���\�-x��Fi��]��rG�t#�%�Pw�ń�ZM�I�ߍ]0x�?�� �Gd�g���j��XN�|�s�e�r����XtҜ�~r�O
�I��|5�N}��}M[�O�]HMX��)��� ^WD����W���K���H�2�{�6�i2�{9Y��)(Q9����������('*&���UI�kv�C��ӭ=pa�NCqO�|�P%ś���V�̶;}}�Q%τD����%YJ����j2��VX�c��
#j��!�<ok�a�~�\������3fMϔ]W&�]!	�-\ff���o�P�W�G��7���-H�abM	�9 �G�G�y	�ϜH ���E��U5[{�I���+=v7��	����_���P'���h@�f����B�[��ڥ9�\��ezcwTًE8Ą꣩��	(x۫��6U��=������)�tg��./��	�fp��vf�4�G��#'�6Lr����G	3�濗l�"������W�2/�fP��x7�*v1�f=b�u߳��c��2T��׍@N�����S罜c�Cm+�x���h���ş NN�Fw8��P̶����p`(bT^�Z�K֗�D���BH�m_��6ܐrb� )l���(~`��H��.F�7T3o�� �50�[ދ�1���qe������V5��<���"�I�ը�b*2���{KG��T����g�,�qu�~l�FeQ�\�Th�Y���b��V��+��p�}�z�#�2����������cn!3���)��)r���޽��K����gY�л�ZP4�/Z�!ޭ{���h~t#���a� ��CH8�����T�U�4Z�,���	�<<���#��]R��R�Y�@�pJ�v�|�r��/����e����9hl������3d�|S�@c�g����Fs�F��9v�r9�#�J��ꯓ�=�5
�or�NC�d�	p��H!Y�u�7t fi3E��]E�"gx���H�b���ބR)�Z���9Ὃ�p $Z�e���tw��ɮ�Kܭ�V��K�>��d^��Mh�hX��6^	�cU��D��F��uJ���xN@�1�4 �`ε�J;��gx�i����AA����gOJ�ۺ���%痫��wfkyl��;mm���~|�X6m������?3�s�K'��ҲL�$n���|c{�)�N�����qjS_��n�3�p����_���ш������{��	����)�m%���.���, }t�m���-y��q����bV/ө�,�f�2�$��Εo����'���o�Q�1	��zd��Ɉ���j<%�b�S�I���^�H�f̊ҕ������,���%1GQ��4/�nA�YbV�v�pA�G�yK ����F{��	OB���j��QcB��m���?-޽��k����b��W�0�.��Kl9n)��b�CA�w�0����'�7��\et��f�U����S �S�?C�j�V�T7��n���`s��~Fz��RCG4H�[�o�楕u4Ҩ��֗�;��U��<$����hUYsQ��j�N����KI"��7h�mB�Q_һ�zJ����E��5X<�PU�튼�~�*Tx�kϧv5&��
qj�-~`��!R�|�8ۂ!*䳖K?�W�E��t�\h���zZ��*7	VEņ�X�\w��ҩ���Y��
�B�#�GWl����Rα���B%)�I���{�dI�m�E��t���n����G�����]]�8~��x��/���x��j�4ۯ'NF�k�8@/O�2�)���"����B��
/�T�."SԄd����s��@&�Z��>�ӻ'����[,�1@S%��J��"�?_����'<f��@�1Rd�J��@�˟����L�`h,uvI������^-!�5D�h�u@�X��`�G��5´�ǝa"욖9�>��S?����}Á��ɟ�mj���^gԤ.ҩ�A�M�'Y�J�}Kg(ȅtn�Aa����A�S��3��~��.?������~eH"�A�J��	�Tϫ��U�/(U�Es]E 1�'{Q%a�NQ��p����.¡@-|��`�"��1BC��Jع��ʅ˂~���@0Sgۯb��?:f�,�Vҭ"PH��j����Kow����M_4U��Sx�/��y���D�h"dbl��d�3=6�tf��/���@���qؙR��C���n�^�ON!�\I�&I�*���(�.yV|&��W��E�z����3
�����;\����Ծe_�c�����&�*�:@|@1$�Ӡ�@�P�䧐Ńo��y9���B��D��C�Y{���4gM���7&�67���`*{M����V_����}��ˏ��Z�2 H	�0>/�Q��,*j1�Ȏ)$u+�d�q�eէ�ɵ��*4�q[4��T��ECh<��c�pa�h�h�@�ܦ�F|��}(����B�2��-\������莏h��ƀ�����OS}`�&�B�·f�-aN���Odm{�md�~���L���)�/e
��(�I埘)+�{�*��>1/J+v�àD��l�zb$)��R�ܛ�����\K����|(@N#6�x7���L�
�^Ͻ��s��� \A��ep�K�4��g�j�M@�M���u�����￫����G�MNQ٨�W$��`p��lrK���mO��k6MyI�?#�9���LP�CQp5â�s���Kf�J6�U+��n/�ʌ���7����(|��=T���j̅�
c��68��������]��(�;���b:s�2�}�Q'Q_�KO۵�="Q܇u�&�����C�<���t��B\��cY/[;BS�l�*Y�:����a��( l�����|dR�
��:`���p���e�Ew�\��Y�4�ya�J�gn��;;�GM=L�%� ��� r�4�VK�E��Η�h^������Q���%(��������h�5�m�Lx*�.�
�n��J<�`nyD���>1(�[�c��̴_r���Zr)ۤs������*��`�|�֖���V��H��g�
٥�H�K�=R�vW��̓RVժe��ȌE3��E\g�p��K�^rʞ��Z�;�p"8�J���0ћ�RV�A��%̖���]+��b)��e9N� ���р�5ph�0��j%,�ߧ��-8�?c��58��Њ�C��$���iQ�����e��AͭX�`}�"aO�NM%�CEI��V���P��!��ex�e,�@pd[����U5+�׫�f��<I6>H���5z���߾��.>�I� ��n����A0y�J�r�d�vI6�<c��~G�Q����P[ܰ.�+�f�2���U�	���繫���~{E9E8ثZjbG�����T�Q����[s::�������6�]��]�F�=dn3�wh/'�iǔi픤�c-َ�6����U3}Hj��vB���_��O!��������^��U@��< ��V��u>{h�g5�)O���;�J�N�Է�
��R<�݅��󋂓Z��ǁF"ř���D��,t��x8��eo�&��>�q�lq�p2}�Bߧ[	.��A¶�xK�����+!�'ڪwj�V^ \��Ӻ���%m��	��`��.�L�ys6e�������f�7��y�q0f�e�������/�dgю�k}�����}�čƨ�-�ZB?Z���P����b��WVC�x_�>,J�A��I.#N8��-Y�oT�%ok�����ȁ���*I��	n[�,�>n�Ӗ��CZ0�y����9��~��w2��1�X3������9�9�Ywϔr;؅�-�X����24!ې��*���y��L� ҩ�ʃ3�IS�a��f�g}�fS
T�θ+��exJ#֬rwَl-gK�>mU����Gݺ^t0����5г_N����`�G{xZy/�1N-<�ce�و�G6'���/�Jj�(V{�Ä��2�<f3�ȉԴ�CT���(�\2.2�GX�\���$%k�mB�����@ �\l�Em�XAS�L�3�A5Sn�x4�߇'+H	e V@��D��`1�l���%�êAL#���%��Ջiz�@�e��/�gQ_�w��'��5	�5��V�p)oD�4�7��� ��o���
Z�{�>���tw��(cY�(�J;��&AT���U^�Wh�dX��Hm���nT�֯E��?.HA��[tb�}�b�I��>{i���4gr�LPP����p(��V�I/ZC�y�P:ݥ��#� �35�u4�{'����o�C������'lC���'fӉ�����z��\���&9�xA�m(|����V��Fk�i`�?�w���ndk$�ӗ.���*�l^<<�w�����I�y�}�PZ�p�\���Lu��i);����:���_W�=�	g�$l�������>��x���b:(X��O��ѷ^�i)�'_7�^+U�k%��z0����$ ��t�����Hw5�gH��c���n}� �o��3����:�ʏ����7T�d��HxÁ���i."8#�f����RJ4n��%7��<=@�NB^�Wf	��ȻJ��q�8���ɩ>��3u��Vc��cNҠ����8 ]�h��(�c-�	��j�}�Nb����ZJs�����t]͜�x_�-�=XB����8&D���`����vn�/���r����/�"���!��Ubl��R���[�s5��U��6H�[���t�A#Z2l;'`��r\M,j5�~K���ZR��{�6��u�ŏ-s�2���?��md�B�Q�p��֏UЍ�Sf�oI1�z�Zx��$�X�Pyl9���q�b��R-R��	㟡�
_~W���O����r$~� :,�_1�Yj�l���0F�p|�.�sղ�P�4��ٺ*�����e/�@X5j=b�lK�:c<�p��{l�n\Zq�{�=*�@������b����,�T5>"���4�NS��xTVT�pf~2��]3{�]�.n��b^8��!�i1Ze�-kj5��٥i�^������r��^ �^�%�N�+6сG�h��+� �=���-��(d}N�l)��YqqWm5�iӽ��߭)10�6ĔUD�͞zvd5ma�����G��ōi�vj�G�%MeN�'ɷ/�	��Q�cc�Qw}y�/�0.o�/	�#�q��zV2X���r#�
�
ϒ����G�X�,wB1pH�hb5c34��ގ4�-4�d V�d���/GDnpIrRvK�M��}����2ac�HS�Ӊ�L�䍁���5�!��e�\�����UA�][3��������c>��y�v;�h4K���q�.�w#}�����<�e�v�/�06N���k�k����v�5��*�����w����<�*�aPX%<���Q����������� x��siyq@��4=?P�(ȇ�<�G���o�=��E^��m�?e
%��Hf`��
�n��Y��`ԞO$o��e4�M�cO����gO��cQ;���"T��C�Ӹ�$0�u�	/��礗V�+^^P�ѣ��������&��;kM��~՚�*������H�5ߩ�!�V��6�1G��llJde@��|�$/�i��E^U[��W�2�9��e�UD��
��Q�j�rU��J����Xq�|�&����l�[U9�B`�F�c�u[m�92�)y����r�1����ͣc|*U` �#�S��|��1�J�)B8P�xW�`w�E!K�"2S#��'6��ߋ�j�3��c�Z1��_�@����� ;�_���ę՘X��ie����>��٠J�8mد�M� �W��"{��ԆDEݽ�8��Gp|��5�j�'[��[�\�F�N�<�HE�Vo�!�^쬝\���n� "�.��]{�͍'r�%��5������&�	C)����AM�x��+;.P�{'�����8X=w�鞫D�+aM�Ɓ/��Qr��3c��4̦TCo*8�Fāƙ�?�ۮv�E;^q�x5.,�� ��~3?4W��v_]����n�^��f��g�/�T��Y�h��
w`O��AO�&m��i���x�EX�lq�p�
N����2FiC�2�x��I�^l��[���y8��)Df6 ,���8���$�ܺ��� dvȁ\o���"�<��]d�����0��>?}���5ƌ�����twy�1�#�{y��K.�~�o\�6͸z�`!��C,���f�O��'N�w��z҇�)ǟ�M��u*m�`4�Z�;E�([���T�X{*�M����=��@�[5s�؎�F�@��{�~�D1��vr��c�������@��u+XJ��R��[D\ҭV�{�����Dpid�e��y��YMD�(�!o���A�6��z�j/��'�6��v>��鞪.�գFk������\_3��wgz����v�6|eO��Ҭ��*5o�7����V�O}(SB�CV�wK�-9��Ļ��,)��IN�2��O+*c��v�б���ɽ���'�h��g���F#� �V������*��]��O����.�'ڏ��R��͍�C����ZZ����f�v%�qK/����Y��S��\�>=`}�Ԅ���صb0��5|�������(�Kä�0>�X�*�;%<9���a�E{��Y�,��&p����{v���x�T�X���rzǔ�U�ȡ	n�nYb.�?E'#�̟���؝;T�А���"]_�߇YSZ�:!(�9t6���Toz+����oL=6��=�Y:-���㌡e9�|.���R�K��kO*ͪ�igK��~�iL.��?W~�]$��ttW�O4���A��Y���yn�{NRD�ml�n���?��D��s{��,�������T�	+Hh��_�\#9�SlAY��~�҄�wNm��ؘ��KpIv>oH-�a���N�/,���b�m���МY�#��P�F�2�8^�+��5�ϼ7��ެ�A�+�n����km��=A����Y�AĮY;�Y��8Pd�pؕ�[Y0�'�K��=G\��6��'����e�ل�����ve_mYQ��po�����L_�����q�`	3���|f

�V�����,C�=�@Q�AmUx���w|gj�<�'�&�mi�؝g��=�r�>(L�g�]@�og���ǨN� P��ö>��)�M��+JL�a���e7iy؆\�9vHі��J�=���|���LEϼ4�tpK�����2�3fofSSs�F�[f��h+Gq#������	��JԘ�D����'is0����J�:��D�An� ����_���L�jv~�*p|�b�zS�<{�"��\�"�z����_v_� �E4�2�̉�[E-�.�(]��vܖ'���4��ӈ=C���اǌ���w �	�6�2��C�F���y}�u����/�k��-��A�{��(O��[7�;}Z�u.� 1#8���K��J�gd��Նdη�����ɰy�����6�
�igP}��:�hyw�x��{~���"Fec�S����3�rMS� <k�0M9k��B��pk/�=��T1�����v�!��u'9����t5)�k ��ٹ�_�#�~�wVFך��v2��4z��q��c��nN�BG�^�B��Q9��nMf
s��X���1>凈9#�`��|f��X�<�p���B��/��i�iː�r��#�O�cS��>���G�8hر��ǒ�X�����.Ea$��n�L���5n9��h1Qd؂E��.w5C�R�����T��ql�2i�i������d����hg��� (�h��I���@�]F|�����ǃ'U�Ӟc�~ҥ�K��r"H� �>�"�S��X��s�O��F����t��0Η>�ͅ�� ��΋�C@�=/��)��l��U�;)���	jw[%8KFa��!8X6D2�Y�iNg�*�s3��?Kn�x3����B�hCV�sr���KSy�#�X�����0IH���˰u	Z��pfDm�9�=�.�`�,.U� ����֑aX��+���g:w�>�[�P��؋�@t��}��'bŗ`��c�;�����VF���Ğ;��X/�CZ�*��Cٯ˹@���>�N��{��HB�Pxc �'�FW����A���*=�������F���r����]7�j�ܘi,����z����ֻ����X�QU�����a��������|׬Sh��6߲B���_��C6}-�����.>7�y�i�L@T�t]H震�7�o{T���!WB���3�*
�r�vF���)늖��z����б����U��͇���Q�bM������G�����e7�d����-��М�!�=r!�=���ډ��x�d�&���⤆g�i��zҁ�������Lq"�H���Ņ��z���Ϧ ����v�jl` W��6�4�۽T�gy��>b}�7�JC�Q{�=8��������ϐF��<18?]�h�3IaK����%w��ۍ��"XQ޲S����0+�>�<�%�]͛� �f��3-Kω��ӏ�kܘxN;B��Vj�~��d/G��Qx��rܼiz�z>���RC�H��|M�p�"���q��u�����"�^o���o�|($Iq���Iw5^XX'��|���l���	�f#9�\Y�E_��?�%�W����{���)<�~�g!�+y� �r��	�ݗ�S7�%����f����<jվ��}*�1-+7c]���P���"��0���e�II�T���I�1m����?�ӹ���[u8�(7?�f6�s�ESg�&ȮܕwA�}�ܴ��1��M6]�9Ú�e#J�d��F��t�ڻ6Ѫy�P�>��)���mP�����7�īL$�� �>�"{qR^l8��\�m�Iؗ��>��K��r�[+�\�PW������L~�I_d��"��Em�E#�q/_i��{����y!s~�<��{ヘl.?V�ńϏ�7�?�Ȫ4B�T]i�S���]T���R�5�+���˨˹�����8��DЩ:�S�@���hH��4Vi�;M9�|b��E�w�@�F�yGh_t+_ű$�-+���9~��6a��}#f�%�����><޴+]�W k��,7z�ŕ�~X�8�������	yGe(����p�;3a!EHOE�k��I�ϷE�`�{�6�A<����~���﷍��X�S�g��%3�K��y�i?/��oe�&7UA�H�K�;_$��z7�\1Ç0��ve�����O6_g���������G$ݮ�X�jV[���̭-Z�ʒTV>R�e�	��|�N8���vBw3��v�'˗a��6O,X�REgD�{Q�x�dή�>�eu���r{4��0��xw��f���e� ,�~z�Є��U���5�	Q �}�r������w8��RRu��-�������}�y`9(�{b6��g��-�[�"agCGj�%a2�NZ{��X�?Q}	�.��L����>~�
�}��h֎�%��ӹ.%�t�W�4�*��,C��8)d�1le�G��%�j�K6��G�q	?ʥ���-N��q�1H�v�-����U�;��g���Ul8DˍK�K�R0��y��W�Er��]ˊ������p������=B�~��"��vl��I���ə��t*'�7���oh���a�:��>��qx����_zZ�kX��o��?��$��d�A��L��#�'1��Dz�sK�c"D}uV�\<ma��ʂnEx&�ɉ����P�f">�*�x������ע��7%��O��z]�茕74bE>:f"���n{Ҩt�PCH?Pi�R�ل��t=.��aL�����&YmWu����I�e��.���W�K4F��O�f�f���<n��&�u�d�����g_��G�-���O6�x�2F����N�m�tGA&;�7����h
(��3Վ/��g�h��,�H4��)&�?S&���f;K��ب����V��C~B�R�%Lv�������{�a�#�7	�ID��FlE^H�0�wʼ=
8¢��c�1��;������{/����Sw�1s?�;Ρ�`����}�Sod��1��<R���O�FD)h�N�&�)�q��9�<T?8)��g��� �/�}Կ��/?�D�;Z�®U�T�?���.$�����P=r�!?�͞'�pX�8ד�����cW��7��"IۂZ� pO�����6��*(l�u��
xV;e��e�K�fF-M����2h)������Tf��ut@l���E�����j�c1�����y�����k�NVHv���`^J֬)T7�:8#V��)�˦I�O�����R����e�u^`���U)d�6X�Q��U �[����A!j�	�SggBӳ�\/�j51��$A_C�8|o �+!�K����t�h�s�_S�U[I\�ˁ���#��B�����7�.W[�a���6�k΁H��WB��O��S��W��J�?�u�!��`[��u�4o㥒��/9K�]�8"S�h�i�����}%�N�F�||��N�X�^��ӂ�H��h��Gxw=!��W`���Z�c���~P�G��N5��'���t	�m�ǻ�Zw���̈80�w����"�/�G��̪�����\q���Z�h�aȦ�Ł�{#o2���#=� J{_r�z>�R}\\9,H�,B3�19�٢���&6�9��o��u$ �~BG��z}?�0u\�}�Z�k�[�-�=���&B	<h���!�f_<��$~eiڝz��ɟ�i��������0����o	%<t�263,��4w�>��� X�2�;v����Te�C��)��%Ǿ�Ri|C��N0Z�)He]���]�;Ns�j~
B�R���]Pah���r���~��t��4���R>�ks{���:�̝$��j�K
R���R�C���j�;dA;��LO�7|bY���w?��_�$��[�X=�Y�[6ԭ^d,�wM��!��#�kV����Eo6ijY��\=�?	�t<A몍Wa��w�ñ�T,H��\=f�"�q�^�L���"ߓ�)�\���םb�~��^֓�\WH�[^�T���
�8��+�4�e��:<�u�C�D��V,��� Di��A�.:#�\����}�>ұv��:�z�CFH��^���/
�]�k�r}R{�LC%kƕj���5�H.9�C�u�_��0Q6��N���L����`ei�v�`�:��e�������&&c���UJA�JG��-{F)�+�������35�1�A�3��⣯-�y���A8a�SӮ��oV�4>�޸GC��y�E�J��t�����E���~����˹�F�5�<���49��!0�P��I���WH-�S^�Z˪��9O�����U&g �3̆*���;#Gg2]ǥz��B1!�F�h�F�ZB�;��Ɉ��}T\��^P­����h���F�
FgM�S�����~|Wgp�tgE�>�t�PTU��v�%�j��L<]<�~I�(��l؀p�H�_3[���*gH�d~��G�$3��iӠ8L$$8�2��A�JN#-��U΅�0םBI8�ε45 ���4����Ks�-<Dj~R�e��g��)�\��3&f&ԕ�J�Z���V= ``
a��_�j'�e�[%h'm��ƍ����=S����ns�c���� ��@��=~�Y�͍�f�@z���,�;V���3�~/Z��qi��~$��ςs淼d���-��
�M��lp�k4e�eN�?J�t\8�����=1dg�>��"pF�}t�H��Ł��(v魵�p�^��+|��\z���B����Pı���>��E�8����v��w\^���k�0�d윝�����5�GN���E�"�+l;>��D�q�XSV��t�zV%Wޱb��
���k�jU�|q������羽e�c�Z:��:ٿ���Q=�X�C3�4���D,#�P&n�w��C�pCۍw��V�dhǞ��e��A�S��ʒ���lq��8-r�94���[�]z%B�� g^�s�a��¼'L�U���J�2���	߄� 
D�U�h�w$r��x� .	����s��@ր4:W���+8��,��<�`��Ҝ8���� �j�nkmCņ�SѢs�r�ģ����I��%�J?��!�k�aC����B�R2�ւ�Kj�h��Ӌ�y�p=0u_�^�����@�cF�~�\c������-o[t�����Pk�i�^�֫,��;�i+�w����S�-�j&ק��~C*�>�~ &�E_�;�#��@��G���a�S.���4"�b����!E�+��E���W��=r��~R(O?�
|�ڣ='z�U�(!w�ą$�L��C�s��Xa9��!ǁ`����[KSY�ƍt�NKBO�n���-U��c#��2�u����5��g}H*�3[{\�H֝m��ZRQ�|s8~S�n��U�1���m�`�tr��B͓�W�k��q1�2<�TD�u\u!��"z_bN��w�˘U	���Y�n<A�^�-�VRn}�;���.�A!X�v���-씦ob���:�X�u�B�p�-șLpi-������#���i_u���1�;�Ao'�0�|N���M�$0��_�(��G�]a�B�vխ��D��0
<U�����[�4D���Y� *��N!$�r�>�`j p�M�a����47,UkA( �N�3�<�� ��:{7��Y���W��9'����դ��~�U G�B��
��?	\>Mm�m�uP������84�B���bKUc=Ǟ�ɸH�v	C�"�k�_%����=Hf1����|u�ʺ]�D����q{[U��C��k��!������4��
���fAo��T�:�6�E%[|)�3z����D�<�:5o;WCX����o�_��L9�o}S~J����	�4I�kU�D�R+�Aǃ�ݯ����0�k��&��l�/";�q9Jj�}��t��sf�E�v�`D��Q,Y�i�4����$mb~��_���#�m��O� Ң�J�G�χ����+����Ho�* ���Zd-(kh7	H}�g��3o�s9�o�խ�V�P+�z����f3&���ar���'�/���sD��E���̩c�w��"	�#&A�d��9w�K|�Q�囂Nl�K�ʮ�q�У�Z���ȵ��`���\ja�ᘩ�7���)z��S�z;����F�4��w�ǚ�QU6�@�uZ�fJ�/�~��Q��/������Nw���E�Fl'D�`M��N���R/���6�F��ʈo/��V�t9���>$�h��i�]��>4|Cw�Ǟ�K�1���fG˅0�c5��O3n~�Q�'��0^�J���N����5�y��4OH�:��,[��P��mi�K�.3}ڷ�=C!O;�N$pK����a�g���;&�m���p�����"%л�h�v-������J�٤�:���/k���k"ݠFRH�����V
��16:������%(��EZ��[I�6&�a�Tla�-AFBSI��}`a�Y��8�y��5w�Nݔ^w��Y�ZB�����QIQ�������w�3Y^���P9&��v�p*��^;��^�c=UW����_v'|�`�d�Ϊn[X� ���{R�w�.T�S,Kh�9��5�`/��Dġ7�u�!������0h�cՕ����M
X�*9�g���ѱd��Θ���|Y!�A�m���:�C3�Ѐ�p���������<J�`IwUg�3�[�V;�k�E��?0^�����^!�RS�-���vPh�a	�,~s�S琥�}tLU�N-(g�Y�m%��"jK�m`Ŗ~-����a�I c?3|٦|Q~�<u�^�>��� ��\"��* �� �w�k�����	�ޅ6��էY�j|��խ�u���k�WAT-tS�7��&ň����ks0�3��KM�;�Tr.��Z�]�7��%c�~�s�y�˘�B2�JW�e[�_b���5;�:�:���<�3t=f��uX�5l��%������r��c�	���H��B��7�Ȼ��H��,����[��Cy�(W�h)��=ȴJ Mq����Կ4 T����Kb�'���F�[s��b��%'��bg��^[K��9���x��`�c�b����o��k�,�d`��A�`���S+��{O�,O0B狮���N�M�^��\\,���XR���b����{m���eŉX�&)=�'�=q>J}$�`8�  Y)�����'o�N����̚dX��uk�p�G;�8�cq�ݺ�ٹS3�p�.��I)��s�!�\�����f�Q�F�g"���jM;A�8��� <%I�������� �N�|�q��ҍ��4�+|���j��po�@+��8�(W���ݥ�R�g[1AMycR{�jm�_|t]�����}���B���u�))"�߷(>��)��Ȥ��C�П�ڤW�l=��X�ӛB8nsa�Ü>�N�is�p|���bwi���n����Rł��yX�$�'c2�o��'����ii���On�ލ���Yg��+<q	-��]J�!���Y'�G���4;Gc���$�B����W�HO)7v����YZ�8�{�.k�R���8i��fX>�����ɘd����,<5[e�\���	��!$���0[���e.c��)�%�Q�̨h}����٭Nc:%�Ah���d�xfg 1-�}�Շu�A�K5��?M���.l`�����eð�]W#]r4zV�o�D�@軤��|�f�-^����$�ܳ�u��ł�In!d�����u�/��Q��c��+$rs��N@(	#/�Dd!�:(uQ�Z����E���3�������eh�X�l�]��k��贄��^d��4�������	� W�� ����+&bZ��y5 {���ć](��轟�g� <�5�]լ����~m+y�P�+�a�MkDF[0��+���gwRV�Zj���"��Ѭq8v�1���m׶���F��C�f��{v���amT��2�<
��'�C�^��/;��B�@��9����}O�|���].�	�����5t�����g���mN.\\�O"`�f��ӷPcA�+B�"��8�2�&�T�-���	W���:N��n(��x$�݁Ӡ3��<���|����Y���W��3M[��ef����ݨe{�3c(1Sg 1�:9 �Ei�GE�H�9�O�a,.�r�<ڣ+�+���kؙ��\�a��7����t���t�Ѵz�@*YNnL�C��|^@�!�ѥ��v5FV�SS�ݭ����zv�s��ٖ�2
���U����I|�-�s%\�o�r<��HzUGɑX�AG�T���ԃ;���jlB�f٣S�iUE�-����Jh4�̿X�PE`r"���k6Sds���Fijr��Q0\;s��P�~!��J�t���cw�����⮊um$� �����ʄp��|s#�����C����~���=���xd1�,'����`�]#Y��t�C�����K�U��~]�`P�k��B�Z�pD����sK��f~�+���Z�(�1D����K��	ŗʴ>05K$ʓ��#�P�hy]&���&�~��z0�^�5 sY�����
^gw�!tE:=��*i������ٰ\�O������O�N�)�>�s��P�5�u�rR�S_zX�/�r�_�r<�m�!��W_"!?�<�_7n�`��[L����ӏ�-�;jyj����2��_�_Ml�6�_�dX�8z��i	F���Q{�\0.�b�O:P�s�o{�X]���BI0��H�;�L����!��^��"W�_��������-B�%�&��Πl�v�L�t8��3�g�\�`"z D�}��$u�8��It�������l,�=/.J�VO@�ub��ț3���/����qR;�=�[��=���%*Sރ ,Z%{Dz��`ba���s�eD4C�����sI��7��������r����s�l���\y��L�81F�V�t���������I��vj\%��?DD f�#ڿ)�_�ݪ�L�U�
�ǙY����}/�R�%��YeRN�+���u�L?��������a�%�ArU+C@�ԃ,��ܦ�
���t��z��^��n���er�^�k.C��4h8Ы�+p�W*#�S0���ʳ����6^�v���e;�5>�i-�`���U��߸���6����,F\Dfx�z�kqs#1j�@��nu�_=X��� ����ΐG��E��Xu�DG��-�q��ϥ��wxp���28�j�?5jD�\�cR�N�?��3^.�j��I�+2�*;DiWa�o��;c1/��aC^�����N�΅F�T��6PV5I}��Z&�=�[�v��ؽ#�{�vX��u7��l�7�-�L.�
c4�UO@���j�čw�Jb?�y`EQ�t2�R�>������
N 21�8�e���}z#s�p1'��Q5������0P�<]��D}fkAW.P��/V���+QL�J󿦉d 1"ә��q[�.x�T��h�G��e�Ov�:1 
�fG���A-�[�ޕ;g�o�w��nj%.�I����-���w,�`/���$���XzڏZ������-�U˵�ܧ�6����>{�//p���a�dǶ{p7�z:q����56;��:J5�j���w�/7�(�{Eb�{��ܑ1�:�m�5��[j���W+��mI,��7�������J���O@��.⁛z��Xc7\/�r�Gn��8wC~��01>:	K�r�#�H��q���;ĂE�m�1��M������x�k��@;$~����[�u �e���0s�i+���D��<\T�)R5�����b�T�O�W��zf7R�geU���U�%e=��IEB� J՝�|��ɭ����w��e�=��$�`>b9:{��4��*�6�F>��H+����bg��̙Rc�M.3$�ƺϦWɆ�,�g/���W.�B`��o]s�VW=�}ʝ@Ά�;���	J����KɊ*��v"X�'��l�Zt�a1OU�9r�	�&QW�my��z�Ȼ��
HDV�Os)��FV�N�xJj<X:��~�ۓ��R޲^�ݓR�}b �t�tv�7o�G���@��?��E�&C�em��&���|ǝYU���p�����o<jh����D�~�Ӄ��n�,y7LS~M�8�S{��!7|�� ��ڝ䝷����}Y���]�s�ռf���XE����?
M�ߍ��kak�A�-�]�mw��ܶ��l��Q�m�7��`1����w�.֬ ����{�z�ʫ�-��3իR@ǌh8�*����_�%��VW�S1`��K�x_�" Aߏo�3'�����m�AP�_�jԅ$ի˞���,�e,�K��o���#�%��a&��S��Q�%g_3��'1���ӱ�z���˾�puz}�\"�kT#Z��I��+W�U�zJ��y�~�U�U
��N��D���x����JK3� �V�]'D61��1�Q�7�@#���MD�Uo��-̈>�&�!���3�G��@qq*Z�}���%��Ld�|+�,@������T�u �e��?�l�ݷ`�������t��K+T��B�TӫsT�2g�ssLk�g�#:Y7@qrN����$�+'��V-C���ʆ)�d`8��b���;_��к G���vb��]�cO�g����K䘾�@�f�kIn�ִ�W���a�kx~AYdsD�b�߂���8 �2��U8���~B�B�W�W?*E�#��,;��i�Y\ ��;@jZK�����dGu�_Z��V��,�r$=�C%�𺥗�L��&BE�?�&��o/{�֗-��rDC/�G֧6����d�\�� �!�I�����@y�F��|$r5��3�=O�ESy�:�G`���.�rf�n��ͥ�Jr'��?a�c�9�W��FgшEU_W�
�\�.�q�%�ӈR���8���e|M�.]����eu��z �ڸ|�|�|�\n�����S�M1��xsW�N���H��I�80�J�<�� �.|�i���R��wB잨PD��7��e/�bW]��>Q4p̈ȰtӖ�1q8Q�k�����b��A�p2�cx�_��5�C�3�Q��T��-W�;���&���͈�p���4��nǑC������Km���K�}����<�?ٸj�<��!��ڧ�"+�I�Z�p!�ܲ�g�
��&��9v�tm֦�)v�kA��@o��Mn��m��g�����2���3����;N�7�����|��>�M�4��Km��.���xp�ڲ�"D?�ؿ:�ڭ��	Q�v�dwY����a�A��"�߅���:R�#2�Ҋ�qNl+�e#��9/���ˈ#�.�=�O�&��j2�Mq�a����¼:�^�Ɛ}��! ���_n��q:~=���H�d,JO��U�s)�H[F�����ɽ@���{�чxʺwS�N!����:����pl�M����]�*+�;�/G�:n2�@C���9D�Pj��qŸ~I�5�ܙ��`F���k�])	��l�"*�Qb�n �����8I�jb>#���K;yx�V$��Go��DʢUv���
������EK����x�~� y����/�tG�W�>�p"	���s5��\��x�WWsD?ho���g��Ra�>� ɞ�6YȺ)�M�jP/���8P��/%l���Уn�����(^KX.z6��Y�;^�)i������e������B&�D�M���
�#��]�<L�iV&(��`�O�H���ȹ�Fh������!J 9�*f��pAR�|c�H�pTsz:@�r��v�e��#?{��a��9(��oa�f) 1�m��c�f��{�:�=˧�^ܬb�\�-�Z�3��ʛe-5��p\���@�N����ީ�9p�˱f���)�u L��d�#��[�6-6�5��t}���zu?�d�a�U��l�ǲV�3c�FIW�PIs�b4�:�n�fL��P�N��b.�Z4���Ә�f���SR'/�P�������F��C���_i�n�$�(>B0��?v��'-����B�=��K��/��}�:��+:�l�n��<x�D8}�p�\K��~B�z" c����G�7�z��E¾��N���/ݜ:󈨠܅t3f�D��x�v)e	��h׆w����m%AMN�&!a��-j8pRAC[Tl�v�P�kԃ����h4@i�@M���TD��$9s��	��i�����Wf0�zl�`��撳͹���95h�M�8#��"�f����hBaV�A�_[��5��N���c(Ǥ����bH5���>'��S�k� ���	����h̾���)E�>��}'�~��͙_�ZY �WL�����nu��l�2�ɪ��sݙ�Yb��B�H���״!�N���#�SMM\%ə/Rć�`����<k�~�*��M�H�lm�p20�^�r��r�9W�:þ�H��-dA�x�]�.��ۛ�?���V�B����L�@�ء��g�����O@y>�BD��,R۟����z�S9��=[�J����#n$�W(�y��4��sge���%�cn덋ĕZ����W/�1�v/Cc(p�q�Y��e��:���cX��S����?6p��@7���C��f9V���p[�5�����"Ɩ?�/+��.�q#���w����8�V��$��C��Q��b��u4x�ps<�:cq��Բ�ʏtY|�d�V\�m�o���Q�:�#��yYq�[-`*�KA��I��r]���H��S��|�QK.^�wB RA�ҶN�[1
��u���U����w��W�x��>D#��ER��>b/+���wVKA�圈�����}u��^���T�+��Y�+\XS�C`�	�%�.�\�F�Ԟ*(k7��5�6b��_!��XL'Ƶ��~��9�~9a�{8$�V�@�u�=�$ڃtF���n��Q\E��԰吏��G��Gb֜�R:�Z�����8�B��Θ���]�,��!U���p�S�\�T%�"P�nO�Ic���4v�S^nκ���/�Dʶx���3�Bʃ��|1��Py��_$���V�p2��h��N�3�t˧�d>]^�=@
yZN��U��<����W#���#o,ڟ�. A�!Z�u��J�6�#}M�����G?�����ҧԘ�޺���;����e$�E��	��t�-����B���D��"?��Iâ�E_Xͬ:Y��i�r�0�ս���"�>�?����ۤ���y�[��l���������*���u�f��b��~g
��X2�ۋ>[Cu\��*_������+��KE���{�����f�{f"���!�.<)���,��'Nz�,�F� |���������(��/�:]}y����	���}�'��P� �o��XuX:��]6jC���������Y=���-���g+!���6�3D{[TB����Vq�=�iXwޑm�Q�䛐����GO���.鐍�%��N�0��F�2}
��ьD�JD���:�H��I����bۛ�u��f)�؎��0J��=bo�m.P�?��)-8���p���n��̸y�fo(�̲���Yו�xg��i}9�����/��H�o��V+怛�E�J2#D���A�hv��7�0f H���eд�~Tǩwİ/�[����7�U]>�� `Yˣ|KHd�X��;Τ�\,$�`L͎O8yY����3�P;��Et���AGgl%�s A��H��(^�ZR�� >rR��ƧY���v��\,�E��Qh��z�3�?���`�T��C�y��_�h��<8�F�� Ⱦ�~��X��LO���s6��!���[X~�i��{<?d�}����?(�˟���i�%���^�@[z�!A��`���w n�}}�ݒӂ�O2=��:�꿱�b��{��N��?�s��q2_ʳF����coRE��@�%�Hc?��I����|!ԭ�Q|4���/Q��hP!�[5��ٌth1e��:��m�n��W�a?_f�Q��7i�zf?bY:p\��0~���-�c� 9��6ז�z��"�,�Z�
r]5/7a��4��3�a��!;p�W�õ͈�\Y.��~w��$-�gJ�a�euy�l�rɍ���	�\�]�`y���a~�Dm�}ݬ�%�u=����ײ@���������(_lT6Y�r�ݶ�rϘ' 5�Y�݋Y���ޢ���=W���'�T�[�rԸ�3�#�&���O���U�� |'���쬓@x�On�H�B{]�-�)��q��/5C���f6�#jώ�O���ﾣ2�R,�L�{�$	,�'Wm���P3�c��x��I)�ҬO��ZCl24/Bs��It7Q��Ho��
��O ���6���+u#�K�g��vpC�O�~���7��ӍE�'���4V��ӣ�;v=l��1�F�E$؇K���Q@)����[������1���Y���t��MjBa7���ݠ�_�������jP��8�+*
�\K���F�5o�~ZѳU��<�ʼ��$��9�B�1b�λ�v�Uu֦��ZN��+y�"`����[H�R�}ç8��¯޶�(DZ�u+�C�iE,"��E��u��w�U�X�t#�~>���޸�O���\����{�S=�� حw�Ӡ��]�_t��eD��5
L��VP��_��F&�2���BM:v�>-�������!��7~P�A�m%B!�h�|�Pቇ��/Y7p�i1�,G:��t�z����]��Y$����P��wM[a��ԪӦ{z����?Ҝ(�(�Q�zv��c�%��h����﹡B�N���O������n���0MA&7����	DH����B�*HI`��:�W}$t����K
�K# ��� ^�����u�޾񗊟W��Ɗ���(6��b�iN��O%��"��Ѓ<keK��#-���QÞ�q<�!7D���8VL�ɣ�ap��Q��I��;�(�6F�-����K��r��y��g��L.΍���������=4H�
�=�T ¬� W�
>�a�mJ���۸667�'�V�L����E7�8�X_��U�"��N�����ڇ78W������	��Z��J_&.`��J�l��Ա�k�C�������.��Fct���[�-�[$@A��I�t���j &<�f&��x�������{w;���?r�o�悢��r��5s+h'r:���m} y��_��=�B�g��=��Θ>��}��η���O���[����6�xIw
���lw".r� �v:����>°�\��ċ_���2���Y1Y����#[dG�g쫷�5$��-W��G��(�L������dC)y��v��kr��χ�ϲ/����`��T��Qb(?�zuq�8������X��mT��ɕ�y=O����%����^%.�A�j�G�/t�p��	E��9"�9�Y�Go�=�%� -���̀yv��2���]��
q�*dS���u�3(�,\��o`+�K�3��>\Ѓ�U��Gd�g�*�Q0K��H�R�)A5��y�>я��y/1�҇+-���!ğ��y��{�6l��VY+�!يy?��[��B��ԣ�.t/UT��]�t0=��:����f��<ێ��j�= ":�U��Ք�;�K(񽽜���	�y����i���*�����a��;K1��8�0K ���Oh�󚘷ϙ���N�
99鈷��F���ǝzqQ�~���M6fQ��X?�����Z�mu|i�H�R���8 �/{��Ѳ����w�"������]h��f�V+(��07Օ�u�����PKO��UOr���0�w�o9U�wY){a���"f\�	b�s�;���K��g�?n[�xU6�v΋<�Ü!����]}��-5Ѓv%zQ�Ƌ�W<�F��Ü �?�e�1y����5��P�P/�]���ݢI� m���[�uU�G"[�X>�pA�j
EZ+�4�D]�,dZ��R�i������"I���e ��d�[k%5�XAz��Y�B�+N?��@��;15�Jk���K�_�n��l�+jC���_QaY­���6=�h��#h�s.�r}`+҅᳈E �s��� �*�%h�
8_m��tsv �s�sY�	�tx2����HG��F�xt��9�� b5�IG�0ZԿ�t�[��gӼ�b}� �)�u�#vO=S*:�<%�>�vԻ6����Cp���M��C��9��:�,� ����y]�[<*^��9y1���5{�N0B:���Dl����jH�5��-�m��kJ��$^SĲϴZ�JA����j�z��	㵋���c���t!hL���|��c��V`�u횺�O�g���oX�����Ќ�[�_��M7Gp�m�~�\�T�\���H���E�8���D~�H�$N�П�|�V��u�z�ߪv�W0B�q�#X�eٵ��\qy�_�;�/3*�qf�"Ę_;bQ�]�� ��&�����A͔y�.�#4���fT浞Q��Cc�<�^�7�Y���m*hc�y�|e�����J�Fa��'�-���_��^KRn=���r��3�u ma϶B���33���eOH���*嚴#a��t��w���E_1���P�i	�YQ�`/&_�C'������?�u���P�6U�uv��s�/\��{�	�Dqj�u�w���w:�U 6���n�h�~��N�`;1���
���dJ/�Ԡ+��4���29J�\HH�q�k�e�P,��~�������2o8�3��I��«��//q�\!��io���i�����`��80wi�����`-g��p'A���Hk>uB�@���Б���������M��2��Qz E��LmT�z��Qlena�`l��PWs[Q����,�� �p�Kk�yNm�/Y�-1��������U԰#�^(Pn�M��86��s;���ݰDn|�o&\��>�.᚜�V�`���5�y�M���^�<���C�J*�r�I�e��ru-�n
	���3�N��Y�K�
�lexש]��G�X�[㛒�i����*�L#v�e��<���!����ae�
dQ|�+®G7�g�q#]\�ˎi��&V�?ݓl�q8m[�N8!g���-��VT���.%>p���p����m��u-�_Qp�4����l�~ⶣ�G~�/�������8��L�F���gR�_$0t�� �/谿�l~���v�P&�P���2U��S����K+C��ݽ>~�9�3�̐�9%D}A���������<����t���Jm��jb�>M����HJ	��/�B0Y�j"WŎ��ߟ�� peݙ�#���C�EeS�E	.*J��l�$�jߵ�c�l��B���n
���n���W�NPhu-�!%�r�0����)F"�=V5L�wxλ������l��G_��&Y̴�J�۩�+4� �A^�ʫz3�Շ�1=Ճ�Rl�iʊ!�I%2�	X��{q��Ŕ#4R�xlw�lq�RS�V7b��;~Y�!�����F� *r�:��s�8�Q#�'�/-O��*�3��o�:w�>�y�\9���jj��D���ǲ��)!���e�NOG��#�r��a"�mS��<���o�G�����3"�Ա�ԥ�7��ݝ�]���{tV�X�h�ҙ�N��u�QͰ@$|������������gj���+����!I�:��b5���_a�s����z'�t����<�9��"� \�i���f���ti�9P5u��="��} �����ߥ��/�>6�Q�y�9%7e*�
ը���ND:L)U_��k�����u5���G4�˯���$�����`k@���sw�Gǭ�\w?24Cg>-Pnɢ��|�ʟ�V�ې#|�)���3|�{I82\yc4={ʔ�XFW���]%��X Ѵ��'�䠪�2���u|>I��f����}��A.�uqf\&��{�vBN��G��y��~�U6~�ڲ��@�:��|g���aJes��N${5��ԓ���Q�dQ�]d��m��\{����C?�e0��+�ʝ,��(�@v�C�����FiNS�z���Ya��ꉢy��f6�[VgD,JJ&�?�m��Ǩޥ��i����4�3�����$�+��
��gT�p��E;���-�z�����km�@&C��
�A� ��ta��ڌ�ƈ	T��B���I�rk �(s��^�ٝ�����_�,z�ςyg����%F���@��a�%��m��'/Bg��9�LL�m��H���'�+�.��/�<����s���du�6<�+�0��2b�,�y<���j��&s�j��L��u���W���fУ�L�e%���'�n��΃���d�~�|����/��G/�eԭ/�(2EvAS��_�W������]��� �=�S�|<���X%��U����@��$�C���.]W�!s U�0�hZ:���j��
��p5M���%[ݑ���Q7ys�����h�P��Zf�(X���� e�`f`��t��A ȕ��r*�>�0T`�g(}��`��	��."#�� s���mQ��L���P%T�j]J�^E���k�EF#��݁,� P#?0r�-�f�_��79�*9�ې��#�̱�\55K�B�����Y�A�٢;��Hr͙�9J@v�b��@ A)�́�2є�<�nR���N�~ҵ�%���1����j�@t+�\
�rG��6�uc��J�@1��o��Dܞ�8,r���?q!�MN,�
�1ac����G�Ǫ�?�W|�{۹z�[aT`
�D�	��;�dó�t���@{��sG�x�
���\K�l��z_!ִp]mE5C�p�dЬ`}3��U�L��4�2V[�_��b��H���=9N,C�f1���ug3cWyɪ��il����Q,�1$��.>��oT܃�^NL2I�C�iT�`}G�l�6x��Хq%�Ɵ���	I�	M$Y�+�b(�i�b��^��	��Ĺ��Du֬�c.�NZڨ�ɑv#P�W֕ﾟ�
���:��s��L22��Z]j����'�x�F��Α����.w�94�Y�����aH�`*)w���
���b��R��\��nd.H���8�I���C��k�v�tc���Fߨ�:�/�zD�j�/A�[�%1��oT��i��k`��$Т%�cI6��(B�i}v�1,������c��9��%�����x�1(�10?����mL�����H�ɡ�8h����
�X#���b�b'����m���Z��`,Y�%V��c�Wy_��`O}��a�M��d�wL;m�z'��X�8��s���U�KGDF��}@?nb�·kzy|�Sŷ��@��@���a��v���~ڱ����r�f�ެࣻ^�ˠfn�@��")��c�neuP	[29�( r�AXe�Pn�f�&�$u%�<ʻ@3O���;B�)��n�t��Yr��d�S_7�k]�!n��x�(�_^�/�n�R�Ld1��B�cx�����eRC�Q^ m9�j~� �dpQ�@�RaYi�밯E1��Ⱛ��$�>)���s����-�Ǯ� �W��Cu����ͽ�7�	]YL���3���A|,�醛%��h�&�& `
�%^�o�Q�����k{�ѫ�l�Բ?���^ ���X�~�%���]�x���$��%k�������D.�h��{`�v�	�;j�o�:S�?�'�����Ic̹��qZ���"�B�d���m���Q�-_*P|90��R�urLs�
��������
�H�2v�@@2#�0
!I\.�@0�us���O�](N�u�D�)�;�th�2��?��g�i|�7J������ � ��K�J]�o�=Op�?�dX�A:�#sT�	��Av��E��^
vV]J�Tk=��۵����b���(�r�+¹Fٺ��aB�Ѽ�`uז�W�O��s�Χ
Y�����h|�aUhPq�\Un�����T,?e�2װ	�D����!��o���-��c�Ns�z�&����[�-P�vK��P8��V2�͉�*[�
sI�__q����1gSV������U���W�F�#y@�6'��8�~f��Q8t�ŏD~��W�}z�XV��j��Twz��l#�U�����|E"1��[�!$_��vP`�}i=x�L�d��X��0c8�������t.�Ћ��O#hb���Z���4H��{��u�0������+�I�
$��*
������@��)g�����7%d��Dy��l��j�� o���Wh��P�u�������t����h5�K�L�7�����uQ��i�1���D#�E_��h�T"��홫)�t:F(w\�~?z�q�CI�5���hƮ�6�F���d����d%��q��<�2�j��� *�Oe�`�Y{R e7
y�e�[����	�zl-�+�^.O����]����P�� ��n�EfU$M�pq���v��������%��#�������p*o �Iӱa�4��J*�e�d�~��4[�Y����Z�}q����6�E�$�\�2:-q�����5��er��zZs����e��9�|�cj��?Ϡ�2�x�m��\S��w�}�4�&��֠  ����G�ע���eүV��-=@q�����?�X��A9�ľ#�Um["�Q���I��/��I?��[( ��
�;M��7N���'eL�u�_�`��������އ�?4[�[�R=>�w�W��~��duer�;X���@��=���D<���'������zO�M�xG�*��M�&���n2B�}���N�~x�i�,�d5�:�Y]�6��`��#8tv R��6�/��4�Ӓd�i�2>�Gfbvh�ѷ��1�E�y���6\�5:�QgI^�Ӂ0奰B��@��"sW�G�a�a��lu�#�x7��C����eg�o��\�AO�*J��#X���AX[�y;S�\紊��rel�^���̷ba(�l�	���x%�n���l���JaJ���=m>�.:�c!���1�#6DV`��MG���zlۉ�	e�ȇ����6;�*�E�i�1^�/W�qm�*�����4ˊ��Ų���T�X���j�oU:v�����!fl@�.��d5ET`�rܭC���ѵ0A_Y�x �6߾Ϝ��搀V�b�7Ɇ�����ˆ����Ɠ���oF���0�6L+����:	(YFI�ѽ�m\U>��Ku"�b:Y�.)?3Ύ,�Ey��E�={�{͹Q��FG����N��6G���I8p톓�5�IT��Uy���R��D�����N|mMqy.C�Or����0���zH2Ut��ƛ���!��D1���#�&����I9G��$��J��baJf���A��;Sp���~i��̉��JS���"TN��2ѹ�1�����&`�Ģ��C�!#O�`]����'���G�C�"6�3�~��*ɛ��� �\y�Tǎ�[�KLg���x����_β�=�^���>:�MB����tKH�D�7�p�V ��Z+���G��g�S�oP�H���iK]<�l�$v>���{4���ۇ�C�eU滤צ Y�����N-K���V�/��7#-L��
 ��aM��c��s��I�#�#�ÆD�s�<�D��z{��M�����'�S���(������8�y�B��o$�Ai�W�v�V�f�:�aw?]x��$Rz�Q���j��#u?N�P�j,�T(kfuF�#o��ل�4]����g��g��H�h�+��m6����1&t���Vl=�j3��Y��?��Q�����ރ.�� ���|B�aro�}�i=Ҿ�"�2�f��c@V�-%ߕW�z�V�eD񍛯E�Z-��By�7�
@MKߩ�s��=�/�����������o>}v��/�N	�q.��qǶ��Y����/F�C��j���_����10!�dw[?[y�q도A��b�,�Y*{��?ǒ��M�������i��+��I�s/��XH���se�m��g�ȍ	��[�IB�&�Q�B���K~���g�����������EP���)���TU�w��Mח�J��BV�$ 6 ��Y�0d�[�C?N��B�X�qT���j{�WWWB��j(�b� ��~sm+9� �W+��m�O��@��v%���=؇ -Yԥ3�t%��A�A���݁�E8�"k��L�I���%o�I\�s7���5Zw<�c�x��yp����no�wg>Sً_���Ul����n�#�Fr��"Us7�'�h.}&ѹl5;v�<��?mK�z�v���z@bD�3����pn�PMPƊ~}�	��ӾA����ξ�\� ��#��T��%X|��V1�H;Ox�R����5ʩ�E9H!yx�����z}x[^^����4��<�nrgkҩ��Z+7���{��	�K�*�?��o�Xʞ�G͵���`Ôj��;0�8����4Fof=S��yEl���oa��r� ����Yߟ $V�{�%���s$��
U�
ؽ�6��+Q"~�PKe�9�s5�O?o@!�2��8~Ŋ�?���|y���W7�����&��f[P��O��οW
몧A�1Z�{!k�j	)���I��N��VO����v�+
�3�,j�7G�m�F�p��4Nw�����aoSN#��
�klf�������V��^h�����c�M�@��o��&s�/ �W��(�x2e����]�e�����%�߂�f����b�E�$��-���d��ϱuf��gdg��g=GK�T,k��-Y�Fx�'*��QK���,�3ho�H�y��Ӷ�f���<q���{;�<��#���	l�8�zR"��|r`'ܶ	�h�1b���!cU�yF�r�"����%[#��dc�CP)ÜE�d��(i�<G�Ф�h@g�tɳT9~��	���Q|��q!�Av��C,g��W��{�=�'?�3?��3������+z9{t�B7d5�ť�e��X��Bc|���g��>k�E��Ûo/�#����E:N���[=��,v`D��$��n�v�p����GX��ĕ�`�cb�ɡ�s�0\���F��
��>��d�㭣��cR\)��(��,%P��d�RA���(Ɨ�+&ma�$:������S��!���O��N�r����<�&�P���P%�j�f��,
l��*��)����~,��G�o�:�Km���e�Hɑ�p�U��!B$�K��\fJ�,^��n6g x�/�q�@���s#� yJ�?�̚I L~\��3MZ�p����ϓ��=W��*#�AFS��̗��$�xm�����+i��m���r���Y`��P�n�L�^I5�G
Q��6X�����li|[�]�;%tI2N"2�pi�;�y�:��0���g<���)P;�C���U�0p���&�i��+p]k2�Nn_�D�rw=��s��6�\S-��u|nL��eۙ��I�$D��D��qD�P)�M$�@e�����Z؝�m����]JO��o��P�
��]�#�ʌ�(N����^V��~lB�}`#��jG���3'�[�'z]�Mw���xМ��g�v[K��iw�G�s,=���⥗$i���BX!HFm\=�N�5$�z��_����B�t35���V���0�?_W�������W����f?���)��g�C��#����8�z���ǥ�Qt����81�m-6M�TdZCC�f�^<�Y�t�O�#�lI��b��i�{�Y)����)'t�̙`�"nÚ�w٘��I ������LC2B�Vշ5���׵�7�d�-*Թ֫��*��������Ț*��p�f�3R�-�2��y<�YXfad�� M�9�<�sj��b]݁1i<�s �{�6[�����"��_d�lqQ<�\���~d(�csƲ o�^����f��)�50�$�&g�	������w1��>Ł�������ܪ`ca��&��g\��"+�L�+�P8��\�̥��J�t�aـ�λ�&��+���%�Ԉq0�C�_fn�t:^�(�m�D�NY�U�IpyZ�P��T�>K󆄞v������3�O�7lS19��4g6`��Ǡg�[���N��O�cK�j{��b��W9)��ܨn�&f�S�Q{��%���������î�2$�;�-�܉���.��H����[\����lŦQQU>�aÂ���i�d�;�>���_����?`�KG$I��cò��aW�|M^�+�?�}�5��P���N���[�Z�2�v�֒��=7�=�@������K��H80{Wѹ1�Gf0�t��Z�(�f@��ᝥR�By�{/ȥ	�q�Q�!��eЀ�5�?�Ľx�d��ϣ��*�[����,37�orE�����U<ˎ�ٽ�I�s8F[�~:�U�/�ԑ���� 6`�-���'k������+����"��κV�eO3��e�p�J�߃K�.�'�7�h����@D�W�b9����=���X��������W��\��N������P{�BQ�xK@�)4<�'m9��ҳ�Ű�M#k�V���'e󝗧'v���m[���!*ݧbxx�u�ܾ�&w��?F�(����EҌ$5��L�o�Ê����z#"�F�~�W�o���L�Y����Zր)�
i8��~T�z6���H���ҟ)L�^6v1�Ш&�Cu���g~�JFn@҃�G���L�1���6�O4��U4ǒ���ƞ�,��ZO�EΩ�u)dn/Nc#@ȱ���@�>�E�
C�p�����Ō��⬞S ܻ�A�l���[֙���ȶ�����A���5�sn��P;�ߨ<LI6�۰
}q����WE/3b���S.
�\���G�dG,!�?���$ ����o�N�H���J��4bj�S;���n��E˸���	~�]�j���7��If����wxM��ƙ�r^]�F��%*?�_�X�3�����7��uP�������cc0��"��[�VJӧo`F��F���?�;�§ֺ89�M0K���Or�$�.6q��<�I��?�����E"j
Kư]��I����a�#&�!��C�u�,C�R9�M��;�7�o�N�>NG�/��^X)�:wq�	ؙB�����<�4�+W�_��%��?�1x�5˧L�Y�j���U�����t�D����U黟��=���%���S\�/�~�ćLvƸؚ���>I�@v�y�|0���h�Ĳ�WG'_Ei�����:�ۄ��?��¦�&�>ĄD6���� ӝf�)w��ۉ$����gPJo"�WODB��hH'4���Ӻ�@L�=f�[H$�g&F5�A����E�l����o��c��(yY3��;L�e����NvH�iH���������@r��S�����g�L��Q��p(�g�A`�CGh�¢���4�dl0r�هЍ-��#:+��7v��Ny�̠�@��ade��r�ϻ>�(�0Dӟ�xAH�&�	��L�6�X�g����:��M�z�����׶��:K.Õ�6k)9�����H-N�}���(�B+�0E'Qێў(}�G�`┲���VEz��W����w��Hke,C'�x(�05��U�"�
Q��p�b\A^�ާ�z��~x�&C�W��TO�j�l�ܯCT�
�4���>���,�����T�Mr6�	㍱����e*��f34�����l�(�m��Y6wgm��W��f�Ӛ��h��~س9�=`Q�xɂ^��#��'��k��'j������n�m0��j�8�&���
�/ݙ	PK��D�吨Z����0"0�Y���ʰA4zloTd�7��D�w%���ބ�d�9��;������Y�¶fp�`�?��i���G���,!�gȞ��[��zoZ�?�'Za���;	��)�({�����v���c!��� K+"�!��b���Љ����z_p��#���y����`�I��,��v��hI�6P��'.;d� ��u�w�-G� ��wH��ϣz��������?�1������m�w�̳STG� e��*��)#$�
��č$�6���ʍN'	��/�"}��]N�p�\���q��C1��KS�F�}EO���GO��ۧ��H�Ɠ����`9������o��-�fB�4�b�
�أ�h "�5It�/�u��ή�v���U��v��%�U'�^�m?_�1�ZF�&f!�b+U���
���H�]h�Po]L���#ι[˫�*D��s��T�@�{��aAv2��?*��JXQ#�E_�)_���^� �A)D�H����Ŗ���e�W/�6����2k��F���!Q7> �f�� X�f	Vg�5V/`<��~���Wk(0$�xC��x�:�<��'' k����O��*�Qo���SO�DG�r�^t��U'�,�f$��$�l��	�GIX�ѕ|����	���C������yG�hi/� dr%Y4�+b��W�GW�,���J�#v��0�'���r� )8Xu��NL#���3�?7�X�2����y�����U��/�^�hc��_Β�Rt-_�_Y*%)c�a M��P�T{y�ҝ:����I�]�S��
��M�vE����!(�'N�F� ҃ۏ�\�}5(/b8�7s��t<2è����O�|�\�7x5:�>)�<��Q���`왞�tO��ǰ8:���,�^W�%SL�`O�K�Ȥ
����'4�5}����dmz�X�`��'p�|`=_x�K�k}(!��i� �2,�ǂ�W�{��ݡ��	&��������婪�W��f�R!R.�1T%!���&2��n�#���P%�[���&��UJݼ�hs&�Ѯj$㣎�i)�=�0�����?@���m�Z� R�Qz���_�)p`s��sh���ŷ?K�5�)�M&E�� )-W_��+���1�$%W~�_�RMGbD��,�E�FczA^�mF.O����W���U&f� 9f:Rȗ�x)��3�8����R�ˣ��d�j/f�f���R[���� '�|5�}�=����7�.x��Kn#gT��a��E��	�� ���:Y�����jPs&c��S�P�>%֝d �Z�\ x�,�����'9.WƩAy�&��y�r��^�LfX1}�� ����a�7��z�̓�u�_U�7gF�pҕ������I*���Q�ƄJZ�T|��r����kk�R@�Rԛ.e2�����-�J�gÊ��F�c߫�vγ���9�W�Q�W�1v�@�Տ�x��5�����6��ߣ�t��!�?R���:1�x[�/�sAmg����/g��q��2�]Kv�1��O�5������O���+�
Ԑ��wu;��\+����8A ��}-�K6���[i�;<���M��5~$ұ'��©�p2��
��ߕ�p�ʄ���q&���uE_���_��ȒN��q��*8�s
��D���E���~ms+�����6���ҥ��gf�oLR��Ȕ��r����)����Ĥ��V�`<W��s\g��F��[�1Tݚ�����y�H���*�س^t�*R��>e��%P]oL<�I���܀cG�q��s�y�;�����[������[{� �Ǯ
�b�$���1��'֣��À��wn�����d	�Z�Ҙ~���'Ya ���**��wp*�ۂ���-T�ǈ&��v1�ʎz���WQ�̝��TW���j�[��Kb�����Ku� ��
�K?$e^]�l��t-�R�}��.�W����g�Sڷ���[�e��b0���/^X=[0��T����O+��t ��^G���u���hEk����_�{6��'l���Hc��2�T�P�8���P��?�'���Cpjk���ӉF׷��[`4��b#t;J&��S��f[�2�P@kb�g�>���EN"s��O�`kD�J�گe�]9>�s��^5FJ�64�I���P�B:�sҞ�Cq��u���/W�c�@�c�~֣�T/���azo#�5���k<���,��LY�~�8fl���W{��>+�~9Eqw�A:a�n��۵��z�V�p�<R+V�|X�m��{�ꏱR�e�W��ȼ�D����$�@�*i���EW�:y��k6�U��\�}(,����(?�%�N�#�a�7�ҟкA�Q�.ku%���(z󻊎�%���F�����	&�k�l��V��)�0����2ܿ��{�	���\�ϴn��O:g�����˂�|-��*�-oHW�"��zS��b&�Ӟ<�a�@�{�4k,��=e!oaX�Dx�5\��PkH �3Ȼ@6��V���B�\]G�.M��y��LX��l�ݴ�Çw;�Z2�8eo�3���	%\��ǫ��H�f�z�zQ�$�>�&��R��y�ț)�	ۅ���?f�� {B[v�^k�� (gX�e>�"=u�|�T�'Q8tEz�V��s�(����1��g+���Dc:�{^��u�`�FTw�c<���x�]�E�`�9�W0��J�m{T��:'A'y^�kn>A��=�I�(܂����~Ð�R�������6�c�q�]�M��Ҙ�p�b����;r#S���M2��z��e㐳����d^8BW���}��c��R�T��C��Wf����k)��q",���B��@0���.��"��؇f�M_��؋Ǡv���)�Ӎw!�[ef@ �b��T�	�ݩ1�%q`ыj���rHZҙ��۶��X�3���ͅ`�@X�s$�şeIT� '|�a�K^"���u�\�����W�Q
%57닺=����7
�84{�~C�{���z�k_���
>_4Q��R|�uH'����Ұt'������"���J�9��{-�m���(�@��/����ּj[�<�75��0�OM�L%&���Z�����=UQ�� �˿x��e0�__bY�n�i-��d�����h���	�m���*/B�hK̗QGc��Xw��DtX�������w��z����Sn��-��%@�>h�b��'�)?O�Qc9�J�Y��ǧ����d�2�,��y�E�	��sO/�*2"zE�|.M;Fs�қ�K4���|UlL�}Ez߼��ؑ"D�.M���y��x�Y`�ӚݛT<��MEM��Pt����N�,�P�5�Ī8�Z���T�����j
�#�r�� �����:w�Bʇ�(	&���LxT�q�a
�*��썏3h0�;��#�2V����xzn[�1�z P��Xw=x��Ĺ����5�^Y� r�_KH�'ȕp�*Y�!Z>��3���ຈ�Fn����XN�C�pґʏ�d9��`bt����~��c/��%��E�E}�.�O ��p�]>�+�{��=&I�U��)���S/"5f.ڮ�-�Q�F=P��Ǵri��t-�)�������4�GXn�xx��Y�U0[��i�:SCA�2F�8l�V�C}���a���+v��rIZ�=�I	ш�5�u\�0�a�:P�#�y�侥m_��q���XC�-�c�U��E+�[̲u�?�xC޹�Wm������8%�/�'({����r���#��~<��:�1�n����3�A��`�b>������7]V��1z$��{6��r�^���\��ʹ����	
K��Z�c�L����~��W�]ʑΡ���7�"��kBU����#9N�q��]߿�fU5�)�y UH��)�2��R���8������c��;�tr�%���"�G�����3J`.q�w(%������0*Əe�-I�:�]���]�B�G,ۦ!3
�#��׳�Ċ�Q� �<8��������I���cb^'Ly�w\ƸTQ`��m��@�k��/�	$��Z�L紬>�c�cN�����V�/9�G��*0�`Ŭz��*�?7��7��������w�/�L���UKQ���+z+��a�
\X9m.S*���%�Aa���=��-�a9:�`T����i��-��[�ף�3�2�-3�nPf(a``O��
*�NpCL�mc��:�V��V�Zn���[OP	Q*��
��I���`�nHt2R��^�b$U��|�=%�џ��x��y�V,_�A�q�a_�������D�"���]0�}�&D�9У��g�t�F����Z�@.ZT��͉.��Y:�\~�o�������#�g��ӊ�2Ҕ����ԔoF�f���苰!kD�a�;�&cd��b����MD����6�0�I�*:�?w��%!�<L�>�{����;h���q��QX�g�Y�)b"��b���3�ӪO����*h��q���N�"׬�4�����z���$�+���;`A�3��aR ����}����猑O�	MbV�ȃ�>�W�
<���S��x����;�����7��p�Ky� �R=V��&������>��0�)E<�i̼3�w�2�����=�ˤs�T�x�k��7�˅���j�o��C]Yf�?�5
�h��ъ5�b:Ɂ}�p�^��z�#�g{ȩ�h����Ř�]�Pc�W�IR{({��,d��h��4��[^&�#�1���6�=��˅^���zp�l$��3�$�Y�WQ��H/$�H`O�	�rݖM�����J��N?Ԫc��N����4F�?�_�F�����q�˸���I*|'l���N�0���z�d�r� $����u�`QYk�*��u��9[��XMg�tJ�<J�jEQ�&�>֯õ=�[���ƃ��-�ݵ|��JY��k+];��b�@AS��i/"���@K��r����<70z��^��I0�C��'���H��_,�IL������b/�b��H�?����~ �QaۈK�n��4ȏ��?���Y�"
h����̮�C�X�#ƻ�	i?&v̾�����X��a�|�����$BK�	���:�7�6�f$���&��Q��[�ϲ�kE�dԮi�W�DZ>�#�"��.�0vO\t1Һ�f�݆�&;��:lq��ˆ�E��N̞�m�WiW������Yeh��I������d����o��w���-3�fgS�A;�>�<p���~�=]�yfL_�<9ݗ�Y
F�`�����|��62��m#��͔���q���CK��jqs�Y�a�����W#<�UM��M��0���yX��x�Ae��KbeI+)�����N~���]7�~�Ѳ�"\H���]�ݣ��D�K���k!����"��,x?�7�aљ]n�0�tn[��w�b?2}1�w
l@���4��(�3=��֜/�1ļ扑���w��eV,h�YR���. L�F���j��sh`xf�{��-�]�2��ͼ�O�^ie�*a[��B��#���ئ��k$�G+e�#���*�t�܀�4�1�_
V"v�c��4C�_Mև��q���#Y�X�� ���� ���t�2�p�4A;F
m��u3����gma:�i\�ɗrF�{�Г�A怑S���� ���Ya��~�wpjI��I?��;��
@TUGpG䩸���;}�ށ|&u5L���b����׮!.~�^�p�~�G�㕎���D+�3���`=�y&�_$�9��N�Ї=�TR���f�˄���S]��H���<;6#��#S*�%��{KFnw涩]�P`��Y��l�s׶o� �^;:�%u�ڈz�tJY��s/��wȿ£���BT�l����/u)m>�"�~+�l�ҎM�#�V���O�"�����3�䫈}��u�UɆlG�V�H	��{�7t�]�~cGC#���o�S�
h��@1�>!��<s��X>��JF�Kz�N8������j��^��eGo��F�?�U<�"�	�H_�¡��p�K�P��l��s�#��/�*a/��0�����3�rC��k� mi�'��%Ĺ�v�WtY2N�7,>}"\�1J��ɠ��B^�vύ/�ʉd��U�*�rEU��͈�T�muuW\Mu�,�E��R�n�t[n@��Ib�E���W��>#Ó�kl�&���/vs��RH��d�|=�P�7�����=J�E�8������?��	Eԫ�ᘎ"�(p�4Rd�{}��x\�#��$�U�(>����)j��]�"���팚K����{�c¾����/2c9u�%�8�$�F��?i�<L���L����?���~�N(��n�v_���I��
 �5K��-�Ux}��>��&>˂�2�>;h�0�!u�]�� �J$K�,? �(A,�#��j�L*�_�n�CiӔ��d�Agq�3�)F]�C���!g{�'n����Y���y<�rbϰ��!�|���9dy�&,��;ý�	�m��
����lȟgnH�IA8/���	oU���\��i�}P#ULo.Ʉ��R�* �DI6̑��;��]7C�[m���tF�m�B�#Ze�]{�Ob|06��cb#x��Ұ>=�71���?���Of{������u����K֭2�?��0WFI ��eԳ=wZ��6 ��%�z�;����?ޓ�VS-���n��>j�������F�h�?��Zz�M��U,Κ,�-+8݌ch��S��T$S���͗��?6�T�M+����D�n�NX�H��v%1�ap���/Þ�
�y��"}�¡�p�Y<Rezٯ��Ty豨��}���AO������˃�}��+`F���[>nJ��E8��6 �1_P�rs�����ؾ�ćs��|��a�܊���C�b	�Oz��6P&�_�m`:
���%޺-X��R1����3�={Y8ƺ��ٶ5��E�P߭�F����-K��*l��t��+*$�R�g���w8�Њ��枖�.�G'e�z��}!�h�{Q�R��^�W�1DE������G�����5)CB0&g�ܿ"���#�)5��h�r���D
�[,ms���*�K�x{��-#�?^L�ɽd�w���CCkܷ�/��ȸ����b8����W�%+�eSR����Y�:r��z ۀ�W���l���2�Z���kc��m/�v[>2�<��|�`n��C�i���46�6��l\Ӄ�&tI��
9�$�Sۖ�ۘ,�ܟ�7hB;7]��B���d�I���Uwǚ��R��pܼdd��&uY�E��Q~�?�E������I"�؂M[i�J�X
�s	$�_�-�����.K�P]~���J=�zwp�<�w����$�%3�Q���n��_�4@�}�Ī�����Pܲ�as �6lsyzjeƆG�xT��I%elZ��?����т���_��}h�̫��bT�}�W��'�^M�5He�˹|޺FsZm�ޭy:���Z'��!��"�r�ș���LS�Sp��C�H*�7DAƻam�߾'|)Mt��+��� ;��×ᠻ��ڶz,�6��߲�s��/Y�P�:�"�eR.Y@ݮ�ق\fe1��U�b����K��X�cg�ӎ��-�U�i-�έ��{��E3[{�O*�^�����.�g5.F�=���4�)q�B�z�e�C�X���˖bl�%&�'�)�?*,V2�����~�=A��Ǎ8�����U��ꩱ�m#h/Hgx,[B{�]�Hr���A�c�ŝҐ*S�ù��3Ć����D��S��	r�W�;s�ng;���(����P���1� I���( a�/Z*Ya^�J"�L��|�_tKȪbd�_@鰊xL4�)*�
d&�=^���MۆH�j'PNd�h�q��%��m��:=�|PڰvFGM�4��Sӣ��H`���>�cX�|!��˒�0�qh��XC�����NH�}��Y�m�Ǔ�o�j�,X�R�6���#Lg�]��]�l�Z�Z3����@�j.�\ N����&o}]�������0-�텻К��@&&G+F������1�{y�B��4:�DMQ�����&8ϓ8uLk:�&�eO�Y�������=�H�H2&"N�T�����ݛOQ97ۘ���H�V(GA�DE��`�*Q�O/Q�s����a���Ql�"P� �q��=(���^���G���o��9���@m�����]�b��ض�gBGUO.Z�A}ިF��!3�z�'��C㊑���ϗe_Mf#A�C�i_#ݓ	��ƥaŖ��I��5s��&�O⑦ YW�A*��6K�h�-$��;�	��cj���{�Tk>xf�� �!�*�z�0��� �6�|-G��.ƈ�%�mW��H���įB"L#*v�� �/[5h"n2#F�h�6�Cunjt�X}N'�{Q�����^�.��g���r�[�I �@��>s�復V�?�k��w&�?�ف���'oߡ<
�ac��x�&ذ��x��H8*`��Yވ���vŘ�^����誜����?9I;��KΙ�K�&<�A�,�=�ƈ�3dOj?d��d��|�t[���R����g�1�8x܅51�@D?
$E�2�	� 7�տp��W���w'D�Ǻ��%�u?E�f���DB�A�TW:��C�]��)#vZ^� ��3\Cei���N������Iҁc�Y.\QV�79���Bפ,K5�rUO]�������΍ ��+������ۓ�\PX���ik�l��lC�����-�E�K��K�S��"Vǻ��`Y��c���mp(�`��5?������f�Ezǽ�`N��[_j�P��`�~��� �j�{�9Cf�nq �6�]��j��p�fd���`2���ؐՑ�Y����87����� �8��g���!�6A�"�:&��,�S�99Ț:���.ɟ���Oi*���ά�,,2��zl��c>�;Yc�8��0��g���Ґ�Ç��w7w�0�1����R,�V,]�ɦ�ES���yʕy��Y5�Ӓ�Gmr/��e!O�h6o
���鈕Ф�#k�cO��6Ϳe:0��|�#./�1�T�~zWN٘rDn�
÷���׫R�/�q%r�T�
eКQ�|�UZOt�O����ϖ��O>� �Y������7ٲ�ul�M�.���j����9����H��h����~��D�b�`7e��\�2��M	V8�R�v�����S1!�0]�!�R��O��@�V�.�y�t���@�BV�'n�G�n�)��z��cEq���\Пͦ(�$��h#�9�(�ʄ�C�&���=K�lr�ً�lp\� ����ޯ>t�k˅A�SAj9Z= �X�Ա�b�w�<��-�+p�N^mX�S����;���	����T��é���~)/��H������E��#= �_fҲ�k_�%H.Wd�o�����d��ocj�E�=���Pv��L�>��X�ce��2��d����iǳ�B�����Pi���zғӵ7�~�ծ��~�:6o<Z�.�%�Jbe�}f�RqtU�G�k^���M��q$)J� !���J]�|18�K"�{��^I�.�J4	���.�:O	���1à>ȫ�F9�	$��i��P>�j�f�pW�0�gv�I ��wj.0���#1��9��g�&ZR+��s��V�̈>���s�k��M �� 
NI��7��8stu(	"��F6u��bM��G�C�1l��k�{>���P����&�����٧�ЩM�蜋�����!��:��Y��"��m���X��u��AD��G��t`%֠Mʰ��s��w����=a�J�}
1hb�'���~E�����9l����Ho��cn�pJZ�ި��K���>n�%��8��2�%�����N��@^r��r�>�xC�H��ٮw?ۨ�m��ր!}���~�j���p��_n�q:�Fr(��3�	0.�W�Y��v)d��,�iV5�˪\s>��1���%���͍&�1����u:��kx �2�+M�R#?�<�]�t����
yL���Ѣd�p���0GƲ7�=И�"�L�"��݈���-$�����֘?���������2lE}���:x��!�EZ6O�X�����^�P?�ߔ	���!|P/�C���œ��'���v�ny�)�[cO�q��Z*6� ��y�o?"�r�D�kݛ�F��X3J]����F�J�0�<�j�m:#\L��l���F�Fe~��')C É�h����M����%�V�����y:(|������O���wc�#�< ^����Kv+�z��7m�Mö�NŰ� Z0��d�dU���:V�i.��{�ŗ�u\�?��ǻxu�W��E���Z��N�l����1�G�,�g)�l�Nn��YVU�w��B�IM�H������:5ָ#"�%�'��+�l����Y�A�
1��Kv�+_�AlQ��ƇTl�;y������}�����_�N�=��w i���"�U�
������:�+-C��@����)�˗*��_ʝ39��|@n��B���}L	R?�~�FQp�s*�O16��y����ߋ)�W�R�<�S�����_ �m��Ӎ���|�o�W��xu�s4s�E��ڎo�c>�����;�Q�!����1��K��������â���NK�z+}�����\:� ,o��f��?��gN�M���fl
����P����c�&�x�л	Ζ>?6&0_꼲��
�K�㶹�:����}��>Z��"�� ��
�i��Hǖ��:VA��q��.���si��忒ѩg�8ɫa�!>��Ӷz�[d "�X,�`���F�^�TNÙ��22K4m��:+��� 	����r�~Aa�bY��{���7jp�b�R\����<��>��U�������ES���/}t��yQc�e3�����/}*g;���M����A���G����� �b��u>�/{􀷉n���&�W=�6�0�D�n\�����S�Ј1�F�o&P�q�6!vش�A�9�#BB�;��V���:y��$��2�M1�.��h٭�z!ag]�IMY֯�r4�v	.foZ*��������4���Ê����6�����2���gq>9%�o��}\뉫����]��E{�C]����Z��`���0}��+%q�Ni%��ŐT~�d $ﳺ��Y�o�z��_��K�uC�4�弢:�d�M@
T�P#U/�����{�C?�� ��:mE(�D]�� �Q��q0Lb������;�,?��1%hXv7����O�u��GnO�������X��C_�{#�E�� }�I 핔189�i��*��gbu��
a�d�F�m0�n��V�L���`�95��Db�n��,c4�w�*�)��=}�lQ43%B3�԰��Ѓ �l����ţk*g�:9��Ӄ���#ϊJ�@�*���j�!]	i�]r�(����4��~�����l(�.���?y������ӎ�ԧ��G<��l��tv"D��LxΝ��21�l�0׉3,�8k)��Y�zB�� �b�������E�v�y��+dA���,}X}R�J�)Ktݢ�=�mc3�x�|�]�B�}��n~��Eࡡ3�
�fm��JΝE,|����n�Ww��:ϩc�ƻ��&�\����#��<O���
��������rV���Cg'�]h@�F>C�Rpy��MW���f���
f̆|�*9�{4#.o�d;Jc�û*)e7J����[�ו�(�e`�V}�Gqx�o�=��fi��uxn}[a3�X��_ѣB�	F6#�.���6�����g�[���dͧkoʰ݉I�΁C��u��z�95��泜��E�Go*fj�/��z0��a���-9�L\E�fn�N��&�_��6lB'�6
���Hk<�z��&<b�l����|͖Wy�W��3�n�����NB33g��$ٓ��Qe�4���)�r��x4�&F�Q:��R{�wSY
j�C�m��RS���6@izϫUw����s���d��քڹ�OS�AIr���m��ِ_0�5�$�/;��Kfk�$<�����(�^�#�^��ܬ(��'�@����=��3W�M��rhQ�QZ������5B�05%vq�F�z�ƺ}��MET� ��¤7�Tk����%(�J`l���r�n�;�F�*]�O��f�i!�ݢ�}�@���U�1��?�}�;R�帷Y��G���v �T�I�ִU7WJ�9?C��)5d����
��y�I<�x'�X�H�vAR���zױ��#���ɛ��%`�wcq�-��
c9�,�3�R�B�� �z!�B�2� u7Y���j��d��7��p�s*����AS�!��~��Q�+Qϙg��}�	'�.J�e�C�.����B�:ХR�W���Ff��*y�ί���r�!��WZ�^�ӌ(=(�I3 '�bO��>�]Ufza>7�Y����|����8#��n���ɨR���bt�vo[��Z����Jdw����q���Ms��Sp��������J�V�]'�r�5�KZ�.�l�04<s����b����8��!�+�Apm�f*�BGT]�����SL2Nrqs��>>�#�璏j�HȄP�
����ɮ�;���n��T{W�5V6�#IH\1JI���c��RKsfnN��]j�|b��y�D��F�t�P�^��"�g����}���=�ֱ����A6��oWA�I����]G<�� wu�PI�_���	c�"��������b���aWD=��r�qMd�����䶃�xA^�a3����"��k����ڣ�;j:3���t��+�`)�HZ�6<8�Jb&&�w�pΊp����7�}����iS�9�OX� ,À�!~�o>��X�:>�:Ǣ0�H�!b��C�z�t�J[�~Q�*V���N'���Or˴�y�pQ����B�t�|��ʳ�a���j-2�늒n[d7��U�9�ڬo�D+5�χ���aI� �qp��jp~5֩��Ck��U��3=���IjMq�N�ݥ�5�
�a]5��O�V�Ӏ#�ݺ�� Һ�^�k݉�'�<�2�҄���ꕰ�J���K�:7��N\ �#Q�nl�|���ox|�	�D3���5a��|h/��Q�X.-������`�!
9����6N��1OA���K��Pi����5p��NjR`��Nԉ� ���^�9��"c��;�+���F�ߓgO�F��iW���'7����[ٖ$v[�����u%Yu�ƝU�^��x�����/���P��]��]l���^Х-���!�t���!�]��/���?����J�y��޻d�#YEB }�0��,�o��ihۢ�Q*{��Q-zڧ]��>�����2��eg��# ���d��.9���9��V�ur�Ŀ(Z�qăIN71<j�s���� aCCSA���$>q�
��h���vd_:�~YAJTk�_�[�C�bׄ�ۣ7�ˊ�Q���}D6��[`f]�(��(')��'�Ț:z"�(��g�V�2k�&�5'��J�v��w܃T7uט�j8r*CB'_R�L� �!��J�4C��P�k������d��^����k�8�ral�tM�>��ܗ)�,�`�#4���� �� �c��j�.�(��_E���Π���J�,�Z��~�\��Qx�ÁZ�86;$�#3�/�8K0i,�-������I�R`y<\��dL�^���Y	�J�l"�9�J�.d�C�XҜ�i�l��s]�i1T�[�*�%��&�
�	^��*R������,��+�WFBbUԔ���#W6�������B�+��A<{#:�U�F�gAgmg>��?�𩉔]�;�k�2�P�12x�P����ںbb��9T�e���h�f�c���I�,���"�7�OG���ڶ����z���z�$j�j!�	'u�����(�j����X)�F�5ɣte�k|�E8�C��^n�hM`���O��P��7>{kQ�V�M���7��P;?��PPvѣ���Mm�x���V9d�:��K��6%N.�<�N�w���r�\*q|ۑ��F�j]����t�Vn�/]Ve=�-$�^^��3j��P��_���O@��`^i���[1�>t�~ͮm��wq�F���� �h~M�Q���\�3���Ng&d��\� �ˁ�Ɠ�y�d���-�%f����۵�:čZ'�����CH�R���*P���ǂ���҅N����e��`8���c�
�eګxd�!]�l�Ombg(��=��Q\�x�������΅ `7dc�/�YD��2�]���6�q�ZI��NV��}�y�s�[s
�)j�Ws���4Y���#����I��n�F��&_p��A��2X���ߞ��ÿN���M� ���j޽�t�N��}��I]���5���˴��?�@jaU�� 3Z��@4��+8��F31F.�X�>��K(?I��.-��y�'Fz��~��.xf;��D�o��.!P�3�GIL�[\U�b��$,�fa�����9q���dH2�c� �bЛf�v椇�m���ra>j�h��Q�i_v�b|��-�1<S;�e��2H�N��#.�]c���4ℽ�:J�\�� ﱦJú�aR�h{~��n�\#)�혬F��^44�q���2A�*�R �7��	��OҤ xd�^,��v��P)�i*�c��x�
�ѢM����!�MW0�+���N�HE�nE�����**y��8v�#��R?�Jq�c4���O	�N���#7R�@C��G�=>XmzrC��g	�)��� N���܂��eC,R�U_�}$���l�����2$="EP�n��(�k�g��B�I"� }��ǕI�1|!�<�-3i�>./�L�U�3��;D �����e�=��y+"��q;���Y@B�+#�0na����$��>3'�R�<`v4���;>!��<ȠI�Ȏ^�5[�K�{R����8�� Qӄvq�W�M���ÈQ�0�nl�;(���x��Nwߩ|�����mTlú_��m���n�<��b�Q{���Vsr/���5�~49�kP� �^iW��s��6m}v\��ar������K�7ϊM�,�2 ���c�V���+&{�;��3n\�,�L�&�v���{�}�~Њ�cP>�9�ss/�Fq̬��D�\�?^t��UT��Y[�v�D�t� m�p%�S���Ȉ%HBt�K*=Q�����c���i��u��S:J����l��c�#�jAD�_����xJ�3wQgG����ƕ&￺�\�X.��J�u�kxͩB��s����(lmP;7�N���۵3тrP����m(I/��t�'q�(@Ӈ��1�/|q.w�Gҹt�@:QHP���gܶ���s��q4������/�}jn��>Z�n5H�`�ut�0�w�H$Aa~�����=���9�� }���s��V�op�4����UC�`-tJXkAC|�^X�.X�|�;�c.�.��&�:���`�'��X �R�Uy�<�?b��T2��n��U#���T+����,j������!��w��
�9��j]ኻ�[1	&�S��rr
�i�����w[%R��}��q`�u�N(���ߌ�&ZK�bc�M�N5
jeزP�zD'�Q��K;��[�v�[���|#�}\�9�$�\:	�x�Tσy��E2�3��#��U�7�ڱ�]���ٻ<�Y���2x���&�W���(d+O��C����_eǁ��l��p>����|$}:�i�9�����)����I���0�`�IBׅ6�Q������3L�뭓B�n�~X�"0���� ��ͷ��lRcG����$�՛8j���W\���yqc
՚��#���U���#��WjOmt��\�|9̎y\Q'TG(��S�Ue���}����Y|���vA"�/��o���'c��kjl�l���-E����ض��`ݞI�R<p�y���>�=��b���-R&�E��]3����0�W���R�!��(����uHV��fy���5�8�̯H���h���YO\�P29N�ʌ�z�ޣ�Y,e�H�L}@J�:;u�ܾ�/�w�5}{����N��s�1$�ەǄ�4M�!|R첞��n8?��W��}Rc����o��j��֎�`v)Jo3���/��A$��������Z���� b��c�oſ9~Y��3����<p�oFP��)=�)�=���`�Ϯ����Lݰ���)�5~�UA%27����ɖ�Z��>(]{�<�����j�l��ba4T�9�쯮^AֺVv�|bTO[vU58m�'A�waW`,Y�#ͫ1�wW��%�P�Ү��[�uވY�z����Ө��#�IPR<�?eU��m��U9������Ą-��9�O[��߻R�������1G�<��D�.ۭ���\{Hpː�;�-�p���B\�(9i6�A�`����KV�X���Wgluh���Pw�S��{����zEO�����׮zN&?!��8���3B�<�=�t6�m�)e�u���:dX)FЬDD�Ve~v��k٢kVw���.�/{5�����\�}�h;0��=rPv��v敬 ���'�Fr�g��|
{?���p��9L��&�1T��Z~�	߱�;����ǃT���ֿ�� v��5�u:3���Gt���ሬ~1	��� (��8oL)&������?.����Ȏ&l�ৣg5ZJOʓ}�\�`�y��N��^�C�uX�}Tb��	�	cW�"T��!(,۟b_a���ρy���SO��AK#�M����U�V()5B�V��١�者_�4�^0���ck�F�1��:�����f͌�w�� ��s�W���2a�E5�3?5����_��!�C$�a�#99l������ĵd�X7��	W�^���5��b#�#����R���D�W޶m( ��OuثDz���/X�4Jv�ˢ�X�u �M�i�P�`��'AN$	sH���|z��C;��g\���g���v�F�>F���Q����l�Y[�=*n.yY,�㢼�懎2P_,�m!w��6�(E��M�a��h%�c�պq�F�3P8�c���fF�;��U��xg�	�#I�V�_n!���[�m62����	+����,�h�O婀�EљD�;@�?Z�H
�ހqK�X0���lS,�`x�-_�&��/�4�9�@�
���n���=ǉN��.a��X~�KJ��3�,�u���(į�Ϣ��7�4�2��Ѭ�g�?�|�uB��P� �iL��!B/��b���;ˆJ^.,�yS��h6���*β�;�~"��Rb��jjR,%��#�L�#�?��������߅�.��yr�1��I��� ����K6Z�O�9��ƀ�|d?��t��e��'�
[��4"7up��T-^E�[��&�W�����2��l>��q�oJ��Svm��H��s�9&������#'�s��u�R���C){�Q��<C��̲�[樏�휱P0��fZ�"�<t�Ѧ�sM�Xݗ|ի����y���o鼼�����s�i������i��'\oF��5��k`�C������e���W+d,�n�`�o���y�:��+N�k�LY\���l��vR�34�B���E�ա?p6�~IL�e:�F���U>k�]{��h�v����s֒Z�3�e�]�"Mx&�Q����}�G$�����`d���pX��mX���0��bd����%ؓ�_����~��a^`�< �#�#@�+R۴c�ў��/zh59�?��8���ɀD�S��m��p�Q�E��G�W4�F��Sw�e�s�E�8� u�\�su2E�a�`-��9�S�)�w���o0�y���5�0Y3;/�X��e����\��) �/�����K6K�;��i�?(�M���`��Tq�Y�ד�����f2�1�ds�سu�Q/G��
Q�A��������v�*����W"��"f
�J��FZ���"�3�j�4~��븂n��$g����v��oy�w��7H�>
�
=k���2�����G���t񷢙�4ZR�:�VR�Ĩm���i�z$(:b0s��/�����?�ߙ�?�/�4�kǭ㵗ӯ
�VU�B3��v[>��Y���/����a�{��ёY��P����c�'�L�3���&f@����X�[�]����A����s���]/�^'�~L<��)V'f(�t�G��G䳀<�]9�������ߘ<�)�=;U��r��3:��>,]�e��ճ5.#e2�Z|�l�e�0���� }���r�>�כ�΄�>�!����|��~SBJ�a��j���g��|��/g5C�6�iDt�7w��?-�h�R�}�ñ~���[��d��=�++@���� CN�:h��E��G�^��9�3|{�U��G��6B�LQ�b�i�����o��a���oe�*B���;��ބ j�z ����՝&A��Z�!v�[��`�9�%�bxE�|��](�m���5OK\/=�Z}\Ȝ��mr�F�eҷ�S6��S\�.	,*�.�ڿ�]��Ə&���A%Ű��9�kԢ��B��x�mp�����w`Bi��j���pR)�t�q5��wx�'����R��Z'�YHIA.`�w\<��_M���A�d���T�b=��k��ϐ��rwSe�v&��U+ʝKIY�g�~%��s�E���)�Y>�X����.5,�:�VϮ�xL�H�}D!����2u!�Z�ύ{i�Y���KR6�o/�s��b����'A�Z^@Tt�-�vI�SZ������۔�p���5�����RQ�B���i�
h��\ܵ��~HH݁B�C�zɘ֓lq#n��V�������^���)r�b�,��*~��{c�MO^k�s��}#�JZ�a˪�d�Q�bI~�	/��H|�i���SCp�S̓Mpw����Kl;J=�ͽpDb�ڀ��o��k|a@a�Aj�5{�9�ώ��tp[���?#�X/�A�!�^˄3u��Z��o�)y���)}��-���9)g�t���`��uQ]���V�\p� �3�V�D�8�����7��I�Z��mS�<�����ݟF�)|�ݛ�����T��R�3C��0�2���s9����� �/jt#*���p�S)ڛ�ĎזB�����.�fx��q��/�5� J�K[�=�i�!?�f�E ��]�e��ɔR��ML�nµ����-�:��]P&U�[mr����D�f��́�q
���<(���7����K3yu��7�)s�Ӹ�6��Fb��r�O�oE�sS÷�+̽{F�C�Tq>�z��lnMF48���4���UB#`�s��碱{M�z�B��N�˼���)et� ��,_j������D���FF��FuRj��ʠ0��}N��0�\�zU��׹�}���[��Xe��.k��f�����.��)l�O1�Hl�ް�J¦M=�P-����Q+\�,o��9%�h��������m�p���l�IFOzN:$���@�,�[F��6w$��Y��;c�1b=�2[H��Ln	����@��� �AX��U_P��k� ,t6�w�ڕk�mݳ��k��F91��g1?��)����uq���%�����^�G�Hþ�?޼�PB�+�W<�<��쨢��˨�uA�Y�;�W��%z44�,vb�4f�&����g[7!�3�Sѧ����jk����-����P��&�����f��zxc��=�������4�bl�囅~u	�y�����l��?*�+�s-�G���뫺�T�8QN�2cC��� �o���	^�D��x��e�a�.NǠ�mQ�|�����F2
�c��ܛ*$��H�:��bso��\[P��-h*8>��4�V	%o�_�
�R8m�dz�T/8����D��� y�sz	�V�A�
�"�|��P�A�Nރ~�#%}��hɊx�����.{��7i�`d���rE2t^��C[�ՂBs��Q�uAĒY�ýq���r�3Rۼo�;�'���-�B����}�X:�Vk� �r,
��4ȕ谦��MCK< d��l3�鄜�2!?�J6_����uC�~��y'�n4���n����ջW�ۧs��k��/��`���ܼ;_L7���� ��݌|�{ȁ[��B��pE��&����oO0�ooRְA��I!G\�>�T�[e!����j�*�4�pm���#���pJ��WM�)ҤǝQ۰�?jUT�I�M�h;��y:�
��q��@
(xb+x�n���������<�<vqj��fӼ�j��B�ܤtI�R�Ĺ!�xO���ԕ�P�� �W�Q�~cKv��ݧy���T�!���N�����&ȖC� ׎zk�g�E�s?�]U�w X�e�zIH�Z���.�����ԣ8RU�ZV"��u�7���-��`��t�,�42�������Hcr5����$�/��D�������&��)q� ���m�U�hIC�!�%HGj��Y�]gyRv��{�'9�R����۟N�u�8��J�y����ʕA�׎h����\>0E��>Z�4n�;'�N�!6د��.B*/����@zS׺��C���݇B����B�;L��HP���s�S���cb�A�'W��V��ڄ9f�ܕgZ�C��m,ds!͎���G�913�P����u5c��
w�#-hj:2��LZ��3�=��L�-�=�B�W���拕��[�����Q�_}x�؋f�e��������[;<��͊?c�˥T"T�kЈ#	=�&.L�T�g�E�?Μ������Q�_�h&�k�-��I����S�Z�`\���'��<��@�9G����}�T�>\�~��UdD�P_1�9M0�$/ׅ���fJ>���%}㡦�����U�%���:���+
�~�f�J�#�c����$8s^���G2_*�]����"m���e4LJ�'8���/�b�����r� \��H{�.��:3���U�e���Լy|2V�\��i[~��f��9�e��b:]��Y�oy_����p_� k��~u+�%�]��8��B��5s��.����,qP���kMd_e���?�{R�6f/�A.V��c7�6�/{�N��t�� ��n���M�O�5�I��C}���쁄m%Ȣ�=Ev���5��R�L3�D�t�Nx��rͦM(-ˤ�JL��E�������=n�:^oZV�V��>k�c|uBA���4m�r�;]m��I��r��p�m4���f��dQ�6��]��߳�m�w�j�7r�� rh9�BLr@��ԻZ�;��"��ֿ����IZ�9�:ΰ�4���=�z{Bg���Y[���o�mf֐�	�5*ly�C4T��	8�F�T-�̂p6$O��e:Wvu��c�X*�����?k�k9�D�i��X����F�)�J`K��O4�W�e}~��3;h6�4�8�O���X� ��n��ǩV(��p?�C`0��V�	��v��]l�;c�#t_C'Q��	�X�d6h$��b\b�;+O8�m[�8h�e��ୀ+7,TxQ,���%a�MJ]�47����xKPx[��K���Èҡy[ "7�?,_��j�E`����]>
O�
���L��iء�떸��f!�?uY�,��
����o�	Ө�Q;v�-wH�_�+���d���C�} G L�����2%ܤ�e����@7��U[BQ������!.>����o�
|�r7\��xG�:X��K�"�V+�GĬ��%��h����i�AGf��8���l)a�F?��1�xw����G��GP'��P��I�m�|j��@,��_���cCX"�y뵏.m�δs:�D�"};࿲AdP�\+�h�+��z��[Z�r�L�UMЭ��<se�˺��BXy�~�a���@A�M(� E�X�)�[�W��g����yo;<����T�n���f���nsh��h��{���=�o��c�GC��=���kL�HH��ڔ�� .#�S�c�:�9Ɲ�� ��[�А��i���õU�o�u�L�V�(,�J�\���3�K�L�\��'����ơU���tss��(��NU�-!5�:����M���ٹI|U�[D,&w��Q>�OFz�G�ۧȚ��X��Ny-�_C�\�@� U���YN ���� o���R%C�i,@]�l�
  l�hE*~Â����a0��J����w�YE�83�r�Ҙ0s�I�T�e��h_�fδ������R�]�ܐl��ƛ���'כ�����Y�Q����p��c�ҥ�>���رUt��i׈f8�)Dw鐰��0�^�}����1��9���"���_��̀�e�ԷK)��ح��ɶ��2��^���	X���K8i-��$3@}�ôN����w/�9G�-c���w_mi~	��!0�5��L`�[����-n>�;�U��ASe�
�M��B 4�e&n�NԐ#�\��q��oܛ�*��V�����{��M���A�ͭC�^V��5�a�ơ�l}��p���G��ؚOKg�F'�HI*L�#|%r�,��$�*�6(�1&�2ݖIF���k{E�ej,Ah9�V�R�
D�p%�Ǖ���mi�R�k�*�ɐ�!�čd�5����u\��>&�x	�S�Az�)�,8|��?IM�@)��Iճ����"���]<��E0�v[��e8��"@�%d��0���P��g�m���ٚځ�B�*�.�4a��<�Rp! �D�X���D=��s�9�	eq�7*`�}�[Oҙqޘ��O�R����F��Bi��ʇO�&�J�	��}����ф�v�}6v�A��J�$uuH\Xr��Rg��\^���H�f��⹱��!�,�HW�_u�n�X~�E�8A�T���� �#�42�yƱV�4j}��|u�QE�ՙ���w��� [#�N|t�u�b�Z&�w;u��t�TG�̌�?�{Z�FG7ȃ���j��y���]��ߝ�h��􎦙Z���hJT/�X�n�E�x�͞�~2�BTvG9N-��+�4�;��o=pP4|6��ǕNi�t�;=�%�B��@�90��*�{c<�#أ�s�ϩ9��75dħ��i�R ?���Av���Z^�8��`*h�@h[X�u�s�p����\C�wF�۳ܢՉ�U/�£���	$��\�-ʿ��S�!��z �Y�Ӟ�ɶ�Xa�m�s��ۺ�kn`$�p����lcx5�9�$�ѭ&��&+����W�	m
��[8؁��k����e*�Hfm�6�"�q4�;^�����'��A�PU�D�Mi1L{���S��3�hlN���axwgыQ�~W�[��j�X(��cz!.��3��S������F��\�zV�sg����B�h�F/U����r	l���ׄU��!�/�����	hmX�:��>���b����Q�B�Tሓ)L�%���2� �4���cU;W�t��4���ۢ!��C���;'��C҅j���C#O�U������dGBԅn�/���5�hC×�q8�g��6@Q�������������!.����]�,ۤ[�Ҹ���@���]qP�����Gw���;92��H1�w��"�^�H7�bA�fAl�Ϥ.��-{D%�OU"�6��y�ޣi�I��j9D�ѯOj��ќ8��|�oW"g�A:ݪ��KE�l��/:�Ů�f3��UIa+���r1q�Cn"��7m��3�^�~�(oպ ���ʁ<�� [%s���&*�aj���fO,�9���'�n�¸�	h��-����v��G,�Z��oW⥋��S����7��jO����q�\V=Y�M�����;��S0b��jŬ)FA{�K�p�4*�V�D
ؓYȦW�^l����n(.r��k^��H�c�j������#H�~w��JJ�*U$�u�EƀT��HǞο-x����v�iҶ�6�4��84����e��.~��t�F�"C�ΊՐ��K��	T�?Y����*�
^��֔��_b#������N�NNC��$:[�_El�� ��U�
k@�����)���l��|�늢Nw~I��t��]Ef]@�J&1���Hnl�
BOj����@�����[��YNl�V�)|77T��8��Up�RC�lv��~�ïo����N�!�~%|ov���W�\�'�K���[��:r
<�4�S�$�|�k�h16����i\���X��e���f&Cɫȵ>'r
��R��	<Mg׈��:̈�4�l�k�R5�/�ܦ����=�Y�J?�'9�f����f���z���x�Mo�5��
U�� N~��̤j�L��)�W��)�z��f���;_Wu�)�VD'W�����#))p'��Ν�yQ�N���}�,/	�LΪ@L�]3�T��ݎ6j��2K�)�(@* V��
|��v�@���lOLH���֭8-�^����V��hu{j�ǈ��Y�:�����\ZY�Y�����m!UV�z]V��><\2�r* F�"�ڀ&<�FM�������6
��c��`�V�|ou�B�_	�]4i�����@�r���h��.��Ӣ��ʑry2t�ee���i=��t���/��wPT��|6���%Z
B`A�9�h5"��4'k����(r]��Ts�ޘ����?C�xC�ۈ#5�4�x����}PZ��"�2R����;��8�j�m��!]��]�ߘ�'jj�P��7���Z�l�j>٭Y��>�y�%NI�4}�Naa�k =n�pS��
fN��ˍ�v��K�JV緖`qG���s���y�NQ&���G��uF�Xgh�]�}ǽ��H�<�����uS mi�]�yK�!_)���f�o��+;o ��{8��DＢU�T��N�*<�qڜ��g #s!X�9�����tk��
�p9\�7��C�L�}A� �=�n�@-ZB�.6k/�h�Z�U鴜cc,����]��l\4OeS�N�5���
�
�/[qn�Nbp7�J�kd5-���	��l0�T�q�`.?pV���Lg\��W�^��7?���h�H��1%�UX���ppG����[�#�6�_�z�N�o�������q-�+��]�X�Q�<K�'t���K1�G�x�����-�{�.���Ք�b�g�fܕE'�����˱8�^����)D�H{+��8���M��� &����V����g�zݛ��Ֆs��L�$���>�(��3V�q�mg5�m��2#���5>��>qb�p��[t:_vQ�1�x>|#o	7� .���:�.!
j������
WhI�H����A�:�lsc�6�.pHoF%��xU�`�j+�{�.B�y˿_1�%�� �/%JlA�����o��f�Rx������^�$���{��l��Vu���)5n4l}�+��b.�m�ox�0���%���%�0�����+���z� �[�]����"	 ��>�v��� U*�w��i�U��-)!�h����(&����y�\���4�?��&�O���MmN���@N���G��~�U�Z�T�>珐b;_�)Ɣ����� ��l4�������p#��R�<J%�.�dEa(��UC��̲K�]�R�"� �=�M;�s��O)��:ȡ/ ��f��X/�$]y�|��S�qc��)\dE|͵=����c��Hk*Z3&������1�
�ڏv;�~�,�v!¶_�Mf�E��,��ć�pq�z�0�I�]ώ��a��yP!�͵^;,������yh.ar��F'~ǰpr���@}1mk�\�]M��V��Ӵ�b�����RxTuY�����l BC����rM6���8�;�(�,�Ś6.+=V\b��l���G¥���t�&�.������F.�Pv̩]��C�6� �����Ȉ!@�B;� v��ǫQ8�N��5#"r�o:G���QW��.}�fs��q�ʫ��I���N�U5���hH�YYu����S%u<��Geb�?85�P���*���B�^���u�N=VG߫1
oV�̣O��6v?6.z���8sAuib$p/,[���sd,��_6��K�����c������g\N_��)�𞲟��Q�5���Zs���Dtmb@��w|&i�'Kmb�M"
���Yв';��>� �V���Q�TayL��w������gJCB�w>
�f�U��~[ą9��'���&�B��X�����+����������G�d��d�e	5��܁*0��X|n���B����c|�L߫ge�[Fi�"�z߬��#g�-�j�����8N�A���/������c�snm��� IAUԳ���9��|	�N?�쁀A3��z�)�!����Y��R��Az.l,�.f�Q ��k�"k��@����9��"ȄX�_1B��8�zYhM�0|�W�cb�I_s��׌á�^�/�ڻ��e*�o�m��z�~��ؿ�����=�(`��^�N��KF�)�1v�l���d����H�}�"�=�B��
��%f��@:��{�{oj	\}ufhjh(Ɵ(�G��Uld�&?C���+�����D��!
��6 IR�S�j���㻓�y�����*+T9�f�KY�a�}u���K�΍ם;������V�+��=����q�+f�i��s�0���=����R�������kNU���+i@�8J��ib�[#)��G��Ub�}n���T���"�c#܇��6;y�`^w�@0�E<f��cW��,��'�m����S�p#6��$�����sn������#~o&���g�E�5Ӧ2�Q�Z'o���}�<�Us����+�/ѝ\��9T6Q�i�g���u�*�cd�k~6�Au�4���u3g���@,�߭"=W0��=�wn�T��R��M
�DX�:�d�<��)7� t#�O�5��$3�a�a�L�*���zc�<���� ��:�떓,�����x�N���]��і}��*�X��G�y��iӈV;51o�'jj����x�h����UN��E,�@�;��0�ܞϑF���WB堹'���*'��S|h3����
��*��X;$�r��΀0��j�O���D��,9%~_>lI����&Νgl�mY1Q�/3]���QY�������x��zAu�qq� ��F�f��c/I���V{纅Ȗ�REǒnb�G���`�	��w�@�fK�MT�"�i�˔�2���4�g���t�d$����QU���@�r�>3�>�+�/��6��S�slUxs0�^Y�H���޿��9�����̶��9	�����ƙ�}����_Q~qv�}�I��+)��	�:l���6(��:Ź�{���X���s@уMAݓA���ŝ�)��y��:�}��)�+t��.��ñe��|��bDeK|ߺ6M����1 uI�A�~/6Sz�9���S^��H��P�I7��T�������x�z�G�v�v��^��s�i�]"�Y�B��w>��#�uXӤsK�q�&6Uo�l#�� �Ôv�5�
{�G𜨜i�L9?bxP�f�:���F*ӟ3�+��p�VX��0#r#OeM* � l��2O[�(���LQ���Ս\��D)��Z��q�`�\��ce7��t���e��92y�v��{���۸��l�sNz��\q��=����3	x" oͬlX��7^��z�����K��V�.�0�NԲ��̈m�i��uJ��i�an�s ��l���͓�Vf��l�8��$T}���pJR�J�F��0j��+N�ɹ��n��Q���q�c<d�H`��$Kh� ��?8�0�文ENHL�c��v2�3�}a/��L����v����F���MK�&����d`��1��<S>>�E6hkm�'sw�`��*�̿*:말ۥ�/�x�t�.�-��&�����T���f�Neq��o�:L�Rc�� �-�
�,�S �k���e*��`~�h T�r.�='�I�D���ԔL��k_���1�qr���3o���� {ۅ�朗s�SIZ��(� "�k#za��舐����QN>���}�zM �&�0�=<����'�<�tn"ŵX���B��y�9to�O1ݳ��K.�o�)��M�ƞ@k��8��ı��>��W�]	Y	�DNї�\�Z�^�L�d{�a-��D�0t�&���*z�Sb�:�'+ª}��5�
� ����Jܝ��>�x�-.�2ߔb�c2���D]�%
�)�%rP�Xf%Wk��1]1�>B���!�O!���Iq��=6����b�|��+���ܟ���r)�	��*���
���M�ȁ(�0r�� [�W��<d�L���+�m�c�8�]�V�wW�,���i*J�b4��X�0f{3��ĸ2oE~�-�]���6~�u����V|U���<��[�vy<5���6T'����0���Ϭ�kߩ�'��6ƒN2�"��_��@�3>vI���jC��G&+���{C���a�wUme����A�kt0�<89�<��4i
�U�֜�K<Nv���}6�����h�p%C��`"*C}�k�q{w�[ʹ*R���H&��=o�����ˡ��i��j��'8a:�߃ �W����.��똥8S�|=�&8K�%��,���D?��Y~}��H�&#N�aښ��'���{�tMP�8YI���6@|r;�7y*��|o"*̡�A��(:��;Kϲ�$�s#�Ǒf#$M��ypH���x��Æ��a+n���6�5�,Y����%1UΡ���<SØ�r�J�-�aWJ�hƸ�ݫ|�6�!]c��G|���=��c�v�"�����m�I��q��ܣ.�C��?f����[�3З̥`�ú�`#8S%`�#��!�2�Ot�e{ݼ��tg������R�JU���H;72d=}�{i���u��沤#������X5"�ߟ@z����ܤ7��s����k>0j
n=�c s��� Ă�}�[����F#\lj�ѣo�;S����B�( �WN,�Ԛ�q[��l�A�C��~��(/��Mr���g���Q����;�8Y��1�&?�F����#ډ��r6Y��'R�2<�s��g�2RЗ�h�~�J+Ap��1#
�4c�Ϫ޲�O��sG:ˤ��xBp)L�P�ݔ�Z�_��|���>#�1!�S�A�z�����!�jY$z��~}:��H����mb*� ���X�
[K��~�#���֜��|@ML365���[�*_���[Ø/�:�p�ks��Q~����	�����%��_bkSj=�7��$������<s����l��U[��?�-@i�d;��-+P3�Je���k��Xǥ�j-�\�S=e0���֌-��
��M]v5P�!��P%S�R�ҋe#<Gc��u]��EȄ��R�O*��X��l֔��])�B���#yL���Hۚ���vu�ļ��i�'�$%��`�=S�űP ��Kq������y���B�' �"��B�f2y��'S�{O���9p�F�ms�G;XV���=( aV�tS�0-�K	Ve�؎�[�'�{/
h�h��k���G�G�������}w!�XHl�bTft��S��Ŵ�ކ���޽ޢ�sLY�-O���
�̢�G�$��?,~^ ��<j4��������L���㓇��U	��Z5���Dɸ^{nB~Uz3�:Y��e��xA�� �)����fwuF��&�t�r�������a'ɡ�#f�;����r��an����PdnW��u�����$*�{�$kKAv!��;��[mQ��� �w��X�*/|�>�Բ�/�b�g:m�M �F�2ê�Z��?/ig�'�c�
�6�����N$�{���)ύ�[Q#Ck��i�崏fG��%�����G�N
xe3w�rъ��w�J�;�5�?8?�����}:�������O��o�G�-B�}���"�4�}FE��6� �IV\���V����s)�2C����x�!̊~L����T!C+�'sk� ��:)|Uf������� �����g:q Yq��L��,��˔��;���ސ�$jJ�3�0%�M�w|;��u������g��j	��1K���WiTp�l�x���X5An�^◒�g�\r�?�)�*�[���8��W�_ļ�K%��kL�F�#KF�;�΂�,��Y�N�e�HV�I�5�`P�������?x�������x
K�ߪ���k�m҂�������OL�k���B�G��ا��#�A(R�#)�>����Z���PFA�b{�Ő�K�@��)_X_!.3L:�2#ݼ�D��z��A�o���p7�a�%�-EC�%�bh��VS��7g&ʣ�\G�-!�h�b[�kcQ�L���[�˥�Ѫq��%a�i8�%�n��_ye���C���h�!�n�k�%A����$��zGq�!_Z�����rh�W�U�w���'�b�D������b�ҵU�@��6���何}2���ݩ��W����LQ|��۪RZ݈Q���r�����Q���$xg<"�Ov�Ox�u3W�h{��C񥂅53���\|.Q���z��mD<��K��T�ι32|��JY14.Q��y>�a6T)�L;o�ϱ��OB��S�{�� Z[<��9�X��&�S����[&��/*$yJpz.������G��,!��C�|��]}���Vwn.2b��A�'BhLO�����x7�����r��$�%<Q�$�N٧^�]�oGDK��m�:�1�0�?L+ڳ��,G������ڎ�ׄA����E2@q���6���<U�Q`�Ռ�SJhJ�,>o�Æ����e��GXA��x%�󼥁�~q�+���3��bC�KJ�@B&��y���g⚻�Q�֧I1��2ԗ�@����Sp���j*��Y���w �c�&�QpC&Rhow����u��Ð�|ֱ/�_ѳg�n�[�}���Y�t|�1悦�x?�2�^~upZ�4�����)�UsN�07��@t��~����C�V��]�s�+�ѹg�P�1f��s)\|���}E��mTh�"^Bs!�����m��H���A�;ĭ>V�D��5l N/�b���vZNC�)�Rzx�E"��m��əm\6�g��u)��[��qu~0ln�5�hS\��!���U�Vw"�-/�H�����ŧ �YR?ۃ�ل��a�s&B�I�QI��lIa9h��� ���1�'kaws����S1%MLt߄��c��.����gj�Zu:����m��ND�Bg��ǁ����G��F��'�%�d��DM����蔗̀�<躾X�`苣�R֍?�<j�����J�r}�dK�7�ǁ��^��J3S"��P8���=|�e,Sp��;�G��D I�� �w�	���Eh���.YM��1=�L����qy����n!Оc:�#.;]��1r ��H8Z�� �;W��p.e�y��OrJa���٭�=�A�i{E`Q�÷'��'a���X�h�2?��^��0���mJ��4駍p�(��KDE$&[{M����J����$�`�����eb��$%VS�gf��}�JMΣ��1����]������|���v���o	WZ��,�M��B�-v?o��\kV���#��$Z�׺�P4��\�Dh�5���j�Ω�ǟ;��M �Jc�ᳫI
���`�x!�ѵҿ١4�r��fO��-�-
�\E�6�Ϗn�<���l��5]!k����m��H�WV���[�qվ��XT�� �Q�7C�`���f��U�ӎ�= �vޏHڕ'k@�G�E���L��S�Ѹh'��ѯ<:�����v�F3-���XxHވֽz��+���g�4!�3�)��7u�hd	�1�Wj����4is�F811C��3)t��:/�H�8�m�ʝ�������{����ac=�?��G�}5i���3 $�E�����[bϽ��W�[E߾�v��x	�	����7�T��
d{������{vMP�r�R��x/2��$�����~t��}��2	KQ����ޏ�OjD\�C�������xWL���ݵ��u�`d�W8N��\gڒ R���@��# ��Э����K�آ�ۡ�$p�'/��!T�>v��R�Ġ	^�۠�<����a�>�p�����6x���x���n���8iH��cj����i�``4�Z�'�������͂$K�A�
𥭗8�����~u��|g*B�5V�۪�D��F��G�������{l�mY�K5�
ˁ{X)�sN�,8��}֟2�u1[F�ԩ��D*&T�>����(��/%޿X�slIɵ�.>r�eK��E`�)54�Oտ(��ߵg�+�p G����Uu�J;E���\�����9�t�3�`�vmt�g��p�]`/%!�l�6����#ʜ��}�_u?*��p���*�"���� �s��EK�I�Ү����K�7�'F���bP��鄚4S�7WF2i�ў���d�������˳�/�^��)���}���,��mi��;yA0��o��E�l��4;�k`���{$/���"������ezLB?�q&��q$[LA�@C��q��~*�7,�Ɍ�{��;x�Y�:�t���!����v�]�NfA�AU´��b�Lu۔�a���/�3I�at�����'9��-d�2�'�pn��.�Н#u �i-c-���݆n��V	�����©�C���z��IR�G(r����>���E��e�mថ+j�p�=��X*�l��x4I Pۃ�>�N<��K��a&>XX<+����l�Ep�N�H���ّ웯.6+��~�)��	<������:^G����j}�&_��dK�������++��	o+d�Ʃ���Ǩ��N�z�!y|(�T�O�8E�-A�^̄uw�K$Mŗ*�
�T�m����o"��TGɚo߶�F�Cr��͜�o�֎�(���[ٚ�A$��X�p+�����oɊ�f��D�����گ'|A����ueh��%����˯��o;��ݥT��e�L%;$|}m�!��p5C�s����}�n�ډ�ij��>t 4R�׉�����B�hziIƵZT�����@�Z��<��cr-_��ܟ<��p�k�@�����q���(h��3��=��&���𶫾��`�!A�J(j6%��ZT��f�ϐ��F�*i��.��-�RdC0t�e�	�D�����ǳ{6{�]3r�����jX���8vd�><V"�aK�&lo�I��ʃ�c�!=`6�mq���q�}�@E��aPW�<�[+�����{m�$�B�3D�C5%��J���Js�E�)O�dr�Buy5�b[$(<���'�P'��#����q�KX\�mT�BƵ��߰-�����\=T�~�N��yJ_�/�+u����������0\G4N���x�
0L:���y˔��7W�j�>�˱h�����d;��� My�=������q��Ap�(��hL;>>�]7E����5�(���D�����и3��%�Z�2s���9ob{�����q��Ɵ�o(��S k�f\�C�e��"���MYFWN5!�y�5B
`轆J#R+:��/k��ف;ysv�A��1�4
���G��n�#��pr������4z��Pۂ�i^pe�L�����h�>{��|�+uq|Ir���W5v*e��T�J+���H���-��Y �r�k���Q��d�O��+�>���#��h��.�Ǌ�C�WJ{_�I���K���Ю �2��^�S�XFm���3L�E�-wQ}93m��K6N�p�T_����o��ƹ)��|��4�?M��-���9v�hܔQQd'{�Kir�B��N&]m�� (�\M0>E��] =^�K���0ȫ�,��8���Mr6�Z���p�~+��m��k*A_�>JT�<���)�f���uk���}�ӧ9���@ۖ��<�����$�?��:5êL�i�"- �<�W8��a3LX��.�΁�:����b�q��hG������N���ɟb��"�pnR�,kҀ�z�`)���.��M�IS}�-��u���܇-��] �(�bچg�sGȘ �+'��X͋"��-��/c�{��|p@k�.Z���Xk-E��Y�O����8��Q.���)@M�ץ��L��6l�Q5V[x���Cr���G������dJ�6�jߗ��0��h���q΢-Z&	�E?�AUD��Wo��T�����?�"�ރ�j�{颊�)���Ї�V~��7ފ�D�VI�Db(P`�3Ft�u�������룛�~-yX˗�P����y�����]OUL���w��&����������aB �y�7V�d�����:2���f�\��%��=�K50���y`hD�/��E�i�#
����w���'M*�(�x���૛J�1��V��p0���ve߉i |�H���It&�^ź^� ���]`�z�\^�O۲v�S	�3�,N�>6_"�=�R(0�yiJT�R�������s��N����9��܏�d�<��*����	����'
��u�%%�>�{�9�1�ar�Pf9&7�-v�y��ŚH�����=i�4����O�C�1����b�x蓱[^�k1�:�q��:ƕ���V �k^��	�Zz��\�D����Uy�M\--��cy2�9���!�����%�ѕgq�t�us�Lzި2 m_T/j���)9� �{�I(�I�ު�u��'�kz3�vc��Ab V����:���b�A�e���d�D����8��5T�˔]�g��؛��!YT\���:{��2Ϩti�;.V��%�<D�! #���Lb�ߞ3bēA�xG�G��[9�����P�@����치!�"�F��H#W$��lYE����	��F+��KҎ���"�L.��.�~��!��W�Jϴ�#Bt�H������E[�d;�IaЀ��o�t}�i2Tᲆ7�Z��¸F�#Ѻ7qcs��j*9���F+�$��[�f�Y:m�
ہ�;y�6n��@�{ ������G�@-�H�iZ� �`8�PVֲY�^�T­�p�a��
��9��EY��1��2��!E�Vs>H�K�r��	k~M=�j"	��\�0�ԇs"m�����$��v�G����`ȚP�*���EN�;�E����5���&�&d��`����)!6�*?
;S�z^;B���$q��QU�8�ɸ����_Q\����ko/+uS��1?(K�2߿ӡ�U	2���P�7A��ϓju-j�Tԃ�=�i�Btu	3�knF�5����`}�oPܬ
�8�j.UWa����X��`�b��`�kOO'�'�hGN�SY3� N��$��`���SY��"���C�U���-�x0�y�����p�T���r�·g�0�(p���&E�x�m��</&���R�ʄiaA3�Qo �_x>�1�����ƙD�2��ț��!v�w�U����+w��%Y&�vlW�If�X$�s���<Y���7�i"�`0�}RP�QL�Ⱥ������ ��~\�E'Ԑ������}�e�b B�z{�[��� �{�.��q��q�$��Ş*�v�G�3��T͟���� Z���}�}q��R{&{�����֧>)�+(	��g$;Wx0V핦�!�t�'�Qˏŷ~�`;݂��3Cf��̞=5�����������F���`<�b���J��w�2�2e^��$�͕QL�bo�U���Eɱ1׼�Ou
��ׄ�6s��i������V��W����R��uqS���h�5��g��<�g�Oh$ak�R�� �Om�[6� &�
�SG@�1�`�+���%��z��N*
���ϒ�&p��V?;[[�	��C����5�ޞ���UƲCɈ�v��PH&�*�Gp9���T$Fa�wjYq/a��8�*S�v>���שwD���t��W���[��������l�s_7Q�@7c�8�|�îi��*�����M��>ސ���g{����HOW�Xk�`�*_%ʏ Ov:�Yx6�N�p=P�{\3/���� �^�Q=w���v6���4�Hm�F.l� �##��Q��ט�Pw�:
�P`�1�V�)�"Αǈ>�*�s��%���xI�
��� x�����\d�TQG��<1�V�|@� ����/�b:����X�pʄC2��p[�Y�\I�}�^�s�����2��j�͙�l(@58��f����J�n�ox�7?����s�d+�ý��>�֓m赼|���`My��p7�,xH�!������GK���+� 2��e��������b�e�!M2���("r��D"~����Y��vXQ�0�,��G��q�˲����b��:��q��O��.�Y�ej<k��z-�Ŕ)�	i��}�Bhٯd6�(��3+�dJ#� �Mr�����h߰�Fy�fn�K!ۊ���[��5�{vhްFp(�~�3�K�Y���~-��~�=i�"H�C�o�1Yp��/�v�w��2��#aR�����Y�0	9�d��/(t�G�i�Ρp�J�Lk���_-K��x�bw�ۛ�V�nD?���� xu8u0���>��a�%�`�ĞvJ��61hI��L2�$e�����`�-A���OT�;�F��/��Wg�՘������$)vDV޻��?C>a?-DVi�Z�X��h�	b}ځdo� ��������Om�i�
e�2-o@Գ�Pi��f.���Y�ȅ��,��y^U�|����70ޘ���	�{D�X(A��D�x�x[� T��"��[���H��O�I�X8H�5������C����l���V,�����=�e��ln�=� N�
�	?1�����z=*������z�F��̉[��q��!�J��ôE:�$��T9��N�W�y�p6��Q�`]������i�n����p��lGYs�:�T��t␴}S��v�N�2^��a�Ud���Uކ{P��z&hx;�>��S!�6��N����#�m�&ؚ�r�-)W��?��f�z���iH�Vu��s�+ه�UP�����2�S;��P~�\�<�C� �D��.���K]voB�r�#u�>�?��I᪵����F�v�@��T	�?fV�^rf�ɋA-�?;�EnY]tu��zĨ�j���3
q�R$��{�`��0���)�'	8F�j-�坤�J8e�D�l��ia����&���d�[*�}��H�ɜ֯pEf���\�ߥ}��L��k��p�2�:+pY}rX!�~�(��o��XuPS)�q�LÑ�v$��0���:�!����R� p�s�ǫ�Agp�Le�o��l�ZrDc�� ��}y�3E��?�N�d�f�us��]���9+�X	��Q��T�*ಷxg�}( 7v��������i����H[�N��I ������@��&�9n8JlRU�Ȃ��im
B��I���4�.�}�8��h�LN!q���>���Y���:\e�}�_����[��0��}'�<[��h��+�?J�qD�7c�ٮ����_������O6��MG���`�6�]TE��F��*�臫)-hh��vcV�Q{�r�k�ԋE����kfm�g��H�|���m=�V�=����<�f�S=$4p#W0X�8�ʸ?�����;�@q.3��7)(���xF��ɫ'9���u�b��uY]���^ᜑ�d��1���@�@��y=���t]PV�ǒSeL�7'vr W�K�]ʍf�\*.(��F.�M�qE�o6����_@b�耍��_<
kD~��`�pW�����
�j��2�+��sNڂ�5l*��_�R3Ͱx-�t�{zv�`���'�^�r���V��k��(1i�w(�C�gP�K!53�Y\�a�lf�B��9�~Y,	5�x�+ܹ�<\�K��SП�QYt�j������I�N�y���
k���@:P�B!nh��M!��Dg�-�Y�ێ���	"�Ozn|c���M�El�t}�Q,p����M1U����2����E��~��ʭ?v�����(bH%X�7q����E�����p$��7���6r�f���{Φ� 4�g��2�}0�g1"v>���&�zͫ0!�E��KF����9ł;޸y�)�T�T��m��{�;�|j;���gK���`�+j%=�^#�7��%��nU��y�� ܣ�����V⦊7�B��5��,*E3S��k փ)N�nXTs����iT^?8�N�l�r":�����+�i:�C�o2������t�đ�a�Lk�8��t;�uR�Y!�.���k	=/�X���rd����&� ��q�zk�K^{_�1���v�s�I�
3i(�"e=��b����p��V��\��\X��0����!� ��������<�	�9�̧�ߎ|~ܝ�C7K�	������ `�(f�Gw�dL��A}!�c�(�mԻ6��8�G����L�oP�Ax����k�������D���j�	�X�H�n��y�`:&�c8T;/�Vo���3v�5?I>N�Y_���`�Aғ6o������_&`*a�g�<d�Tq�����gڒ^_1�jt�+�����q7Ҭ����'��s@���:� �����#[���>�> ��o�����%<��BOߖ��:+�sÇ)ct��#w.B�9Q�I>�|2�1��f�~\������OB���؜�ڴ�G�E���Wnޤ��7=Ce�~@l,�N�D	m3�T՘�XK��9��D�I�����0���~q;z+�M��NY��Z$�8����3�iec��n���.:�L(��ʖ��\�����2��l���)�M���`WkQb�.cG+����Kx�VhwS��&�ӵ�ZxP;���j]��8̕|>�9�#����dF�F�2r�w�����4~�b�Dr���C�d�OU{��½S7�Z���_��%ZU���$X�F���F�y�t���Q��<>}x�=���<z��*-OT� "�q��$��Ȇ�0ΛN�� �v���e&�k?��v��|�� ��k9��<!D�?��l����}�jwrhB�i�D�Ǌ+Ech�y���x�Fq2���Χ<��LYr���+�flX���J���T�tJ��a�,�A��Jәe6�	 �y�8cv��R�����A���ޭ~#����x��$ے���H�n39�
"	4�{��D5�����S��i���s���G��l�6G���i�At�}�D�/S*�K�&�&��4�� @��(N��oSJ�=��ޣ]����f�I]IV&w��q�.p��p@=�zI��� �'�Z�d��^�RG�8w9��jF�Z��}���.���ӵBg��G�F>< x`���L� �$EQ�'@&�V� �@C4��njAV�8x��-������ӡ�3�v�ٸ���Mz��d)��Y�M�4����d/.E��4�7g/S1D32�Y����A�t��;>A�\~��_��#|�3��q��
Sօ������j=��~>��ȂV(i���o��E�W�w�+�6��O�/^���Ǘ_X�L�@+֌����)��7���i6�ԣcsɷ�<?�p���Pӧ$��P��	���[T�G�UQC���4�e1g2d�!��t����|Ī��q���O�g2!f�*���K��߻����:xK��*y�<��1V �~�V��J�ɷ��hs��|�M�Ē�H��*�l��܆D���WF�}
4����w��Q�to1�,��&2k;V�m�I~=\�>'薱lSsA��P]��`�'O:?�r����y'_�L++&x�RM�r��~�mr�{���>yùua�5k�s�A߲�h��:yk5����U*bnq�0cQ%`W���6d��([��a�m]M�Bw����k}"�D�I#�s�a�h[�u��p�X����KQ��72:�t�y}uE�G���E\I��
�}�5MV�� C�O����D�+e��@����\�ʏhײa��1�f�\��sp�2;>f~��0�|�qX�3���	��@��]=�}��1�T=����� 0�CEp�F<�&�䠬��^w$o���E�)t.ܣ�!��A��r4{b͝>��o<,�TlXE��X�ҋ�#���ڐ(/|�EI	������e���w>
��it��E��H�$���ؤ�y�Pr@��W�6v�-�{��	��hǋ'�W|�^,S7�����B.�X��gB�Y6S�������2@���|�\��a"�mRYh*A��6�8$j�
�N?y���:��YSG�����"�V��@�����&����$@ ��)��߿�F�>w4.Y���m{)|�6��"����<�H"4ݢVǺ�·�B=�C��<�@Ђ�C�F>���� ���ct^#��	��{�M_�$��r,��>�b�N�BYc�^mZ���)7 �t%�׷;$����^|����_�W����$�����@Y���Z�f`���/TK����L����m?E���io��0!�O%�� 1�j2��!��ޕ~�y�y�=2bw��a�թM�Xk)�܂c�yǯ������o� 6Q��zn7��\+Ȯ�i���{^�	憻�������r� �]��K���=ӟo-;1�M۽|N��"O�X:@j��^Eh�mZ���l��uBX��9�R��ST��%��5>5�rlG�2��$�Z� �U�PS�	c���x��V��˚�ota�t�zu������E��s*'?1�k�̈́�3�IA�|�>�fj��q�q����,+��	"���5A�-�sZ�&��������V�����Zc����Y���U�6�>T��!B�u̮�����)$�Ȅ�8J�.�=�t��o6����cc�h�����Å�&��lֳ��H	�Wd�E*o�pP��A��$�
*j(8k�lpx4�*Lh.��R.?��
�m��7ȹ�2�?r��;~Oaz�iD�\D�:�����QKmi���.�(�V̢w��`"c�YT�Q���a�K��=�'�;TIv�8�3LU.-�7|M[di���X�Z�h �z�e��W�<�IJ��^�"�VĄ�6}5�wɘk]�Ʌ Q.PUq�M��%WڌP=8�<�V{�y�rF�gъv���6d����!��J����!b&X�yb�t,t`�������McYٵV�Q�T���~��#�L`6��#'��o��(1Q]��m�\��)ֻ)���-({�)�0" W�8��\����
�U##�s8t��5��-��x�K��1?F�lN�"l[��Y҉��Sx9��I�؊�dJPC�[N�8bpN�t��!��yN�Z���#�X�ԁ29q�4���1�"�w��������"'d�ʖ�*�n��%�% ʹ̦�S}R)��W���f?ט�P��v�&�t-�1���=u8�&ΓA���䲖Ff����W����tsы���$�ŝ��!8�Hw1��!�nq�m'�)����^�C��Cp,��lqP�t{1>x��߀�@��Lc����g����]�<g��Jmu�<�)�:N���'N�)��x��'�3���
Am#���B���O�����"R�a!'��*�Q�g���5��l=�}9ǌ?��g�{?�M�^6e~FKB2�k�\���%���H�����;v�v���JT��E��$Щ��o���>��_�Y�|�2��nndIm���֏7ۤ�Ѽ�(�R� ��I
`�������ʷ(\�0�m�m�]e  C!H�ҟ�ѵ,���+�uP
R���i#K�8Y��^����T����aw��D_���;�������7��|q�~�ss1z�_�X,PM�Br��I��	�$B"
O[��/RA��5濤!�Pi�]������w��2��M�>̮�f"���c���p-�ߑ�aw�k}~���A�kۀ�\�:)54�Ӵ��:~��S��ӓd�2����b���e^�B��n�&�r�ό��W��$�sx���uz����sbpܔ��L�
E1�����hނ����u0>�;����-��e��5�.<���&�U�t=�<��LkY!<Ia���!�d�����ۘAV�R\�	
S�-��t%�b��ͳ��0����
5���M	O��޺���nsX��?�R��<�H
�Ŧ��'�e�R9�O��U���,f+�n��}{����~�@����!聴������a� ��h]Yj��;P���xʠ,SPh��b�D�t�:e��8�x^�b'�y!�&��q�U	��R�M���x���W��LJ�{���4�rD���g����b3H�;mX��ȡ@6�"q�Sy�z̛���/L��oTbb��<�H�䫛y�WW��A�r"P�5�f_3��DL���-����b��Y>Ze3�����#��P�t��l>fz-lB���OK1�EK��A���GV�>�!���!h���᥿��m>Xp%K���kz��//�>E�֋#������!�e7]i�u�8�1:�x�)�V�XjȲs��!�_�ܘ�_���r�56TO����=�
����j�U�1Y�'Po�3f��|��N�K��������Iȓ��Y!���(ÄN
�%�ĕ(W��c�'�*��
'?x�Kw#�c�A6ur 2#/&v��(,���ɠ���ƩIJc*��3���s����r���0J��c�Aa�}Y>!#�`oSc>��S��~|W_JM1�Md���V��˳NE����!DƵ3�a'ۓ [����2=>�A^iQ��� \#0�|�D�t�
`i8x�?̬�\�&+~���y`�+�ܑ��F4}c���S&�5�z�Y�A!cE�w���߶�7j��Ti*ض?��W�G۵* ����Zq�*$?���y0'{+��1�3�� ���t�3���q��!Rc����A��-:���͠p;�D6|Vt�Uz���:7�й)sۮ9��0s�:�=����c�CNzp���v�'W�W�f��o/ϸ��"1/b8�R����:��%�iYq>Cz�!(,u~�H�ڔO�m�t��ײƜ��c��o��2�yk�vo�΅+7Jw ޷fO�S=����F�Ж�z
���Ì|(�#�K�q���Sb߼�4��c����7��)���L`�.��{|�:�0?>��X�g8I	*�K4�U�����8��z��x��(�*j�
�ސ�Խ T�	���`W�'�u����.�f�A���0��� ��.W�+ہ�vF�8��$�勞K�=0�}�0,�o���VM���o��p󂤞3�/{�ք�:�����6�V���~ �����.T0��]��<�G�{�JY��\	�̊�X���9�i'�~����'�j��7��<8d�z5�ÈI��a�+jTg�Qt�9�Qj�)���蚔�a3��N�ҡ!)�wޮP��0��o�̾=���	Cl�kIi����. 5�N�{R��K�:�R�͔ާ������5�h�։��d ��� ��3H����x���CH��3��Ty�K*`&"�2�� �nU��F���+��h3���Ę줻[u�pf��)~˩3rK��$�k&e�tw��q���y�
��A(j{���*b�Ƀ�փ#c@W����i�f�$�����/�Y~����$�^)�r��a}�J�H)Cn�B�o8�J!��.����f��A�<���H���~����
z��`�H�>��&���n3�8�7im��|�p������6��	�B�y�s�~�ߡvt�<������r:�R���ﰵ7�������oC��#0u��
8�<wD�$;���$_�Q��_?\ ��$��<�ٿ�y�U7��m�É��m]S���cg�Y�X�g���a��_��إ=�T�����)���y�V��0�d?YO�S�����J��s���,�����2�	��M�r�Z�[�4v��71���J9�i��x�k�����3tā$�\��{�\�S
:x���_h4
�x��Dܢ�{��CG��v�����Ւ�zd�b�/SՍۮ��ߌ��:��s�cņ~�y��g��ڮ^R�W���;?��J�y"��Y1����Z�����6����WY��!��Hg�X,�d��ӊ�n!e��ho~�c�����_�e^��?I��!�I����+p
������Ғ�Mɑ3w��6����m��t�������&��a5�JN���
��LF9;�E�b��@R�Ϧ9c�g�ll�{�;!/�U�N-�^Q��,���YS�
��t[����U���~�����M9�ߊM[d���Ʈ��-��D��Hz1	�|��zt,�4[���';6�g��p��\,Vr;[Saʑ�=���W�{�"O�r;�O
3����F���J����L|�-�/�%ObU�n�WC�g,�+Rwb��PzٴK�tXә��1�/�zi��/���bn��6�LG_-�g��~��U���pWw�0q�L`l>Cxw7�m�F�bLN�j	�g����Yy�s��ܽk<3��_9:�U�
�G����bi��0�Kp�I%�>��K�Ɔ�{�[�����N�g5�I�䲮�9��>H֘�u��<.�;�[W�{p��y��"��%$��$Bw�䤬��4�1�{�쯰�헮I���5��<(�����U�~�[Z�����$l��r��"1`_����[�>o����e8���h��2� ��)��s��c�_���{�>`����QT�*���)��}�^J�
Ӵ��/I��� ��9�9��W	�zԃG7FLy�n��%R�:���m8�V�w��1SR�Η4�~�
���-���
�=ȳ�j�f�M+f`r��z��gu��3���}�d�>��ޝ���Lq�����,M���1����j1Ƹ����cg[��]�{R�(R���0  �<�Y����=�� �Z��2ljA��l*���'Ј�$!��hA�T^���f���؋1Z�c�JE<0
˸�'5�a5�)��3H��nfƎ�1ɐ��s�����
���WᶳJb>_5$uO�2���&��:��y��,�3�4�"�[�޹1`ɛm+}��3kULʯ瀚�އykD`�΂��q~�s�4�N�ņV�Z.��o���x�NK�`/qQ͗��IΘ��U��fo[Jtq'��qx&���P@R��)�,ؗ݇@g�lMo::D�����EX>T����cێ뒪�S���w(� ��#���kJ���!Pu�}H�
�|+����P%Rm�D���R��ܒ>�Og����S2��w�C�]�u���;?+/��7ploAX�l��A����\��O���w]�jAjA��P�ƕA|*8y�X,��	y~��^F�!1�K
�/�`������P{����nP1BU�"�I�9^�z�����u�]�� ���)��i�~��V������IA����S��(��K��^^1=8T�i���������5�޳� 6Z��U-R=T��N,B=�`C�9��F���Ga���i�i��DS�������~RU��R�;}A8��:�^T�yV�P~�C����P��V2̧��3H�p�Ђ���|�sk�|`����~F�h��~�б��@�8cFǑ�ꮊ�A�Tz����7Ti���ɹ,Z8/pB%����&@��s�
�L��
���zd:�C9�h��R ��	�J�y��������O����ג��P��%�]6.N���Y��v��3�e$�_��#��0.����JB�ڒ��U���w�Q�ՏR6�4=w�z0.ދX��H��u���mC�r.%��Hd���H�n��8v�>"U5��(y��$����A|�5�=�F�u<!�SY|q�F��*������O#^�)OŎ\u��C�v��?��%��o&5�L��5[j%�RE6�D��u�;�׆��c&b��'z
_�oAo ����/RR�A�@~I��RU'D,CK:ף�5�o��J��`X�FC�R:��Tf�A8���#��#�kr�^:��:{y����D-�e^&x��byG�vb��p�t���ћ:9rj�Ǻ,�8zTAǬ�֓�F��/�J��r�N0.�������E�ч�����r��c���,����T����.F$�Gk�����C)�(���$���Oh�k�WMX[�2��q�P;��U'�������̌��Q�N���&dp�a �������'��~��]�I��Q���-z��1	�0�E���	=�h��!�R�Z>L5�l�H��@��:�wV!�̝4�Ǿ�v\�O�R�"\[��i�c�ʻ�$&��W	}2��}kpҜb0r.��Ơ,aB�r{w�.9�#�_���*R|�Z�Sn4�	��ȇ-<�Ĝ��|���a�f��}٘I\k�i���A��
X���'W�h�~�?��㺢5�=k�o���t`�&YKj�o���<J��^	��a�@ڎ'�N���!�Q&��ުt����%>ДeR:ʑ9i��?�~�B>z�_"O"�(����lw�֍ �&�1�ۓU���A�$���'[�Х1���.�y��WY��)}|�V�)B����vJo%1[����[.�+I�c���16�->�� ����*�r+��..B�"Т�Xc��;����B$Oܺ�<>qE�2�
-��5�+Ԗļw�	��	�B��(9��Ytyc� �UyED�-���/�>�{�6u�N\���|�|�e
O����v�+3YQu
�x�����yܝl���(���+r�/�B�s�~��FBN�d_��MS�65��6*+ҍ(+��-C7����" A4�ȥ�z�.I��sJFW�NM!B�d����Oja4J��ܱ�/ʰ��4i����<����H��lX_�)w]�k�ݩܵiL�w����[�8{��)>!+_ܡTI��O⏳=4���m�]x��>����wwgP�s�?���~�<T.���tqCq0ܒ1�+e�B��[Q������1=З���0vs���Ｉ\P�z�s��G#��Z���E��jw��0���Y)s�������w�O:���
G��tL儖�x��])�k��R�� T �Տ%��^,�1���B���f2�F�l�jLae�=&��%�AG��J��Ց����K\_�7��Fj��Ӝ�.�=e�>��4������J5�h����-K? (�	��a���"6ݲ4���þ����ӤnT%���@�U"z����X�c����'��q(��,e�,���Jϝ�?�3iJ�@$���W#_J��e�g���6����>�p���!D�����%�K��o�g动�����˿h�9m9�[4(%P}�/�_ـN��i(�D��s�'p�7U�Y;�!���c�aO���<TIC W�y[��;q��`L`&C���E�(�J1�0��3H�O�&���!�eiv��Mwa7��sЃ;�!�È8,���n#�C�,�r�{b|c�9(o�o���nnPIk$)N�ߓV�<�֬xJ��˞ڬ��nï�)���}�y��!��//�H5ė���V�Y��f(��=I�Eҵͳ��2�<e�'�]�i*����>yji�٫�>2������T�n�D���3������VT\��E�:0�P�4���Z	�l�L����Ъ�h�CD2��[��t�W�K��i2�c�D���[�d�1���{3��H!����y��6"���_��	5��F�W+�߭�8h�?:����M�R׭��6�C8����l�M��Z']��B ]��GC>_�v� �쎋��|�ț��� '�ov����5U%����4l�<yfZ�m������)#$�I`�_�]C5-fR��Y=D4��������#0��UU�Έ@<����A�1c�EVqδ?i�J$+gaYWLXWh�N��C)Dd�ZE5$&1~��;zj1M�T���`���O��j.y����2�,⩜�����[,���ǲl��A!�6qѺ���� )���@ӎ�INx��d��(sJ�s���Ϩ���.���/�{��-�<��5i�`���m�ki��=T#�y
]%F�uЊ@�|�c��MD���nħ�|[����w� >X�^)�|Y0Gw�h��/2�S&�w�fX&�^ԩ�9��6�"/��d(1#����r/�U�a���r�I����-�nE��>_�����/!*V�L�q�Y[�Q7I^�0h���� (d����cqP3թ�k�t�eOy3��Ӗ�:�o��J�� �y	`Q�P2>�9-sm~o��uAX��wa���:�	�P�����~��Z<���x��'{�f�od��*��N�, �w���b�.�WR�t�_s���en�0��V�g�� �Ӛ�ss}��ԘP8C~.�vuP�:T��8������z�S�~EwM�7�\b����֊����� ���6X�	��`+m�c����e�$7I��Q%e�qz?��a�~~ A�"��]�� �qAEvQ���d��rp|2o��z������{���(.�������U�?�=����_wD�o����D�~$d��l�Y������Z����Gm�a�0��t֗
�I��.p���!����y�<���Å���J��'��Z�$A4E�&�y]dc����m��[V�f�����L���.�|�����F�K~^���Tk�F�2,2�ԝ�e��%q�I��J�zi� ����FJФw3����4~�q��T��T��cF2�]e�;fTd���XO,٨#�K�"\�Cê���h	��U���V�u���l:'GC���r�H�ө���FA�@u�	,Ɯ�U�B�Y�C25C�.��aQ���M<U���J��S�ِ���3���7���Ǩ0���3����h=���1�`�I���R��	�����	�"ȼ�����1H��>@*~ ��y���K�<���e<� �3��]����Q=��:�gH:ͦ�5�0Z~�G[�x�=��j-����X�lІa.8���z<��y.���n��Y���Ò�2��ϯť��]D�EkC����@�L�rw��ϸ�� 	����<��}� �Lߴ��1? �Qe���KQl==^�/h���p����::E�b��Q���Xm��0�� �9��mYk���D:��E�3a4/��M?�fd���ۍSډ�����>A�$���_�����x�_��X�=t��ё���LP�+��20��!mJ�ٱ�j�1N��^6X�4�T���ǆkr�\������%Z[�`K���t��(�;J��8��q���|��4Ȗ�r���R��@�i*0��k��N�'Q�q^�T�Ľ|�wQк6t�Du��1�\��/��!T�!��T�BX�~UVb���k���\*yl���w���~�/�F���FgY���:����+�I���ZJ��c��m��'�WU�M!�����F�Hw2��&�L�A�q>��>L{{Xt�|J����;vZIe�A�"M���L����4�B������n�\��)5J��o��?x ��6<SPqb��I�A�4��!�Y��Ȗ��&�C��j���P�#\�4��g�۸���ϒ�啾g�R;��|G��wϺ�E�%M�0��h��Q'�v�V��Q�a�)If	���߄G����{��ͣɜ�?��M���X�)r,�i�C�Yh3�d Ez�^c_���Dȁ�&�.�����>�Xy���Bˑ#K�>�����mI���V8-�����¿
�X�� �[��h(1ĉ��1�W���^e>	����r_kn�}��I�m�䊺�2�~���Z�kP���	$l���Ui�����a	�4o�k	<ޘ,�t���WW}���_[y����-�
�w�aR��u�X�n��?>M����ȸƽ�)�l����OhA�I�T1=C���d��1�6)�K�a[M*���b��ŨVU��j�fV<��7��B�C�у��,��K�(��N;�I �XO�T�[�2����6B�̋D&ic AMP�\��S+�Ld,�\��4O.�b������Q� \R�����O����".|��!�w��}wĽ}��g3�j5���1��َ�vX��ޘ��ΛD����˫,kF�su����o_�
"�+�����_��5���?El�\�e�T���q����ڦ��!z�-��k�ƃ��+�(��)c׃�r����k�9��|�-�:,�}���vWʝ͹�� �Ҟ�&�)����MbL�Y��mD6��ִ+����~$
&��6����.�#rѾ��V}W���2�����k�+�r���SN�}6�]2�6U�l�@�^^���hV��aB�S�p�����I}S��i���0��\6��&T�2dO�M/	P�5澤a	ٟ���ߝk1�pMT��Ħ�͞a��(���P�|ܿ)o�j��,g"۹��Z���՜�IbU� ;0q�`O5P�$6x[�\�E�_�+�=�1�-���)7vX
[9|�,n���z{����Aw��FU�VJNO[`;�E�rS*����L�%� ��͓�_Px� p��9dR& �g�n�ED	�I6���;����G�j�w��׸#���?r2Q/Vu���f���k�^%%���7���9����j�_r�O�{�AW9Q"eҸ-(��:%f�,M�  D��&(���k�p�,�e�Zo
W	�^�-LSBY3�IO��Z8Ѓ�p4�|�Dds�JS9��&�5e��I-��?K�Qac⹥5z!2������i`L���Pc�:��hl���,Wqė�R�p7&ּ��b$E�@�A�!�߾��0B��?\s�<���B鷷���P����֙�ŕ�(�B�����b������]T˕c��JE�Hj��)�:�9�
�	vFǼ�;P���/�p���#��19�Y�r4�cDm��y)���8�@�l�z�>�no'cir�I�w�r�4H'��@1�%�F{`�"L�ԧ�WFc�xd�p�8h�����w��M�F�%�'�6Mh����$�a4r����2�׎ ��v
��X++�>A�D+O'��T��[��_�A�_j��ǘ:*�e��Ӭm߹��� ˾�,����xv�,��N �2b33m�-��@'q�+���t��}e!��Ѝ�����
O�Kɑ!��J|�2eZ� �krЩԅ-�s�u�};�3:��c	���p��tnf�2�s��xp8�ՊNm���El���c��;��#W��aY /��~��G,\Q����䠂���q�t��)h���4�zb�eᒠ��t�c�5��>|
M{i����a����ѷd�P)�����s����&"J@�gt���o��͠��a�"t���N3��TUܒ2��s��f9�>*{�1��L`�Cَ?Ԙ���y�!\׋-�R�띊F�@�����׬bQx-fmj{�p��MG��!��a r��ٽ	�'l��w��}��Ī�t���'tc���ë;��n���U�G�J��\� �kΎ0��)fq���t]�6�Ϛ,�a��`�N�	t�O���)�k#�f<NC7jH��PF4@i>�	�C]�DT�n&F"I(�<�H���9tB5E�F�0yI	�J�LNF� ��e+>��sfڌ����8n�u�,a��w@�w�^��{�C%��a�s�f�d�R�Kr�x�K�KEeG�e�x_�T��N�@H�+(�g���������pv���f{���m%�h����w *���6����JM2F�����?jv�����|�I@Pw�Ԯ�k�l1��⏩�.�� ]�~E�-@eҐ�ƁHŹە��u�ɬ�B��R���In�M�����
�3�h���fꘜ
;P̩ݶ4M�Zo0�H[`HX/nc(��0v��!��8��<��b���5���33XꍗC����7��G������i�����b=,M���9x�2���j[D󚕭Q�Sf�
�CW���_X�O[�����غ`�nG?G���0r{����<ù��ы���3���L�����TBR^���%�X"͛ �����J���>עm����Cߖ�1�`�7b�N�miL���d���C��nu�¶�?<4z̶��WͪxӈB�4 ��`�*8PX8���v��@�w�f���G 
7ed][�]9�A��ui�۪�Eg�C��^>�7f;�|N�'#�����`���Ze=HE,����4rB�|W�A��6�=�)3�l����R�V�G}������)6�t�8a�Z5�3۫)��ؕ���t:�8�����P6�7]�p��?��UIk��	�7�a�7����	Or���2*���r: �0�bs�.��
Hp^[��H�?��ޙ
<�� �w�������X��l׉�~��$r&��۵hԊ�XXGɴ%"`���|]�et���K��+:�l�2�q�6M_
�j�@�yZo��Cv����d�p��4�pd��.7�,2��i,_�nَQ��D:�/p�d9��BpJo{���3��7t|����a��iz�ѺQ}ݢ��ÉA0�ʢk7�>��c$2��S��=�N��:��&���A �/��y�i�O��҄��.�sƐ��Y��>Nm纾�=ڐ�Ĥ��4�k{�䟔�ڝ�.�d�$'����y>��7'�X�ҿ����LKW�3����#��JL������\X�D��0��e���� �M��C~+�Y�*�@ț6�!Tc�u���g��Xʵ�?C�+!sr�J��Ψ�S�sq����a�C��i958h��>�U�gó��E�zP��xز��F��*M+^�u?���dN~��D�� �X�N����� ��~�EM�/X5�2�݅X��.WЗ���[�d06��L��I���x�}A[w�������M���v���v�Ys�6�{|�/�^��Ο���q������h\0F
Ȁ�W�t`'ܽV
���t$�aO��Y�h:���Ӭ������	�u�bqz��\3X�rC`�#�G��[x����b�3�L�
�/�zh�d���q���8��c���H��O
�D��w&����ʿVz?LW���Ǟ	t���f�9���k��g��}��eX�q�6N5��`��YѨq陏W$�- u
�2��؛���P���Ai�P-�M-�d���AS�~]�d]�]�c���8p?#.T<l~��R�7#7#�QPg)��>p����`���NPXa	P��:����H��o��!�ϒ JA�m�-��T=�1b�j����߸ے�]�P��u�v��������n���o�h�u�l�S�ƃ%��s��k��D	7-a���V �Y�J������=���e|z�o,��ܠ4�H�����Sލ��[�����l�$]� I���[�,
�I:V_`�Y[�#�F&��Wƛ�HE�V�{ڷ*��1�?u��'�uc`��7ڠ��>́�0Y�s �#����3]�d����5�w���ЫGŒAN�AT���ɖjR5��~'�m��&{]�8�ķuP�~�{������t�Q���ZG�쌙 J�W%j{W��x���jY~�up���d|�ʹ
�;{P���U~b���ADsl#g� ���+�$
�D�y�ErR��0�*�C�UUn1]�_������C\��uu���l'�44w:�`�!8ǈ����H+����&;�}in����������>X��v�܇��F^���K@;7���V^����>�T\r�����N̏c�L��c-jW�Wg���P��Xm��z)Rs�ij��<=L`
��v��v6����=6��F��!�̣[ΐ��j
ɓo)b��(�.�8����c��ؑ(㧯5a��0z��r&ԕ��~�^�'f�ҥ}`�0��mxQ��4"v�V^�6YZ��tZ��;��"����U��x�79��!o���z��1�Z�R�Ҕ��Le������s�K;�b��4 �J��`�	e��:c!�j	�ԋk���n��H�f�M�}@�Ҥ����r(-i��7f�}S�S��EK�Խ|�)��еy_nY:nP�[�t����1^@!R�;D�4쑊��|�Sk�����	�MV^q����G��l��Q����e�:�KwT�h棔�,.�ޚ<�g/z@�����R��[P��=�ó�����nn�po��4�VrD����\�b�weUQ<F�� �\=�[����=Y���K�׭��TP� T\�����kZ�:��cc�匀9��ɢ7�Ȑ�ܾ����M�Ý���U�����[���	iؽ9:i��DȖ��P���W���B/*�_e�~=iݨ4䱆�}��{�"N��Ҳ�K�zN_7m�U�p%���Ǥ�/�,������,n�+rF@�h4��=1�H2��}V��p�t�~�%�P�\D
��޼�׾��3�p�;�f)�����̙�)�)wc$��:����nm�`nY)�GU�;�SW�x�ݦ�t]�\knc��)���P4.��7u�����f��[�\�����*Ԩ��(��L~��g]��5�Gr�����BY��V6ǛIn��X�C�Q��+h���<'��8O���G�k|Ë�u8T�=v����#lg�y&���i_a��[	�!��0U�DW���i���)՝�"4`SӼѻ��Q㐖�gW��	�����ul�X]�͡���kUe�OR�g�����	��e.�SVG��4E�^����-�y�l��^׹~����-���b:�I�rD�#t����4X"���
xo�'�;��x�h�����P��KT-�̭vL�X9plݢ��{��:h�Y'��W-^�8� ��#aO�-�B�������(��%��)�+g��O �(A
 x��]H��Lʣ��'R�a-1�K��k�4� p뱢D)�]M�p+���f쥓ĭRyJis3�M������Ē_�e�.F�̽�/,�[F�ţ��_�Ǩ&���sr*B�
��Vr�������J<C��#Z�!����شٲ�ǻ�I1� �o�R��cIe�^���F� }��(��Kh���hRKE�/ؚ�Xr�6���6��Ԋ������{t]ؼM��� �X�Qτ�U]5̧�O<�iėU�Mv�]�@;_�p��hU8a�Uܧ��u�R�WC�� �TE�4����H����͹:)4���<y���#�Em�*^֖B�ӽ��~��w�	hݖ����K���-��+��F&Ox9���� ��@r�íG`^��~�1�u� ���R.���H��~�]<�й\��`'~�C�ˤ$��d?/J�e@����>M����X�I%�u8�on�Z�	��{���guh�[�_�-"��Uw�����qw�����ዪr9gw�-([�;H�,���O��� ;�?�����]��!��`l��:���	�M��f���-f�tLR���ǁxTТ�rNĜO�������zD���C�?7R<�3��給��x
��<��|7M��� �bZ�S�.�`�d�����cn�E$��o4CtP�X7\ !�[������4�{%.֜�J�;I����|%zuD�^� <d��G��t�������a��y�oL,Gꩫ��屻9��۪㫉�-��^J���3���stz���e�4c��0�Z�&R0ɷ�9� �i���B��na����ˉ�3�����0�{��݅A�?=*�,��r!
��gƵ$Ǫ�����&,7=���B z�m�-
z|��A_9G��'(���ng*7�s�.�:u�8���I�w��8E�Ӱٚ{�4<2��y��B�U�~��0��͘ůl#�M�J���i�)Io(��D��sK������&�G��K)y��Aa��5ֺ�D6b��}
'vo�o�VՕv��.^�����y����G���r����
 nN��g���Aύ�S"?��!&�Z��BF��fܡ���s-[o��	�'�ޣ!-�,� ֯�_��lL��X�[G��$�l��v-�9Z������<���Y���h̢v� C�&� e4ps�TF�³{�@�6��]�
W�5�<�{�����v� C�"fn?�H&�x��*�|X�ɰ,�al&��ؙ>�(tǽ�~9�D ��u���{��e ]�)�>'��0H���%� �[��i����E(pxPW�gXJBO��hؙ9er�A��޸������tώ4������H�%��+����>f�V��L���S���"�*�҃�7zUL�$��[q����HYc�T��[������yM	w�����2o5W�*���Ӂ?��O{�yȁ"G`alupR�*�FF�����/F��kǽ��R�V�<����jڡA�?@gM!�|��4��~�Q ��W�8ǂ`P ��6�ɯ�|����Xc�`�2�{����q%ٜh�j�
,�Ez����]�Wg����v��}�I誢S�W�S/��R]d�2�\�([3`��[v��bȲ�E���m�){I� ���~�)��~�mIC�&�a��r*к��?40a~��aRߐi\���z���PٿWi�d s=��(p�(���b�o*r�4kz&=���$��Q� �m
�K,4!4�>T�f����d�zR`��@���N/��a��E��:/��k���3(2��M���`�%c/����*��1x%��D,��7�{ٓ��F>]0:v�¹�_IJ��ж�R�\qE�4A�gZ$@ސ7�P^�b���lʥ�g���De_w�Vp��̧J��:��z���N��3�s��}����B�:����6��(s�3���^����җ��	���� ���zyQ�3WQ�fw#�'�i�ew3v��[��3��UȢiN�5WQ�,���������`~'X�bx�{�^���(WL�h�j�-�̒��[Y���͸�s�I4��o�����������)L ��� XLܣeLApI�h��R�~I�y�,~új�[j���	_x�O+�0bJ�~��t��X��Ǳ�:�HӘ��5?������Jj��#*О�1�::����:��9M��L���f�~o�h��<͆è������Y� �}Z� ���|.8M�G�R�/A8Km}"�9'�\޹���Q����hk��_?
J�l�x����Ի��6�a���@[�q*{�#CDF�%oՓ�b�%-]�w3S���_�%ľ5�u+
�Ne�,���R$.�x
WLEÿ�"'bM=6n~�n��t?����\���߯_�����8�Vp1M�W���&�oZ���G�\�.�: w�#����`���o�h2i޹%׹	!�`܇k�䜽2e:C�,���&����n2�%��@}s� �1Q{|��w5�|����uUR��t귲8]���n�:�G����}���ŅaH�u��˃Mx�r�F�z��ۣ>f����9BW�b��v}ҚK݃ҍ���N��i<���OC�����8aŷZ����G(0������}�"JQ,�
��׉��4�I�P����丳:��D4<2�j����Z����h]��Zm*�ɳ�D������_�&���O��ʝhB47�i��^��\q�N�2�Wğ7��Hc��E��7�D�X�in�}�������4���
&�z"f۫�.�#��Ŏc����QtoG��䵪DF����o\�ކ롉ȹD{n�	:�qm*�}U��ﺨ��M>.�9pZ�3��Io�
�O�H8���Y�-e����g��W=q��,��Kb��ұ~�����|�ugY]�^�O�e��_1%�4/�]`�K��g�'�~g�ͤ8$�p4D�����-��hm|2!�@�0[v"�G�H- ˞��i�Zi7ֿ̀P��BK��YӡL��Y���׋�"X�K��ȅ��U�$��\{t@No����ɗ:v����QR�;�v]b=���F��`��L]�S�����aG<��;�1�=�`��K9��
[ �x*�e�� �D+e����q��z/��5��hD���Y��V)9�qZT�Hl~��[�h�'�$�f��S�jcń5���gۗu8Z�]�]��������p��$�g��G��*Sh�-�"t4+�rM�����%���ZZI�2�3�ڏz t�H9M30d���� �B�au��#,,/ Hi�:��J��V���c��
m@�-Oo�T�)�=E��h~���G�
h�e�5�%9,`;�a�V���a�F.��>�I�L������=�>���{Ԭ M���P�}�!����(
�v�����'�ć>qa�<jI��%�1z����
�@���!`K�G�(%T������F�j��Ü޽�P��@ڪ�\/�r�<�)�U`e��-&w]w�;>T�kޮAʰ6m������>S�h���M]�T�~�.D��98Ug{;�C��|0 �گ_7m��~ks�����}�(U٭�� �"	,���<�7}�T�����|��rGç�.��Ó�읂.`b�k�q�O�L� �
?zp���"w��[�c
��X^���{�\q��6���NR��Cz1��?k�{�M��ܽ0�K
�lV��@�d}�6�a<�"�"� �H}�ǷL?�F�>��R��9�@�G6���R-݇>����|�B�����!��%�t:af����iЇ�g�B�h�ǟV��v��W�޾�\���"�T'�+a��"Ca�i���{�=ty�y4���8�s������
�\g��c�S�_�#�[���H5*�\@e�����G������;}&�v�Qi��0�P��
*��7���M<^>C��=�g�Ap�c��i��8���E_��A�^ߪ,��oR�c�D1� $xA'x��ȇ`�z��+�`�G�sF�e�F�E|����!;�+����r��Y�aJ�I�w<dB��|Ԅ�W�;f�v�z{�*i?џ��C��vf	���T�;g�ө_����m��`˪2tE{��t��~������46��U�M�>�Z�A<r6{���*��qb�T#J6Y�%�m����-������P��?�T>��[ �l�8��^���e�N|���p�/Ů���<�O_�A#��\��Y��1Q�]�ܘR�B���a�RB�l�B�I��8v2�p(��9y'���i�Ӻ=��22b��0�t�mR2�أd��AL���)Q��V�PtA�0 �0�~�mpD�ZD:ғ&8K��sd���E���(���"�~>B堛f2g�%f�}G�1>Bޑ1���vLV`Y`���B�ĀC�C�xԘܔЀ��Y�,��-��g�����ZfōL��v%�o�
&.���hҒ�=��i�a���F�k��d��X�=W�����=��Z�a�h</j����=�awy6ă�WO�Ǐw��q9s�[6�X`����fo�6Y;� �7Ot�Š^�|w
m� �AT������6a�c �����>�(8�Yw��u,�� B��+�J�.��Ys��AC��u��]����M6�N�</X��yZ@���D� �ࣤ<3P1exɉw�5��=-?��ӰJ�Y�!��5�?���hH#%��*�4�v�J<�M��(Dv�ً6�������~c�Р����'D �~�|-"�r���,���݂{��� �h�>�\��f�#�R�a4(�� �Vf�S#����dB��t�5Yʶ���n��_S }��j/'{J�*y�%{�<�G�ld�]�.C�~���18%>��"סk� L�i; �X7.\P|y�V���c�Y��cyo��� �6V�^9@�:uY8� ��".�
B��Z�C���0v��`�l����i���9B�p��f>���m���u��1Z�)w����	����P�z�.�ly���%H���Ӕ�MytĹ/�S��ǆ��nO��(S;{�M� >^�,P����'��{�È���[ˬ�YP7�k	����c�� 4`ݟ�Cلl�\T�T��0"��Z��01XS������ϯ���}vq_�
[`�*t?��(�g&.5�N��s"�x�:��� ����""�߉�ߖ�丬�7C <�`:hc��	��d�/��9�b{�N��,��C��{���R�:K���g�,�j��l�3�7+����^�1ʗ��:�(�'@�:�Uu�
�� ׇ?$���H���)���]35���N)fӪ!]m�|1&�1x��*�c�v�-�	����-Z�2 S�D��s�f��Um�vR�DS����s���,����A�=�xWV5�w�EXέ���V�����nq�D�Gx�ꇅ<e�4lU��yz!��PZNp�J��h�A�cQh�C���N�N������(�����wG�t�U*FP[�aF(y��?�8��Yd�+E6b6/���7N���r��V��`!&/������Y�T	�#q���Fu8ɫCiFګ0��ݣ�^n-~�D���:_Ρn5���^��	�����Hz�2��~0�/}�Ƚ�h
Q�%���jC��B�� ��F9�X����(f$�'����'�,o��<���2&�'�}�l��Y��,1��'�g�=~mU�'�~�+�)`kj��IWn�4�c��S2��ߚ5���n~*y��;=�S����jʕk8,�n��.��e�EC�ٓe������9Ӑ4�gB6%��n����Ӗ/{�0�@�m6 oĖ��!�^Qj��	�@X��bY.VM=O�������c�z�[����̝9��g���:�xإS�?R�jO;��g�]�ڤ|��:p9,����d�&�#��s~�:�h�ZS&�{����ɣԞEM5�0��	���7���2(�3x;���w�K�.2���o�x*{ߎ�Y�t�a�|���n��e�BW�-����+K"�=�HѣC�����W<�u>�HlA�RK�{���-�U�z��;��8�¡��]�*d�[�{��
~�V��)�"ձi[�d�����v-�� .x�~ D'D��s����5}��M[������T�D�5|G%�z�M�V��A�u#߻��|�ZL��D����Xː���Z�5��Zw>`��;i�J&QCg�z�'��o��y�w���ɱ�@9U�d	��8oE�Z6Z1n;݈��n�1+���N;����c����~��<�i��2��W5�����o�N��Z��T��`�4�C^���4��9��#c�к[{M˛�����;�{�ڮ�42b�) y���I^��׿2�t,!Ӫf�KьV���d����q�ؗ`�MY�tm���˪7�	�$e�:</��߂�C�a�_�y�r�(٢"�#�輶�)?�֚2��^�n�z�|n�3t�+t�u#ZǸ�F��LѼ�Z�/�_���/ YI�%hhnN/��'������*̤��˟-M��Hv��]69���z���O��n3E��{�����g����!l���N)l$�RA�Sc��;�bu[��U��𼲆�,���+��|����K�x��U�s�t	��;�`|S^���v*��; 0z𿝦M����K�@W��)�ȇ��ku$"�p����Wd��������U|v�Y��^���*X�i��<^�����v�W�;�G�����/�-�H��W�&��-��t���V���6)[P��@���] wH$�H
'�O�I&^���!����6�&�k�Y-�.���waYG}���SD��$!)�B�e�>�4��|���᱄>R��Ǎ��4�+G�AY���M� ��3�f�f�p ;�?��t���)ݸ�2��>;E8#Bft��;��B�M������EI٩b�.TSK�]{%]�qKî��;�ܠv$%'��y�F]Y���3
!Uj9,�O��4|�~���[�����⾘��z;��C�Q[�SU��8��e��a�F���	d��f�\%�9�nc5n����:�>���MoEn�cBnL�v�Ks�k�+.f��X֭O%>wS9�!�}���2�w8�y�����!0�
Bc���}�^��.o��u1X_�Bg����,#~��Vx��5���; ��g�~�q�����g�'՗�!������E�n��(oE��� ���XZ�(��4�����Y�q��v�³/�ۊ��Ki>������X�
f���Z�޹�����SQ3i ��h���~����ui+C��s#����C�
�s���I�p����qSdI`�Q����Ds��LWS:f�Ks.�y��}L[�Ŧ#��������A�S�>m�/_"6P~�������/�}��2cU�4�����=�y�=�7x��#��K`������;��듾VOJ0���l�+�l?�f��̿�f*���S��)��i��ܨg;�)�� <xTk����1�Qz=Ҝ���Yp*%�?;���%M~�!X���Pڦ#`�Z��D�O�b����8w���)�$a+���3�za	d�%[$D� Y�1��wvx���bv�wWy�e'��t��ɖC��������p_jݷX0^G��}�=��D��¬ ���q�B�F�{i���<D�:zf�yw����|{�\�#��(�гo�t��p���h�����4ci�n���A��
Ǧ�	�4_��*�U=����*�d-f��̡ʲ��M���
�ow-���Iu�E�iPw�ho�((�>��n��:�D�<(T֭k����F_ ���L�H�%��:8Vi|�Ә�4a�ւ����0�}:n��1<I⸗iO�&LcjgH@�G�:�e�7�i]���#$W]���ظQf�C�Q�Z�=�ѶŔR<�`+������N��a�6��f�|6H����gF)���u�$��YZ��`��+��ط<R��ฦ�pM�0A��Rn@w����ʁ�.��De�"y�h����,�T}���}q�7}n��7�X�V3k=�˚�I��rԯ fC�4w.��6��0Z?g=R3Q�[�E�d��ҽ:����j�:��F{��=ʜ��[~�No�6����as�N��X$�O��4��@��� �
}�W��&S�y��TbqX��8��]�=蠣:Ë�a(Cx �ʨ��gicE��M���J�Q'�;�z��V����]g��:����Y�]s38(Ÿ�L"*$1B��
���_�8��*��ɟe6q l�sx)&u�H�x�#/ٿ������U��XKV�qZm 5�D��h�S2U��V�2�hlԉ'vz\���������)u�ʍ�3�0�e�6`�7}*S-8U~փ�Q�P�8.X�8�����9���d�����vf�L�����rZ��{�+y��=Z@Fu��v�����yC�r��̖NuŔ!�JK˚��0�哟���&�(/�K3F	"��I���<i�a�/7��9��* �SP
E����}�j�`*2��#�O�������sKi�q� �)�0�km��j�9��|K�y!� �mxG4��c=Äz/*P�����.cE�|��������ī��x"w5׋-n�d�]���KF�z��yG ������)�wp?���F��l���t��+a��rtO�T��Ӑo_�ŋ�5 ���-Oe���g`�\�����B*�*<�~�X7>"��غ	z�L�\�?z�%��L{�dxwF��$Iy�}���:;}C*el��g�'�Xi���Y
7�ZoՋ�������U�Q��χ�츨L5&����un�����P*�=�JT^*=2O�X7A�؁HЬv�{~��r����bd�b>�>��f���Ql���ێx�G�~͇���7�ش'y���ǣgg�N8PJd�Ü�:��#=Q+4K
��#����F$��H�
;��/���8(UU�i��-=�쑑�y��<l�k��K�|���J��|�oۅ�55#�-�By�G��w7J�\;zE����@��ѸP(�\G\5	�u�u�Ўޜ��e��tj�)�?PQ�{��jh�L�L�j9�s?l~�悇���f�2xs��h��8E�TY��"�.#1��_-A��,U�+��a~+�~�V1ۿ�o����k�_�z�A@�=x��t�S� �>}4�f�27�L)��5z2\�)I8�}����c�!��)���1��-'����{ib�z#�F�=X�&D�.�Ua�b]�$���t�=mb���U'��PV*��N0#=Ru�v��-d}�2(��A�o-~ Q��b�5i ��Y��m�0/�,`��.��oK��4��D��"XviOi��{k���*}�h� hZ�qƫ̩o����&��Wl0�����L�Ĩ�^�}[m�����*�R0Ȉ^ΏVP�5u���{_5��I=]~Z.k��pG���G�q��\M,o��i��gr���[ �x���y���&�< �>���=��pzԿ��4���@���������]�ϓ�S�8�]�{�����ҙgl��#C�ֽz�|��	������0e�1�� �i�^�	�i�-��;l3���~+ko��J��Ʊ@��6Lʯ�i���kZ@�louq4t����'g�]�W�G��"��Ed�Ɇ�[�s}�R��a�T��B "��vM���1���+��+��hB�F�H���O]c^���҉Hsŋ�C��	���_P���~YQ�+�}���ڌw3Ar̝�������+��q�3\���'�?i5�m��g��p�c�=�@}מ���@�������,ť�vj)���Ω�d�N���'���I<�w��Z��lR�FB��Ӽ�W[$�Eh�$��(�ovr8�&�P	��.��Z5R����eO�������M�H�e��%��W7����K�5�:�O��ƌ���"Z�<X�r�,�w��x@���5� e��L�O(9���U�ۛ7Q�����׊�_�*RcC�_���g�BW;�*&�]4p���`��(�: �5�p'�"�������!!�fQAN�l!�߹�.��R�>���k�a�HX���{���:9�0LU���=}Zg�d�Pit��&P�q�_�Ү�����ӆP
�B�'V��L-hV�} �F�\�86v���>��),��=8*cfh=PWSf�j��h ��;u���� �yV��R�H�����6��)���jޞ\l`�|_9�&bH��r��!\��ڻtjvim�X��*�"ZYj��'Iw�l���!�as\��?j\Kr��|�%���.T�\��&�s��Y���F"����dj���Z�ӹb������H��y(+G��P��w�M�]�?��m9Ayj���Ba����<��G
Z��U�n>���>kQN�0�=Gm��)�[|��r7�Ǯ�)�,U��hriC@$i��Hd7��9z����sA;2��~݊Y
�d%�[S�q���*t��㦖�17��~���.V��SּW@�	�VC�:LC{���!/-�640�ƭ�K�Σǟ-�Z+'sg��q���bv�k�Д�ݒq�fD�J^-��W��R3�z�}�Fj1>���\
?	��d��x+�B*'`7Μ����������(�k�sYÿ�@�Z�zO��@��R��H�:A�%.�w�Ǿ��р^ZT;�u�g�[{*"K�U���Hθf�WÖ!����׳�m2��'R�w/v���˰1��h��@���^�L��V��C�_'��(�)*L ��	DoS�y�u�S��j]��!���� 7_>���(�"�n>��S�y�>L�F�Wo&Q������L�c��h�*�RC�%X�������?�_t��m=�Ex�W�U"��y4 �[Q9x�)�}��@'9x.�0		�����HBX��q@���3pɊ�Zzw�Buԉ�e�?̥���4��+��//¥h�g�Z�(�Qu����H�4���4rQ�x|�h��z$Fb�x�w�?�.���-�c����"չ^�P�ݻ��!/Xʩƭ���|' |�m��|���ʱ)vh�e�)eD<�`�oMi�^]��\�g����������Ωȥ����xZ����S��K���q�� b��ޚ���!d��bD�OYe���X�F�n(s���D~�[ݲ�bCun���<F����£��!�N� �>\��W�1IX��)��"�b�	��K�%;��E��ș�����x�SX"�)XX��Q��F��}�P���iI��I�}�fM�n��<7<�/��8�V��J�����k�f�CvM("p�3���U�����Pފ\ד���ރ��x�������N�i�xt�3L�����,��������r>0-��f;C��͓�-���ҍ��6�!�a��s�g07�h!�h�
H<�e�����:�[�U��J�W�ܒ�m[����y�n㡉�)�??���	L�m �+��zMF�B,������.�T͜hr��������[�C�|�e�ە{ܽ��N�`�+�Fa՚u�w��8Uҩ�����#�r���ɰ�$Z~���u:����*D,�>�͘��ԗ,T��x��q�{���7��<IOq?av#�Vl�O�,
�$U���[��/��ܒ|ma�`r)'����(���yB$y��
ۻ�+PZʺ9��v��?oAb��)<����K����o���h4#�
'�y�=/�=��0��й0��_��6&.��*]�8�������e*�[G�f���f�z<��[@j��!���4�O����/�U�X)��oTAQ��@~M}0�uD� c�LI�[���(c��2�E�^r#�\\�P���n�J���9ҵՇ�1](^��N�i6�K��`m^��Z�OC��9�4y��ވB�3^�3D�2�$Mvy�7��1U��`��,�4M��9<b��D �k<�=5�C��� O�y1\lX���v�Y�>�գ`f��>&Y��ܺ!L=@_�Z�Ĥ4@��Gq&D��[��!ҩ��@k[�(j(�85��L��;Չh�n%ċ���}��m�K*e-���D�����b���!�r�x�I��rH��T���X`"�0���r�k�9�5���jg�9.��M�]�$=5��������y�ʱ˸ˡ�]��"'k'21[��Üꎆ��-�\��W�ӽ�