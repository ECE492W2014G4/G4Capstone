��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+���]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�O'�yz,�_ ���)ZN�6��dQr�p�x�y�C'�m��H.@'�!ѽ��Ќ����M�����9p��s���v���	a���y�A��n�M�1%�P��Jl���� �k�
:�q(T�F��l�F�j��;*Sc�e�op'Ho��$��'�*>��e���y������@�%X�9��o@����&RY/�~f�C��31�qĄ�J� ���2��:<��-��q*J�����>+e�!1��]4q§ �]m�ԫZ����v�����F�q�S��8�00�F�ړ� ��5���5����Z�Q�!�&��^�����'Fdf}uQ��z����*��>1���	��k.A_wa���Dky�G�#�,��*W(<�����%����۲Ȇ�������J0i�}6(�� ?Rvt�=�8{����dR��冖�kx�BZ{��$̐�,�?AvvR]5�Sڔ�\�4����j��>,�5>�-������E=���Q b���k��s ������c��Y��E�̒;�[����5������A�k�R�U+IM�"�JGp��w��Q*�|H��2�c�o��MP��P�W�-�0����9�Y�� �~~'A�wёO��/�ϧ{%+�)�8�B�F�H��l@.��Z��!;OJ�R	(� ��P���P�C���^���J�yӵ�����)7�ߦ/�L�������vO5ك?8=� �$N,�N����C|��(��-����l0M��Hs~��d�#:/ ����HjAEMi���~������1d;�m	��ԢvO�|��H�R���v�ta��;��j-������6�,�Fj�Ͽ��9�Q���T>*���	��B�\w��������!*E	f�z���݉�8̬\	�v�ܥ�Bf��PO5d�9|�.��e�E�]��/��F@ķ[��՞�Ƥ���RXYb̹�}�4c�:{�U�m	���	^�.���o]b��BZ��E��V0��+���R
��6��������פ���N͛"��O��	��F�Z!ޢ���Iȃ���B���0� �����J�T�2nu�2�M�)�!ł�n Ŷ��t���t�����M(��'�sg���g�]j�z�ɿ�e�얱g?ջƝA��Z��: ��AA Y5�f��M2Um'(���ρ��R�e�1����L�<vU��e�&TD��9��H)�2�V��{��%g��kl��[���)t`�ȣL��ni���8Ж8
ԓ���KS���4��&6�������4���~��`o<%�!�qK\_< �8��.�l��u��$a�v���i#��_�0��c������
�S�GV�ْ�	��k��vT���0jZ��#>��ćW%�32?��m5�kB�?]+��V{:x�du53"���Y"|�>�Mny/L� |��c� wM,k���(&L�Z6�X*x������U�IU��\>(hW$��M��B�Sy�0U��w�)��_[a-�U��X��y�V*�����T�.��~uK84BIf x��H�?���=��M��xU�&�fc��b:y��6���(�ޕS�F�{��g#��e���Z�㸎8ҵ�n�g3qD���/�ĮY��۵���kk,Q�����U��|�]���B���K� Wt�u��H�g�D!��>�0�����3|i�:��I�c���#��
�J�[�'������І$��-�s��p�AW��Qr�v,H�8_D��iɓ�5S%�6i�Ǟ4�Qv,d�^����[L<�ݜ�����t��gt�� �lբ��m�3Mj=-�ih?�e���S�ƫR��n8tC>s��j�jL40Ȕ85���.���(����4񺉰*IS�xb�b��*���.���uT-I0�Y���jR��4�U�2Ns�q�T�j8Eb��GP@�����R�x����H8(��"��Ԙ1gK ���{���v�
��fʺ"���xV�5;H g9+m�$y���f@baD=�@��B�P�����ĕ�=,N}����x�<���k��V�cm�˔Á���F@�M�����M�G�J��@w �pH�o4�4�E���Eb|a]�x�-��qL���j�Z�}4��X��6I$��G�$���ՁB`��w�w٨��xS��J�=�M�����;���s5��_�Q�u%ԥ|�Ǵ�z��?�R���Y���ua�Qo$��^{2<�/����0�
/J5M���G�Z`����Xń�L�m�tmv��hm�Ơ�t��9x�!���K`TK,�Ad|�M�^3�T������",ep	��HX��4�ned$���e]�ن �2�6U%�����������gI���3��Q5�m��:�V��Lr}�����#"���Ꮶ 7��� �[�cM9=��H@�_�=,%�NG�YMl�WGp�UoKli����Zy���r���P�����EH�3��K,�g��<bɌf��������~x肥D� �{+t��=HN�yQn4�c�K ���{���M�)�h4���2��a�̀�����#&\��<��Er�:f�d�I[�B`I߶_�X��
��f*KeB��6��7���RnQ��*�NNj'pֲE�{�>��'��b� @7��xpt�xM�w���E��D����~�=˿��fpYKTt��9�b���\���*�36\���l��h��MB&G!?u*�.�:�V��Ë4o�!���u�A��@+�J�x��5Vh�+�#�Ta,���{(�%52{�w{�I�/(�ʮ�3�ʂti��j8���c�97"�����ʘc[Wb>-���@�9�H���_4�ܺ�m/�>n���d�hraP�&�j�0�
��kG�d,e��8@�� T�̅Gre*7Au��S)j�R�]E�;3����������`�ͷ�E�l��)K�
z�6m������������H&��q�;����=��� 9�a�Y�9
��g�j��k�k`p?�:��:����~��4`��z�h:�����
�e��ޜ�u���&6	-�t=��w3�]t4���i�j�gw7Ҋ3��F��F�笰tE��[����D�f6|`-̵ �����p˰�Y�8�����UK	�hP�~\P	��:PĻ���V*4|S�Ξ�R��Y0��ӕO$@��;�����B���ߓ|b���}�ǂ�|I~I3��U�^]�,�����f[jS�lO����e��u�Õk���8�s��f[�l_�۽�"	�P�A�2c8�,omA}:�F���ف\7x�#�[�sXi8�Gj#�͕ڑ���V�.�q��Y���j~�@\.:"8��;7l�R��?]�%7�M�ڨ��^,���B��?��ڟ�s�^��6k��������}���˽~ d%��ۢ�|��S?�'0��IzF!\��Ț�LL����	8�+)�jz¼G؛�'�Zq�>0٢�d���izɼC�)5��<m���gM�h`�{׬��3\�E�����O
�0V@��V��I�r��������b���3U���WJ�m�Ӗ�D���)���hj��3��EL�z�����"'Z,��
�æ/QhMQ�oa������.��g����8Fy\�S��a!�� �>� ?�X��qS��v���8�xw��%�v��S�q�i�Qz��>Qh�	��t�3G�O@��ğI_W�E�J�*x�G͑E�P�_U�v�Cܞ�LWh6٫�sq :"A	��]U����2t�[J|�I�[^�[����p�ì�@��f";嫕�q��|b�g�7��y;��Iw+n+��ҵa7����pkM�/�e69�v��nġ�A��*A&�fԅzN^is�0|��r�s�ֽ�a\�����>.���鴗?��(����+��Z��!����y�5d]�t���gt�:�2�9�.9:�p���o�c�oi�����ڙ��fco��e�����#�H����T�?�7r���_�nV��j�(+9!S���OMY�^�wj�V_�iu�0&'@A��R K�JL�~%��ۼ5x���MU��N�E��48�gY&k�.!-�6M����x�ZQ*�����хz'�<q�-s�%��a+���<5wC�\��E$S� ?�玪 �E���]����M)|�ub>�(p�N��{���M�w͞hT:�.Uo�'ѡ
�	�"Ǣ�-���R�y�u� ���1���b���lm s*�9��'��,4����P�7�7�Ê��,��z�������Pp�a�d���[(��E�=�%ǟ4�:`兝?s6�UL-�y��@��E �^ )*����D�S8z�A<Ye��kވ���
�3�R�Kj���I����W�I��A���a:`�~����-�@�Ox+�/�̸��L���C�#�8��z�F"߸���7�Ҡ�����?IO,��L<��ۊ�k���}�|J��t`��	,�]oKI��bzK�}>�c��/͘b�j�b�[�����QI	(] �)����P�G�^�&9��q�,�Ӕ��	���U\0�F���`uYo����V�1�yY�R[���W��v��`E�_#�0���5y�'�(2	e�1���	�x��o���5��nʫ!�B�u����K��C:Y�\լ�'�4��K,�OY[fW,�e�Y<S��tl�&ɕ^����a�v���	W>>���?�n�B��wi��>T����{S�i�Z�wgE��m�h��,���X;�N�,��V�.�l(�t�PX��O���ռ�ȅپ�`?!��(��"��������J�;�N��+�����AK8�j�a���;^n���6����jzց�s�C�k�d����ƭ -���p)�-^�����V�	1�W�uxw��"a�DF��e��`Y�:{o��@dU�T�}@Pf�Rk���������׊�&�eJH^�	���N���]Z^^�r�i���a8����)�$�m3h��DS��W)`���:�QZ3KN��'��Q� �@���F��_b[��ғ�E����_�ѫ��
2��g!�Y��zo%���L^/ݽ�k�t;�uL�UH(��9ڣv�2@B���0�����E�|92~Y��Ѯ"�9��>y�󵻕�V�V{�`�+I"����������/���x��]�D�^B�x>Kdx�n����`���r[Ԯn���<97Qƞ'8�Tж|[��.��QVH��b���H� �>;�i�b�U��gmܨX�j���	s������mѷ�� %����3t��״���=.�N���!X�`�N!p��Gȩւ��H�W�%���:�q�m�`D�ٶ�6@k����cM�*�޻=a�G��|��P['�԰C�yU-v�Z��%;����,6�Ӓ���\��?\߻[�}E�PҨÏ��
�_�i[�"�E>eu���!R�	&�=%�h�.�~��7���H��VbQ7N[w����'ɒ̕��-�`��u�ǋ�A��6��q5�YM��3�<��B��cz}�EM������K�I�a9G��H!=#�{=�}�z`�J���ܥ8��{�t����K�whYh��t9,��e}f�Sz9v�g�WVb0��7sa܀���仍�������ߎ�X��0�}c<L���i�T��H����M��8�c�_��,��9��1��V�;t��=�[r^�<�!.)ٳG�v�5
W��q�1-�&5�Ǵ�a��+n�н�#��!�������	P`��Qj������U��Ο�2��7�de#�3�ﵙ�����v���pu3S�l	�������t���VUJh.�YшK���-6�TsF�愩�c-ݐ���#���rM3À�9��\Jԑ&�ຈ��h44��0��-���i�I���5��K��R�U�Aʥ�Sn8����eE�>&a@ۻ�k�y7[jIqj9ͦ���&��v�@��#Nc�zW�w�DS�Y�A�ƅ.0�wɵ.��Gj�&�z�z��
A<��B_�p�L�����C3&�f�����8�!�xfZ�9��<��bb�p�I5�X���C����̊+��9����b���2N�	B�G�B��^�*\��5�D���-�Hf�{������� )�
��b�=K��INDo!�oIj��)�����5Or~�'�B+��.#/���x����A���K�(prz#Nj|����g�=��f镥�.e��)�^f�&a�:G_�N %�ȱ�Y{<����$.E�N����'�o[���+m�w"��k�7,��c�-�"dPHn����k��V��8���+#�/�����Hgc�K/d4�G��NBF�N��N�Ա�������d&��yI�Wd��#|�S��@�̒qY#��G��R�u��v@JR�ՔN;4-� ���ƌӨ��F!�p[�id
@�\�beZ�h���DPP~jEE(���)sd��K��-"5�@����5��*C�@��@?�-��0됶G
��YրZ=Yէ�c0��嫰C�W`�7��$����Fj��8�$���gK�*�@�нͼ̅�����D��5��?rS�����^ v�"2�li�^N@)��A/簷���׎Ѱ.�wT�����5}�5F<Ӊx����3���u�=�

 �]&��6�ʛb�TD�x�`j@Uݯ�����b�M�4���TM*��9�ޅT/-��k�~�;h{�I���>�J�1����U��Q^D�Pp�r
�~��ًw�	[��/"F
��X����&�N��
����woߟTSZ�B�N�(a��~�!dٶ!4�M5r���v�
�E��\�h=s|�7�I���>�F��v�}`��	�A�򚑷iF�V�r&�̄���#���J:]>_0�<��Km��9'N�.�3d_��O���8U������~L����f������g�X��8�Yof�u��@"[3 � n]��ـ?&y�� �<
dXA!&�-)��6��7ChҴϪ U��`��W�i	�1C
�^����fӴT�����+=��6����Yc(Q1&���Y���[�t��C��)��7�Y^*�cl��3P���i�e�O�#շ<F������oS��8��p�i�,bꐕ^~�#]��+�;�OJ�WV���8-�Ǳ���~�A�x5Co��T�1a�m�"6]�b��~�k��WGm%Ǜ��6�oJ�X�������Xy0yuk�rș+!J�ɶ�)T�u���J~�q׏1@�%�LO����c}R[�յ�#0ٔ���v��<�&�˒K����6��s��B.;�H��R��K��RT��ؚ�)m�������I���1Ε_d�E��oa�'�z-�ܗ���!"������f��*o7��ޒ�G� �����]�������.�j@�P�q�y�~��a:�f@w���K�q8�"p��<�A=�ŔK����/S���������aR���vV��嵸$��tB�
7��ܟ�9׺�	�}?�SGA�Rq��BO�s����*��*ˌ`(�����C�r9���� ����!�k`����\`�����"ܰ_�������N	�|�?�mGj��Q�AG��ES��H����}r�1�tEIQ2Q�_ ��k�5m�2�|���r4}��\��p������cq��,��W��/�@}߷/\��_8"�!�m��o�o��_F��}k/����#@�+Q[�������$X�J�?�{W��b�}o�I	��)=�OψV\-�[b�e8��Se�˴j#�c�J]�O��=�h��X8��x��ǽՎs��U�[�]n�,`P=��S��k�Y+0���)))�e�|2����⋞�ͧ%���縔�����"��fv�p Tdb� �����,��Ӿ���!�P�G�w�uN���u7��.��6�&� `i���#
���}t�I']Z�Z^��n;8v��T<�I�PAb��h����Ӱ?�aW��q���"�ޟͣ-Jͺ��A&��A�P�UH[�������@�#���Ѷ<e�dt���d�U��7}����s��D�\���)��y�� r�@�M���6��� 8Y8,q�-��O�.�.�JNVr$���eEE�<��h��^�춐�Q9&�xk��$Sw��Pu��{>�o��P���P�6Rm�����Wt(�=��ؽ�oLE���,��t+�wm�6_�G���[�%�<�l�t�#���x��_b��3���N@�hF݂c�z�jw�a���e��	�}F�������|P�^W1�mn�����j����jR�Y���@!�B�|��߈�����R�w}ցZ̳[����(��6s�m�M��Y�_q�⠝m(��
uO�R[��D܈J��Յ�`�ă�)ƫ�"s �sV��1��֖ZZRT^u�ܥ!��F�4>�ˆ��'��%�����:�Bs�]��t�~���3��� 8��P@�uH�!o�Y�=�q�c,ֶD�G��i�&���/�.��|�1Q,%�[�j���i��Ƹc����Ɗiڿ�F�pf4a
�1Qa�h�*傈hX3L�Hb}�=�X��,`� �v-�@�g;���������@�9�;���W:"+A�X:��`�Z0�c��8F��m�B@g�%g�hq�1Gq����P�-ֺ��K��Ώ��/;���
�}B6(������*e��i�^x��3���s�?%	;�7�۝0)�7Ӵԗ��o�N�yɺ۞s2�Į\1��"�+�M�/RX�*t4�"��wۈO*�Tm�E�	��c/�1'"p���1�ݜ���I��R�?�<��w�L1��mW,ҝ?�i�v�6E8��z����*x���:P��u���>L}�2.�����k8*c8m���^p};�ȶ)�b���B��&���^j	�㧒X�s���d�-���+�fȅޛa�U�1��X`����ǓG�C)��-�����F�>�<�]\�nش��#�$�E�fM��Ȑ�Ȧ]�u��;���8ۛP�J�&�٪�܁�,���;p��"Y�0e�{?N�τ�����u�V	ǜ�F	t��i�d�+��Wn�x��#X��:3O���>�t]q�_QxC�KPmUYHu��݋��C �ʗ��PT\������ycͰ��g�M&>Ȑte�XJg|F��%r�S0��1�	�Hl���;(�O| �}_=rLf���>���"@w��]����׫����Y�!o($��m<��K��`�=�W�زƲ��Dcca����N���z�"�`/s,�񩷫j��`1��k����s���}w�RJ�3bQ|_Q�N_�((B�*KI��Ҭ������~�u���̢>-��	U��I����z��iCJ�� ��&?A�<*�w͑��\�L��MϏ2kHw��R4Ms-4d�S(2D��:���6:rΕЫ��1�0s,���V�w]�qF��}ڕ��e����	d��<$�*"j���{��'nI�#@c������/#�(+y���J0�
w7�T�i�5����s�e�b�YP�ܤp�T���`%]�-W�}Hp
Ze����>�}50⛣��9a��b��CcE�)'�rޚ���%|���/�T�\�Z��jvڵ!L���������*��FA�����(("�?q=��+�����#�5��t��ι|=�K㎊�,
�I����M������]�"�:x����i�y���kw�*�j
�lg�=�z�������:��Z>'9f�y8Kg{�+�qF����]������s�<��\�E����"u�=�.�ևl�]�{�dj�����t��t�BB���*w�6���F����n0�Ԛ��f��G�/�u;�e^N����c�E��=N���F�@����<������얌u��k1E�7q��Q��4_�"mpv��
���5 �fTR�"�W�'a�}����Y�RG�������~��K���S>���d0������MP�z��Bb�"�H�z�B���<�Z%�Y��\��D�X��l
Ύ�8L�����=ԛ�ҙg��x�R0�
�)�Ns��B �@@Y��:y\�ٌ���Tpk���-��S�<�D1�<������ZR���U��oWΦ�l�|�;A��x��R��?��f�Ŧ]�H�J9'�V	Wշ�	�>=L�w0E1�aɅ���.�����?����r,Ď�Wj���!ջ,� ��S�B9G)�;��0��ዡ��&��#�,���8�=�Y�Muf/�;t�sV� ,[e�Z�����aT�l[yw���V��{Ё���_�Z���w����>�7y6���>*7�mN�cC4~��_�/T��ԕi(N���+����@̀�bl�K�0A"��h���K�g�2`e��5!�;.I��cyx-�}����$�Cz��Ps�	�|��bh�����͙���X_4����P�ٯ�,�d`bw<��o�D�r\:[s�-֔"�&�0�?��������6#��[-�慳
5���}��gI|�[7���C�������Ţ�"��Ar��O��`v�G�}�3���`ѳ�D���y��1��|�z1Gi�V�@8����������
2i�BZ�b�յ8��n,�`�T�l���ݣ��E��>'4 ((T�#�e�~�05�Ort{?�Zh�IH�CYq�	)P���k�'����&��������h↟b�)�c����ւ��ޘN�m�jH ��Y4Ě�Aap�i����X�jw�o�;�k$���ξ���p �hd�	o)N�nr>����R���C�k��}�>�|��PkuU��Sq�+�vH!�	(\��t�!j����_���ϵ�T٫&���K�}�X�����֒�Is
�1%�����`��JA�\ZtNQ��Պ��&�UȽF����- ѹ�v��|��{p2��4�q�,k��}ڿ�$`5���I��q�3���(MYۅ�v����$�`�z��ӹ��r屾�1��v8��R�$����r-���<�W_4?�"�=`k�E<���{��+�z��O��-�m��e�������D����dc?jH�v�U��C�p�*�C�G>��{���O���-5��hh��8�Z�l�~:B��ԓLc]�}n)<�.X�E�r4a~�p*s��t��K�r�	F?J��f����ㆉ��Xs Ĵ�/e����R�(2��c�.`0͢�G�7L��0���P"����>W�_n�i0�3r!��ө@��b�q5ԏ�?[�q�A�e$�e�ɴ6%���-5�Uh��ۘ���M&�/	�l}6s�-z�����&�^�J�؏����uS�C�K���k�?;p�#7�[�t[�5�٧���Nz�Y��������X��8�C��?����6�R������]�<zpa��\��R��H,���Y��:B
�PO��C�l���2\Sހ'G�E�w[�����[\�g�~pT̉^bu,��b6or�R�h �!h 
�6�`�5' ���4��B�K�M턕�Hx�`�ǗV���Ȭ�u����fp[��!�Y_"�l��iܚ�$�=�/��\�4=)�=�Bg4�k/9b��qB�r�Y�}�u�Z��l"��cg�#�xx�[|���uI%��Z�O^�j˓A�YB��K���~*&��������1p�[z`�\LP2\�L��u�,��8��Q9E2_B��j'Õ�6V�7f����<��Gs>9�R�؏�d���V�;���MI�m���pCP��\x".E��6&(j�B�F��wL͟$�����mH���u%����X�j	���m����� 7,~��� V����l��NS#���_�͖�j	�җNk-��߁������N"z�Xl�0�H:U�m#D�"J쮞=_D�>�4M,b1;a\�ݜ��Q�h��w�嫦�(���jݎ�!*x4��4��tu��`�W:���~
�Q3�K�VVd9:c�?�|ʱ�����Dr�֛��o{�T%����R�#7~B��< ���7����Y�f�م����]���0/����,�o��0.z�'}��t�:
h^�%�>}�j!����`M� ��ݣntR3�����_ˇ|G���
l�磍뙻��[Ɗ�4=V���?r֮��OQ�Ĳwc��h��=�$�M6��\��+�d���y�B����+ ��A3'A^D9_ҙ��U5��I�������l-�)o�dqfI{�����SC�d��
L��@�OC;����y�i)���.茡6���Kw�=��	�$��ո"��g��$XHH�~�G��O��"nBYOv ��yϮ�[Bt�JQ6v�-�S�1�	HRK�3<I�R�)�\	�oCd��| y�f �b������}18�V��sG�4^|�$t����x`hu���GS������~+�i���B�yܻ�Ӊo���Ab�3��#��"�o-H)���=m��i3A�H�:��o�L�\�I�nh�<5lstf���5DOڃ��5��Z��ӥ斢 8�����`m�P舭�I�g�|����D��u��kN�g�;e�Y��0ɑ:��ϸg^.��]��⚞���0�#�2�vZ������U��uR�����5w5@�"��4
"u�J����׻��}����p|�w�<4$m��#ln�H'���uQ'����=/����.�c��ǋ����?� �����la�$t*����7N��y�R3 �δ��(�k8-��#�:S#W�(���7���봂�i������D�\]G�7b�d�#�a$*TYG�ƛ�H�U�`2	Z���l޹l�9�B�e~6&�@e��y��:�5���<Q�9֡Y��!��1C�P���m$�8�8��Ɖ�*���Bы��c�<MnS�)3��w���W3@�K�:Qϸ�~j��E��-ǧ.'d^�~I��̂a@����p�Y�u!�T%"3q�����Y�G�����Z��.s�Gid��j�]���[�˦MU�j*��b����Cѓ�)��7#���p�����̟�e�O�����k���˴�����6�e;�#Ȍ�<����5�7|c��@�.Ճ�~��V�?˫M�RCtV�
w�@l�����v�n���I0�(]��D���}���x�G�hy=���O��!��d��+��+���6�a��1z  ������%��CNA�N�w:�s�-�$�d�#��0��RϤ�nQ�h'���e�U�>O�W��.��͍.����s����־�!Ö+�p�3���^��tJÞ�Kf�I�?�	�9 @�;iK;��9�z��mo>#�?7讕�̪17Kk��}NNF8�S�6�����G|+\���lQ�J^L[�3P@Q��{����U��z��s�]v��5t�-�Qc7��u����Q��}1-�: i :){���x��AXЂ"���V	�=��躺�PF��&a'K��q0�&�-RV����k�i��O����S�h���Q�b_,3E�T�kCr�E�V3�����R��UhD����s��_
�Ũ�r�,ADn���ܨ{�`E�)w�Hgq�7J<$yY�?�~I��Ѫ'`l��~5�OKc.�,?�-�Ӷ���'�>���I5�j0�J�����;�(�y�b�!��b�m��(@%mI,<��Qub�ӐB�ǽU����� ����~��,5�Qzv�]��A�u���P��Y�P<=X ���3E���I�5J���^�J���
�h�<�;����3���ГN�y�`�:����,�^��RUf!}h:�D���5�LU0����q�(���#�O�-�"<N-n&O�x��r��  �7�OU�Ӊx�G�l������)ek�=�f�0�
q\�ƶi�YK�1f�����jUM��1�j�2��������|(���T� ��������7|cY�߃�6>ɴz�
[�;?�Q�ۛ�N$�G�M�b�[��9`�Ry1,m��ZKބ�΀j���G�J�3h>��ެ���a���ۢ6�������}���6¾�y<g��g��V�'�k��v����������,�Zh�͊huW�-��'�J���$�a�n�4𦻞�t�݇����3�N�$�V�-���3IMO��Ή�+3J�Ľ,���埳
��π68
W&';�8��W��e�Ý_�N�6H.�..DvX�K���=󫗹�8��*�@��Qé���#�M�J��2|{�r��,J|������.�����}-�#���=��$�u�m��X6 ������ b�t�1� :�N�m-b���f-ߪ����e�}#Ht������c�2 ��~�ETz<F�R�������B
l��%IDl���)&��P�[/�[M1�
�ۋr�ԑ���н�L)�C9P,<yM���?�v�k֋����jj:C�!8x�݁��B$�!�l#+0�c�:���ꗟ�7�@"����M�K䣹PJ'tm�j�9��e�A��)�w$�nߊS?��.��G][+	�}^���m9����oW�x.�|?{Eh�[_��}z���5�8���n>b�l�����r�#�O#�J�-��-�|jo�n
e(�FM�549���N5�j'�Y.��%$��R$��'�9��ꀥ�O�=sR����2��|�SIoz"��V�΃�2q���D����\=|�N����45�q.4Ű?/ܤN�&�>��|�i��M��W��b�-C�yyn2�y��2Ǚ'Dn֢g���
ub��OB�I9p�<�H��/M�I���)ǖѪ�ED��>y)�|�Ɖm3a�p4�ܺL��G�-�w'�jZp�^�մBj�V檭R��*��zÔ�]��=�q��������y�.�jMI!$�7����*�j(]d�]�O㊭�9�U��\ڋ����3��%�񄍴#z<J�{��}n]>Q,�wYsm���ۏ�#�^Ğ�`�0�Z�t�6���A!���#B�=�"�}ǒ�w�x�G��i���z�"U�#,���J�i�**Tۮ7�tL�$�D0"�%	FZ-R�K�{؆��ޟ�?���lO��~%-�D!�;�C���Şf��Ѣ��8
,���Ż��!���M�&�{�j=�O}�4��{�md�Qg�O�	���z�V�v�_��>w_3����D���O6_#�M�qm��zGv`�x�+x~�J�Ѩ�fW����`C��%\�{:Z|� ����J��Q��li����ĉ�w��0�� g
�WC<�-�a+��>z��Sd=���~ӧI���,��8��-VP��t�_�!>�>�ם-#>��R4�9fv�[Jf��<d�M�#��Q�X~����z-������B�/>&n&.�J�-c��/z�s��tT�#
�i��0�\���S���ˋj2�[��Cr�ٻ���X7��uy�lb�,KJ���A������G����<�K⿟c���V�b�FO�a�q��\	�I�;�HӍJ����G�tq�*��4Ơ���9��h��-����b����ބ���6��A�hMf��C?/�3��m�nҭdꌌn��N<)!��0Lы��������ﶔ�k��rGH���:�!�z�v���S>_�+�1����g���-ԑ�-ۜ&�ukGM���x�2�Ӑ���!\�}:D����%,� �r6����v�A�}?�n��ܩ��{�T|^b�O�6,��f�Y5���t�8�����'��V��T�Te)N0��*}<}5t�3�x=e�3�@\�[���C��'�<�|���*\7
��yS:RӋa�ةDb��\FV�^����S��N¬y[���#�*����%h�������w�f���}ż��R���8�_m���[�\3�q�~1v�[�.��U�!p5$��e>��7�r�{��'d}�	�ϭ� ��,�1�_ڔ_R�Q[��	H�t	��O� ������0�т�+K*-�A� �]+��WBc���p�oa��lf{��A�}�WXH�n��u�
�<��"��C��Y�d�h�q�\�[��q��RT��@N��<�{��*�.�|`��\����єҪ�"Q&8nZ �.ə��[5��'���������7�_4M��h9	х��S��Co涴<��d��~��?��y�mNmKh�|O��OU�mP�x;�:L�Gl��c�B�����
���B���y��J����� ���t7���E�?�0�>�Sp�oK*r͹��;4�
�����˽,c��[z���u�ˬ���/�JCbd]�����P��N���VW�ć�<M.9q�!ͱ�D�N�F'˂��qv�ց8v�Npdژq�X��l�D�+]@2S��7�����y#ܥ.�8�0��vC�i4���1&���ݛ��X��f��Rt��m�J	Ȭ%�&�D�:^BB� J�G�i䠿��S\Q�PGz�^�JA�p�=�R��:}co�o�
4pÂ��n�+�1gi����B����(0S�.�?m�AM�=��k!�=�t�Yʣ�6R�Ս�Uv�A!���ӧ�ۇ�{�Mv�����	jI�������FѸ:ۓ-�6F�g�]m�I��m���fz���������������U�J��U����QF�Z�T�{K:@8"cM���?�+�&1�hXD�>5�yE�?p �=� ��S�����gq�|wN��h4�m�H���A��p���b�LԉJ��c��`y��cD_���L��MKZ^�8��⩆8���n��W	�BOr���h)�]3{�|��M�����B�?�E��>Ad�v�&[B�1�d� a��@h�E"\'�mfƟ�J9l�_�0���3�>���s�; .K���!NTI�V~�C�Oi͆oL ��8��r`��'�O�e�����+y���v��ko�n'��@UV���$�x(s1	��2f!SX�N� �E�G�O���� ݆ʘ�g&���\�#����`1��b�	�^��T%ш*�mV�މ��� ժ,BA�����o�PZ�H�z��?J���c�Yt�]�5Ӄ�:�n�'�fMV�o�(�G_�dvzQ`���εγ�/v�b�&�m�DPT��b��ظ����Q��qp��
��!4p��L�������t��9�n��-Q^��@���P�1����v)��Pw�#TD�J��UОb��~�Q��R���M@4bjз
ۓ*���-�����E�̳t�h�D2�g��^Z<3�#Z��ȕO��n#�q�i�c�>ļ��0���d�f�,+r�p=T��Q-�`	���kA$/���&�	56f�+��q�Ba`���H�W&h.���m�i�֐PzEh�p��A��~\���k):;�"X���b�7&�a*�)�+����O҉������rM��������I��=5Ձ���������E
WVδƼ�����{V|H�Fܞ�RC�i��ӿ�^f7�r?���q����B��aM�NY���e�=	h�T�R\�Q��[��]��㒤iK/U�k�7�G�'�4�__�C�����A�3�>���kY��A���q�4.�US��㹿2pt&z��W�8�|'�{��:�9U2���ՙ��ܔ߮�{�O�7�݆S������VKJ�>`}�V���Z�c�%R5�X�'u��M���,�Aď+jJ�M�%q�=�������J�-��d��M�)D�	�����6�?}ˇ�@ Z\�+Hګ�� Ja�p�nF��Y�@�c��<��VtQHu����(�,��uv��4jb~HKlB�
��s񆬉�������2Z�/��QI���uM�Ǡ���T������W��6�O=ַ ���#`�q�-2_{��ԇ*Ɋ�G�|����Cu�#�Tr�ӓ�ti�����h�-ش��S��zO�/A6E	�ٶI�:-�11+����-�����A/�fO��7��JC8��[���W�sA�^�5�^q�r���"�*�`��}:
E@��Z�	����g7��S���FS �=y}�ͼ#��2��;�0��H��Y�B�v���MQ@�����^`**�r<OX�"���\��o���ͺF�����$$���ؘ���k�	s���x�5VvJp�D�N����qd�ާ�)G��5;h��/�$���y�X_���r�t�YA�_�=�ν�r�_�)�%W����͐S �Y��8��T�8�r���f.����"�u6�Ȫ7��g��P?�J*�RX�c��8�Ida�ɐttb:�X��{`�5ņ4�7$�S��p��-�*�H R_�W(%-����R
��<gO�}[�I]m��u��I�ų7";��Y+z,�9��#�>A:�
��U,�.�H��7T���j�?��Hjy�}��ߣ��=�m�*+s��B4�����|����+T�yC-�b��X���E�	j������i5�cSIӵl-)��y6YU�6��k��\�0h��ʜ"^��x}��I��8U��A&�AFK����v� �HS�A�Umw���;��x᧠�6"�����^|��Ye+E3_�����������ƅ3���]�i���!|]��_?�
G7%�8{K5�Z��o�@�� �8��a�g���"��Z����pW �s}l���B��D�j��[ؚ�4t���Q��oNE6:�/��� �Y�{�Z4Y���_>��h5���Eb!��+sIF�3��-����V����*��#�:�7󏿎Ӈ�ܦd��W#�B����Z9��[ ��ڧ�	��A}1U�ا�m�;-П�i���5��i����|"��H�������G�.7��r�7���j�v�����*��iO�Egv��v8�3�L�Ϋ�:�~�_�!a�ǯ,�)��o�E�Z��� �9�'������X^��
�y��e���1�T��_`�{Y� u�i[\�N�eE���Q� [}D2��W~Dh3m���SR2��U?��Ⱥ�3���&YV�uQR<�Yo欝��ٗ�z�����<L.��W�#�*V=M ���j1Y�$�dI���?�l�vJtL6�~���}������ى�~n`Ot.�#���6&Z���W}TWOa��=K���~�,:��)}���d��QeoE�ԏ�1���'hu����k��A���
���S`@,�a~��@snI҄�:��ku0� 5��F(?�P�X�.���Qu�Oj7�P�6P�ih�L5��i��.L
#�n,�]����w.V<1�#�����:ݐ�-9����}<}q��&�%�e]>�趡ۧ���*m��C��z�c�1�y��G�݋���ָ�O�����Lz�t�� d���88�����'�n��Wq�z��p�EB�K#x��Κ/)�����i��NجCU�	�Vws{�qhdDL��|jAӽ��e �ł9
�[���m	=�Y?����O<J�~t��c�-M�.+5��:G��l�|tд���ɀT�!����پk6,L�|�Y;�����.�c�m#@#T�-�PGd��=�X���e$�Wxa+i�z2�6��)�2(�Ug�&
h��j�;i��6��+�z��kf���+�����H&u��H��I=0�/�h� ��{�4���c��Ȯ�N�7)�ˍm�t9qVfAbR[z�����Y��t�h���uho��G3k�U����f7�-�4C;��O��b$Fv����^�m�\#R�I�>���p�E�Вʣ� D�B�$���糃�{��U��}<QHW%�ÿ`1� a�0 Tw�h�U��'���M�TS�����oܶ�[��?�z�P�z��U>��;mS�Dl�8�l5J8�='�������/�k�+�����^�����jI�8�N3;	W\��:0A��/��|�%��՚@�S�^�����I��z=��ֲ-���b�֯+�x���@x��aeH�g�|�s��p�9�-_��%��ٯdE�oU�$���y��I׀�a�l-�6�Pf���th�Bn�t�L#�e^�DM���1��_�! �|G�O�,9-��2�59ʰW��e0�r��YY�5HG��^����^��!V��o���#,��J�RH���s.y����۳��0W�4�i��,����}���aJY�_���S���걏=�4��og֖��%�p��({��QXuH�D��S�*�P�(���E�rk̋�
 �T��+ �AWz�@�1b�?�Ǣ�W��8������玛q���4��u��?x���q��'�<v��LrQ�!�(H�����k[��1�j,�V�dS��ə亷~.E�q~�A��J���&�<����������JN3�
+��7�6n�r�]���$G~ڮ�c=89�)���
=ư/l�4���
��4u�x��Y��
\F�L�h�������fpTK��&m-���B-�O��Ј�
�n��)�:�2�ikضd������|m:��dY�K�f�m����:�m�-�LB��۽���p�<��w��Q)��^�SXeQ��0|t��4ׇ�\�0Lg���2��s��z~��IKx�����F3C�9���uӟ�ɚ��0:B12W��� z:�u�J�a� v-����Q8�(Xd4nB��x.u�?t+��j�3݃s@_s@S`�|r�Ԩ���� ���f&��ך�8H�l������d�ێ�<�̪d�8\
���J�5F�=��9��Cd٠��Z|���XX۪��7v���I�U� ��q�Ì|�8<q~���4�/����� &�����b�]��+>�8��i?S&�B��خ	J-k��wƖqc���8,P�g��Hؖ��u�!愻�y�&��m('eL�,�^`����xP�l�41�Np}�uh�C1B�5�FeP��F��]���]�~��6�.�J�t��� �����ӮL}��M*�� �?Ic�Q�=|�.{ 5��g)�L���pdd��ڶ@���&z%i��oo��w���@g8;9�u��f5������>�Z�o�O'�;��G㵵����1��7���1�y�@�.����M���x�Ǹ^�Q)8��U���bA?x�t�օo(Ά�$i��yIUC��t!iӪ��Q��F���i���u������ߜ�:�֗�,#L����a�F���H��C�dT�cL���v$��t�:��
aF�����O�n��Jxr�I}��ȿ �CNŮօ�}]�=S�Ե�a^Q�x{QWGt�H>�3��d�����;s6�ˬ��Y��K��J�7w%H���Z��L/+�%����{�
'u�a��v�o����yhA%�"<���:�O�f%�^u���A=x	-�	��Z��ŷ�Ph�t���s�[M������ n�5-�&�R��8^uq��VH��O
I��#C"5��%QR	����ˬAc����w���>~���6�ЕWD^�m��{t��H
f�9��U��Le�0�H��+���꩓(`���}P�W8li�ٌ��~Շ�R5�|�>n͚�ʥ���B|U�����w���H7]��uM'D!��`r��>����Y�ӷP֟ݲxy�Q��y�$�H���*	��?�ʟ\�u]�&��/�].�nE#O:�|�b��#�����7H�?.��$��P���uC]M�é���X�����Ay�]����4Q��f�<\VAhZaBX��G��r�����<_��Ty'�qV�5�x���1��PP��w��s�	�$���>y"���[����]��p���)��&���?F����$�c�Bn��,E�m9��;#\APe]�F�ʊf>���|�VBw.Ǘb���Ub�xTT��Ëu-�J�������㺂n����n�y�Xx���zO�M���1C�oJ��],�u$z_ٕU�j�mmw>��k>Ww@G+�0H�� ����~&Ii^�X��:� oE�Ȣ��%�n~uR(㏹j�*�r�Z��'J�k����U��~�ڞ
�T��v�Id?�1��n{QBߧ�6я�+�� ���a���P�v�(G ����Ԑ�� �q��eF���g��e����M�pet!Mb��AF��(�U���W��^�TN1��I2����<U6�a^�^UK�3׽�_�Q7�Nz��������c���&o�������r�"����Y����4�D�c*�s�TزV�%�{+�6{?�U�f��zd�]�g�ó	�l��j(Lb���$�G�# ��S���I[�j�M~�pR�]������[�
�YA�k �R)m��|u���~n//ڇṙ���^�:�W��X���4ٵk���޲m�n�Z�JQ��+g�]�B��-:��Ϳ�=�K�ܿ�
H0@Z:0 ���Iv��}<�@�]�2�b��*��\�vp�5w���$��v�E�x��݈�mA�O�^�T&׎b�TA�����k�Z�i�Kb������EGp��ɢ������(�^�X^݄�l> �yl����I�bf����g��o/m�Y ��4���Q��t�A�{;I��2�#����6�����Id)�ZU��h	P�6�c����(�bш�W�~c��-�=����Q���؎�d^#�M^X%%���,^�>�Pgl������`M	��Lb +f⍀M==Q̺,�����: �ȓ?��\���~9�F�w?N�тu5���Xʏj[u���"5H�i��gUJ��Y:�E0��/xj�|��l!�.;#]�E8"d(�Yf��	���Gf��1���b=0g���6��.rW�؝g@�F�zm��_ݤ*Y�e��+!oW�94�����(����+g"�ڀo������>"i�!SS�u�S��E��3�0��x�5���p��5]����(ށ�)Wו<s��H�e���!��]l���F�r�+ ��K�x�QM�9%��V��Ȍ�EG��X�.�C`�%<��w^a���[0Ck��r����0K�jxg�M9Ghy2��m�
���v���ag_�+�����_���.�4����������u�?�(س�C�	>����E[6���:L�����q���g�L1e�ʔG,G��-��)<��Ǽ_��\�]٪f:�(�q��w˚�8��vʅ���(��T2��8�0����pw��jb�B�����v<d�Q�U�2*>��5�ٴ��K���H��0O��[<�P����)��¯	gG� U��V]�]�Ld���x�#,���-p��Gw�[�'s�߭c�,
�JS�}��L���ϥ���I�5����>:�Ӷ�v�փ��1Kr�h�
>#<��F��"�w���?3C�`��T
�iGh��?�F�_��N�/�c��ւ�a|��H�.��)on#z�F	������[M9�^h��g�/����}\�'�8�z�7m�
�ft.u�\�1ɾؗO,0�ϘM|�lL3ہ:1���zrq��b�����E��؈1�j����i1�ཫ���Fb��$,lۗ*Y�*����U�g9�ǔ1������W������ ��:�i�����4c{�H���9�є��̪@F��~����N��cY�b��5��S���t��1�?��OiSuς���u`8{���&�:�n�G*�����ៈ���{�{��2���5	�Z��K|v���b�]p��������<���gK���U	��mg�<�L��H��FGcFf�'cՁK"6Z,��u�DM������z�֦!�����Ք�N�
O��*���T�vO�$7��#�#�EC�j8Ts�s$�K�-|��ǉvW*���I���5�d��r�7���a����ٷU'S� 5 ���^@}�SI^�C�Q���A�-r;�3KD厰�
��5!>����*�6�t���S�UEC���7��J~�n�}/�VS?�(
r���Jt�y�-	�+9�d�LxІc�DBO���M��>������{[��Q.w�3]b((�`����h:xǠ����P*h�mg	�]��U~����f��������z6������yW_| GUl�Qtk���u^z�#�l��D҃��F�y�[���@D�SˠO�����KJM���C�1�
�B�?��d���](_�߾4�O�4�"jÞ`�=�ˑ�L�g,�����!U|}���4s/�����9tuJ��h�/�XhU>��*0�@~-&��&�m�&�G4s;<�|�%�_I8��[���~��M�;tv�A��eL�|ϳ�Af$�u�����u�X��1P�9vs3ӈTo|:'�]i�y���@\X�%���b>>&=�T��ǣg��l1���Zm
�9�9���������CTr>����/t��$�\���]qy
�]c4?��U5�P�������4��˙�aЫ�SK"�Z@��b~(M�7Y��1�S@�s/���&��dO��|�s�d^��z�[�����M���d�l|R��<������R�rߎg��q��'#�3��C�*�J�k�իv"P������7�e]��O�����s�>,�Ѻ	�dT�h׉ٰF���ҎA�* �����[�J�+~(\�p��� 27��#�ܽ��.�`�ަ�;4�'��#`k�� �g�ݎa��CdՌ�mo�olc�I�-`Jnd�Uǜ4�W�;���D&\��+�\$��J�#�4��B&8q�,��O�f�&�Wޡ�U�"W-4�^�<��o���� �6i����X{�	��Ҿ�cr�<��=��ٙ���z<�p���&���.��w�rqi_�:^+�o�*���/���N��t�<��?��k�x�π����;pk\�P���_7<OFdLj�e�6+��9$`T���I�{6��U�)��Ӽ��_�?iE�Q}��B�N/
�9D�9_��gu΀e��t�Q3w�x�7�?�G5s +��2���Ns���F���\�A����k�ȝÇ�?�s�%H����`��w����$��/�Jd8���b.4�� L��,��e�&���1,&�>���x��1�9g��wi�|���uE8�ь?d�h���H�)r��-��$�%�kC�۳]�v}w5�~d �j)�����Zp/�o��e���j���eA"�-$���*"��$�0̈́XDS_�3����=���`���gˠ��-4dH!�6�e�k�C3*'1=G��*��;�A��SrR:�����e2c��aҧ2\Ә��-Wh��o�z.�'j�%��-���_�gt��9��60������륏�v�x��ߡ���9[Ҍ�������g%���{�0!��4Z��X�@��rz&�HC���G�R|��1����+v[��)�8~�P�4�^	��JR���.�hN��v2M[~�,$氂|�ow������cQH�I:���R�Q��l|�=����I���`�Qk_� gM���Ss8+DVA�ߊL8l�X�W� �kBj��^!�(/Ut�G��I����2������"j�d��c P�5_�\��#?��i)6P�	�R��~bX7��A���LZas�-ڳ�T�? �v�*���Tוu�a�)G�� �d�^:�L��.R��o
V�X����S�9srT�����)XmmnɐB�o:m�[ݷ뼒�\��ท�G��v�_���k�Lyα�_������!�ꁞ$M�}f�����J�pSn6p�j/kdwS ��j�N.�ǯ�-M۞#����
7N��	z�� ��W#wXX�O)1U[V��V��y��$�4~��)gճm�
#2�Qf����Z�e�t�BUK_�d�8v[�F+vp�����Ԣ��i��!�ע��;(�K��C5�d����S��q�/�؉ �{nT�礨�y]Cf4��3p�e��Q{Ģ'�s�⼽���jA*�#G�Qb ��Y��I�,��D<�Z�t��r��B���ܓ�p7-�K� M3$g�Ýզ'�����p�@�~��>)��6@�����P�͒�iUH���3��Oj<)���J3g�o)��%d�P�J� .O��8^:��N7M5A�:g�p�$qQl�<��OF�*Ձ�1r1q�}­��T�Q�D����l�:��l�L$��{c�lW]bު���OP�üf��M����p�p\ݒO�`I����Eڡ4(��6б����Ǆ`%�^��j-��N�u�����cY� ��LE�-Wӻ���dq�4�K�Rg֢��}�H���l�ȿt,;�F*d�ha$8��Ub9)#�[F�>���;P~&�{{�"\�v�N�����V$B�>�ڪA'(�N���D*+�E��M��Z���踟0��h�NZP��ў8��̃�/'�F4�G�
���vl��)}>�Ѝδ���90�	����z( 죧(;%�������ۡ��P�bt�?͌��*��UK%u���4�(��CR|,E �]��bS���E��(0	���\&��'���s����~QF��/��0�f=e��!�#�<�s�1��!fx�e~TQ��R����9�������äT���&г��J��2j'�z䣘�� �a0�|�:��JS9�;\'j~G0���*���W����w�~��JVR�щ'�?� 7���RV���L��Z���d��}]��ӉX_?��SI -"8� ���%T3�\'����.c��.O�@���-��Gw΅�ECo����+���O���H�����i�\x3����/�dM?�ZR���=�~f�L��P�	웂�V"\�(J��l�;�g�������`��c!b�|�9��Ѿ�G��KF?�
�ဇ�q�`}�dc�P%t`��>���r������+� �7b��XE?���{fNO�Jh,W�Bח8�{�o݈��9��V&v'uzU����&�{��q��2��ߑ�����%N�,��s��~��;/i�2dx�ڳ���R��!��<�Q��u��x���ksZL/�ʖzI䤂&��4� �U1�K���Z��"�|\%Z����V	x%mi�!dC�h��.�"�e�Z��,�&�b��0j4}�Z��S����'�Uɐ�&k�I�ٙc�<�o�[\'��6�G�]^����?z= }���rJ�Ʈj���1��㈆��vJ<�n)������$%O�t���B�zQ_<�Y��wr
ҹ�،?fr.�!Pn���Q�2P�b)��$�����k_~b���^TW��{�n�7��������:��������e�"E5�WWqħ��̲h4?�,�����w|�9~d�E��G���P4�	�(�9�Uc(�M
?�܌��}(T�o�H�-���=�7s�尴[�SH�N��q& ���K'�'���C�r\&bE��N7�Y��
�Uy����/�?O���֮Ө��wu�KG�C���7a.�J��8~o��#��H\{E竣���:����:�taʛl3R�%}I��XxN�h���vxZ�|�9���{��_�$��o�y������(	=�IV�;�n��)D?D�(�ܞS,�%?u�=$�$N\��b~/�!�6�0�4��u��vj.��p����=�M�*��ݞ��ܐ )kN˨�"$l���1DݹJ�@����cB�>-}��6�dU��|!�%������*������ʎ_��,�(5RK���n�}���Cǐb�e�(k��� a����H����nu�4x�P����ն�~�l0/�jH��^�Vc\�E?�wf�:��_�F1k~�� gP����E�ܡ�Cnet���W)�Mq�
X�*D��tZ<f%&^2�p���X���}b�R��N3V쩁{~��Pfz�~]vրm�_�J��(+0B7,+V��_7�i�N���EV�Lޔ��J��|��f�q��J�S�aIc�A~�g���s���Q~�ʗ�r露qW�-%[�����-����P�ώ/����r=�͌�����=[�u�t���7G�R�5���qf�h�,��*�<���\�a�O̝`�g���}�4�; ��E@�M��(��Dݧ����G��=��䓘�SF��cb�����l�F�T������pˣ�[6�����k�0/������-�/��a�S�|�.b����}��\*� �M�w��ǃn���t����5�O1|7�K���r4㚃��>u���o�9�Ys��s�������Q�?���t6?I\��4k*i��P.���X��`�l�1#��0[�β��2�=�(��@����˨Xs� �y�Md���ɱ�K�^-�(<KԽ����(���>�)�1ǉ�����+|�$�ڗ�<�%��{�wP^���!���R�!2��X��2�ex��(�tb�K����O3�v���%S=|���RY���֝e�]\:�犥y�N	ւ�\e=� ,���WJ0����B6K�C���ob�9�^~����‸�4#�F=�n@������s\`��?oݾ���o�v��� �%AS�cP/�2'�Ő^ ;ҥ��a�HmB`�鬄�����'�����԰9�@M2t�{8w���T���<!_`D�;����~tr��
1���~�-�OZ:6��@s�ׅ_�-�l�����/���'�%E�[����-%pJq�͸�!�A��b��%��
�(B�gr�n{he��^��U|w���R`F�1lrP�������Q�KW�F^��h��.����ܡ��®LD�6�G"��!���w0Zl�|��^{��^N_���c�z�zr��L�[.u�}t��q���qު��.�آa������X��K�*1x)��c�G�<-��2@�.B�a ݍ��M,Vk���jd�k<��,J_J��'�:�2L��,Px'z��os|�cܜw^ҁ��"y����������?0j�.���^�7n���=�|W(�I�٪=��8�6LZ�}ݑ�#'&ˎ�a��T�o�5i�_e˛�.s��Q��>)9{�T��!$lFr��a]n�����Փ�ݝ>��cL缷}^E���Z����F`��4��e�s[I�;���r�yӅ`�`���b�i�C�d����qW�3@�5�z�]ga3��)A:��ƪ,Gj�Ȗ�&��]�U�Dfi#��G=pK�������r�w؏4�tz�{�h���M(������噶��U�,���R1���1�m�ʪ5f�,<�E����U��ָB��/�Ҳ�]���U�.��Q�1΁�1�����Y ��^
􁴐4�9��A=�`������(�YF����UG��	����RK�� �[�cJ�V']W@�FV���!�U�Wn6mg���2i����#S���3aH)L�UM��G�sN���3��,Dsr�ȵ�Wp`���3��{�AS�W��h��}�U3X�0�>p`V�P�@Kg�H���N��'�w�Ѭ<"M�T*�BBȢ�;��r�o ��U��$=�?��m�\?�+�ط�.�U6)m��C����Ų�8�j������xq���<�3s�_Q��@M�jT�
y;i��M'�tN(�r���|�{�]<Cbq�$�eZy,�c�|���`C�B�>U���)��w��c��R�^V��yM�0�>�5I�5+���(�����t�=��I��_�X*��/HEJNjn^]̟0!<��͙,�� �b���s��"�����%�,�e�7�$*o�P�Z��_�wFg8��5oIݟF���,knt��t���\��$>���HM�-��e�V�a�=,4͛+<����B6�@�En�Җ%L/`ܕ8 f}=m�{hf2ڧ�zua��� ���_��4�R�����&%H@�m���> ,B��	�4��V�`a��Y�3e'�Y����嶧�eZٴ� JM�35�g1G��>ZHP���4{��i;��$��I*��
���j���QF�8�?ȓU�)�(����@�]������X]t,I�J��<SO~��j)�ł��f�PatW8�u�@��x�'��<�R�]�G�N{+��Q�p�x~�n����#+Ѳ���
X�O�4�e<ٻ'3�-,�R��-�_iw�0��݄?o�L��Py=�(���x��Z��}6�&]�w�%1���0$�x|�����4�����J�Nu_���w��Ej��Cj��y��}#��u���<L@����#�G<�ʮ)�k��#�{L4�T��(�8!/H͢��+����;u^���))�he�n�*���b�[�辧�e���@J�.��c�=+��
�%\�L����7�ɂ}�W3��L���L����� �-�m�7�w�Z˖L���y�1o�u.!�R%���fQ�B�f�	���c h�[AT������)L	��{gt��8c�*2SBlC�bX+�Q~B@�ʇ�N�?X6b���?'@ห �j���1ݐ�o��ܽ��B���*Ƶa|3V�v�po�*NXZ�|]����_�ޠ����6���q��݃*Z�hRᶏ����x<�1R�t�\t������0Z���6� hZ���˞�������
��OeV� #*^��G��q˄:��O��yr���cr�y�Z�o@A���|8$��*t_/L�٪_�$I�����]f�����J��v�����A��Y��x8�z�
_aB��"��Dz|�, �@�3ܳ��E�f�%ι�[��.���'��[�v�,	��׽r��2��c�ѻ�q�J��W|�9�'���w.�C���$n_ ���f��̚6�0��]x�n:fJ�����ϣ�i.��臂� ���`�P3�Xc���8�}�7g��V��ނ��S�c_Vw�Y��:�='���?�b���. G`�OY*x��n۔��@�:.�Ɠ�ސ2���x;&�6<���R�:���Bq;)h-{�9V�V�.�"��s�]��"�s�H�(���|uF����1ՠX,��X�g��iQ��[���ko��p��6��G�a�4��b�g��������7�Y#;�E}�_.�g2�����)y�8!.ݿ�u���U��4+aS�������=�n��. Gε��Q�k����@���>jE4ci57ɀ��}R7C�_��ծ-t��c������ϹI�V��)�H���pnv�R�����������Dt��T���ƎCT8G!x0Y�7���Єj"o>���+M`oS��r`��1��h���1�#R{.J��u��/n��s9�毋�A����%���Df4��ꄀ׌]D�7��J�r)@���
E����j帇��"�7)��Q����Tn%a�ٚ��HT�ر�d!���6����e�F��b���@@�jv�#1�~98jm�F�3������)j�[6E3HP\�gG���j��+78^c�f�8�4.ʑc�fE�ҿ3���0�+���S�k����1��D=%SS�96���O�9����U��h� H9(���K�x��cD�3l�@�y�_9��A"=yv�vr��jS@m�@ijR[:=g�=���X �>0��Z%U+�	��,�Ν�|�^�|Pp�I��D\@��������V�����T+h�⟤�����P��g5��k�~��z��9��Rt,�O�$7�%�a���,ߣ���+f��Wf��4�^އp��pSB�5_	yƞt{h ��~���ƀl
��f���3��I���":�j�{���"�m{���IZ�2���O�r�KP�e��V�~��]�gC��A{�Q�b�AT�B���꣒�jA��t���[���,�0h�oܞ1��r��a�}�Xx��ڱ���DL߻�g�����l��������0�P��ZY9�˝�:�λ��x�݈|W��j�7��K�uhފ�m�o�	�CSlo�CE˼�t��~���>f�=�΂g7���$�<;x�<�~��{��9y�WP-c��e�~{P�1���v���D
ȇy�G��*94#J	��}t�k�=I$ܛ�FQ��#����^~0n��V�E����^�7Q��-q�
x�����[6K����ެT��iq��X�1`�[�VQ�������;n�q/%A�.R��n%, �ɣ�,�N��jp���z�]yk������wt�~+�!��>^;�*�����3/�'�����ޖ������(�Xh���XV��1����Y��^�Z��SB���Π*�u,�P�RhА�MTg����\�����������ӗ^"����m�9�?�.��-��X"����	����`�t)��m��L�� �=: ���8S*x��tp��G�-�}��E�G�}��b�xKکE՞)~ ��O$�}����2���-���~���T�	������������]+�фI����?�rmdyk�L�/�riش:韼�,�8v�ز٠�P���W�;VSk؛I#��6vLJ�nq���>�[�_��b�Z�S��N
���0��p��7J0C�#�#�d��+WLE����!Ǉ;ryW��"?!V;��!�j?zO=�I�4��������ڡV-J f�Z�6�]@D�-�'���j\�B�Ud��q�ΣDz���Bp`c�^����v�W�-n"�������Kט2��Z&$`�Gc+�;�N���	����&�%TEa��)U�����O�R�4i�� v ��h�HQ��f"<�/�t�#�oœ�|��β�[��юBYm�3�$���\��� �!�pR�����j9Ss-3���ں5��S�7���n)�ڈ�ǖ���?{k
Ҁ����k;��Bc��Нh��[@s!�/�p���2F�Ik|qL��@��о���;!#	Rs�c%�!zE{�����ax��&�lM���Sd�YYd�7_��^֟|q����G)jF�qZ3Y��h򛑉R�Bc�vxgb4��W$����7s��a�ѩK�Vϱe����f
c+����"JYFz]@)5�a�h��LD�9�>T?��qm<aZ��0�u٨���+qt<<��O[�]&W;�A���?�$>�$�:�i�g�6�ꑛ�\�|��7��/�c�V�o��RF\*�y�T�����b	b���M7���b-�i�Qw��AO��v2	c�%�.�zX.iWn�.�y�H�k�~�g1�T|V�/σ��6�7Ӽ�k���#GV�@K�@�IM!�)���~U�m,6n�}��"��Q%t7���m��U��G|���yxx���)g;E��WS�j��w_s�����j�47g�/�B�{R�)�nV��p�t�R�@n/�� Y�ܳ�/Y[x@��7�X�,SMt��:��ޓJ��Ԡj�����FSXH/� azR�߉���}(A�VQ�m�S̫���]_s (�D� }.&rQ��I��-l-v�=$���d&l���>��Mm9�.��;j?�\��d��'�4r.cCF�k�=����z����!s����_}�U�;�<�B��Ґr�ޓS����(O8^C[���R'�2Ɯ���`c��*��J��	u�X�~��LF=��P�4}�|N���΀��1�q�.�ׄ��	�?��Z)CA5	SJ��Ϧ�<�r�*a���jD��éL�_i���b�h��WN��'�t+L�e�׬�)����*͈Y�a���)BHb�v(���,#�:�ρ����l"������.c���ɷ����ft%	�A١ui_W�?q�Ȍ�b����͟������fz8�1T@S=$�Oo`�����8;	vmd����+�����!�F���И�k���׏��T�Y)���nQ��i�E�~��l����fS�&<��8�O�����)[�7�X�N���>d�Ɗ����QB�z�����}Ʌ��(�� u�#Мio����|M���l`}�[`T��dTUK�m�Y��FckѤ�P�b�[�A�G��3/��+�^'�7$%��.���\��VOwV�"k��;r��>��qX��ug��_a<^̮ϗ������{n�Z�OH��Ip-p0�������jg���3#��^P��TsZ���!k��3�=�r�t��;���dP���-:8�b���F��푆�[�<H.��LuA��,?|��źڛ/\���������P��A�QjsI��dz�qmޑ>�3�ټؖ}�e��(YN����Y��p.�-�Eg%XV���`��� �dCP�qވ8��y�2APm�,ez����~_������I~��b�-�������	&�yBm�C�3��e�/���5cݏYR<�[��% =��p*0Ao���A.�+/a"~7��b}���\, C�D���9�uWgtl��&�����,D��P����E$���m�����&�卡��[�ʷ�|�A�����g�B|�M�Y5p>��o�8�M�9���Ħ�Q��6�Y�ZbW���0D��q9.��_��	O���j��mt�L:(S�2���6���*<��)����/��_�9V /ު��;q�ghy�2C����;�a��[ue��h_�� �O��9�����g��~ˇc
�h��B���n҄D�C���^'�'Wj�C��C��!�
%&�� ��-F��z�U�UTGI�Gd�υ�u p���SϭxJF�%��7G�	ׄU���Ey�i��>��y����a�U ^�bW�NJ��B��ĉ�4�����s-�\ў	Ʃ�{�&+q�⪋��1�הiokJ qN�FVٗ��<�[�]���7^�AH(�E�	*%� #0��RX��IM�z��Կ�6;�&����%�#e�9�Sn��'�:%��Kt<�̀}�y���ɿu�*�	<	"����>UUJ8+lѺkH)�|��ń�Dzb�.�c�O5]�#����Բ���a�/-�)t���.>>�3|���5'祮NZ�C!�p�,:��R����Y�2�����z�#X	�\����ezcq�'}β���>t����Q�D�-�-��a0ޢ�z`��s]��{-�f����	�VXa(K)v@��e�� ��P7�՜�x\�Y���T�3׷=u���oJ�� �fj����2:)�S��T���6k��3�X��t�f���pr� +�A.9���c3A�Y���WI����~D=��ba��y�4��Z�#3�3���p���K�I����f��bx��Gg��%����Q.uѥ��Q�����Β����*���,6��}x��7ȫ��Z$D�Cx�*��^Q�ln�d��A���� @�l����s4�-qBRh�`���;��
�>Ʌt���}kH�t�V��dPj+ҍ����agr��xk`����v!Ƒ��Z9�Ul��S6�T.�^G�����U��H_}~��6�%mW�-����hړHQ}�d�x��
��@qAj̋�QM�	/����� �zw�|G*>���x����-b~��*�%�N�ڜ=���섟��Hё���	\�:p�<B{ V��b�ssNB�`|g8�(Y��,Qs�3Ͳ��$[��_HQ/|�n�����N2�$��b_�OuX����SJ%�ޓM;B���V�1)�U�}U�����'w��]�i}(�HT�|�ȴ\4�7���b#�f�[�����s���W���h�u���hlNN�:��������b���X��l���.��@��d/w��ѠVK��:O�IGΔK�H�\�����U�;J�Y�hE3�X�-�-4ɖղG�u{��o+S{9�X:��3_�) ���]�Vl�z]��㠭|�֓k���|~Z3�魻y�f�g!Wc��bŤr��8l���u�¢�|%I�X~N�,Ma1�š ��k7�P�����E4�"y+�+��f�N\B�1�
�\����Gs�Ē�[Z���\C��E��GjD�#�@��K��9�z֕B�,J��UpH��+��~��+'�a�M<��H��V,�0��U�u�Z��:�nf�B��yO������>UZwZ�H�@�s�(D�\���W��WI��Oe�.�-��:ҽ�������V�&�k���f�����i����t���F���h~聹��1Y36I�9W5�Л��#����r�h��T�,}-��7�L��Uߊ���6��V"5���x�N]v�Z���h�'G �~X�ԶJ�ˤ�F�9�J{+&��������}ON)ˁ���aF\%[u@%�y;�HK�	��	��/@��w.(1�9�\c/bCJ�@��g��BR�|=�ayp��<dP�P:��:����;=~)�z���&����x�5ģ�w�x?6�su-+Zt��w@q
Ȼa�LXi�]y��0�\a�;¢����$��rW�WhV�^q)�'3�ܠ�v�d��9N����h\39 k�����:��~�C\o�y�]IP"�ߑ
��c<�}_�b^��9u
u�_q�'���G8]Q(����R�R̢�rK�"f�N�3	b���R��2]I��7Q�GY��ߴ�M���u�Q7ۨYF�O:��~��m�%M�v��+'&�/6 '_}�0�8W\�VMM�YUH����Sy�F�ܖ\O���<��N��g@,������(9!�p$R��ԖN�88����>�~c"��}ZgZ���d*{۩0-vܓ#$CZuܵ���\l��u��{֋g��6��&�����O����p��S�,����#��:!"���0@]�]fCx��/ʄ葲�$������و����'s�T�����@�;�U��tV	��K���r�����-��,W�6k�UÊ_~����7#����%�L�!i�M�>��aZ4do��
�ؑT��tyH�cIHT��H��������>KR�NIl�ڜo�#_]��>�0�wҬ �B���iX�`��8p�aۓ4Ϫ���E ��@�����?>��P�j�J2%R4qV���(�� �[U��pF;6�A�Me4����>�1v��j>�2;dES�=,��-��$meu��Pt��[��4�o2���"�Zo�a�yf�ҸW�[4!os�4+����E�{�[��sw
]ZQ�L9��𽑢s��w�/��|�x�1u�L5�9]���I�s��$�����c����&y0���Ϛ��>ۊ�Ձ
��8,5�tJ.=�ED���h<����6Ɯ̶�4-Gcī���^�!��	_ePb���e��j�b�Ӄ��a�y#�������7���1&in~i��~ΔJ�C�\X�qy��u˗�������c~�bohʴ����s�'N�:׏�?,���H��=����y���BlC~A���3}�����B�F��af��5 �x4 �Ì�3W@�m����
6-m��l�M^�,�.Ƀn���nI^����).S1�P���>x�G�� 7A�&J�Z�%'�)�������x����{�Kf�7ڴ��܎��Ay��'�E��(�w��B/r�Y��`���YZ���M2*�l��쒃�5�J�sv �Ոx%$�N�tE�:(�3*����ׂ�ղ�N��Y�>Gg��z��_	/h��,�3<պ�@K��@V��sPD�X�����'�t6���� ���->�j��.O�;.���`8N�J�=���-�2���xC���=���e����'�`,�=J�f?�J	
)��_��VV�.�����M�W�S�"O!�(�i[aqڜ"�d�hҴ!_*.�k.��[��-�o,��Ò1�5���RMF	�<6)i�E;�*�|�\��q30�,�C�����=L۹�2@E1٥1��h-��;H~[ Т�-ĒӠ�έ�9F���}w<��Ђ �7�8��{O����\�6���u]��MZ��뉔F��P�Z��i ����s�]w(���'��dq׽*���F�sc�t]��;�购�������ٱ;'Qh<@��j~:��rS���g�[�l��J�@��r�ꨊZ�6��.m���.tY�j��mp�䙤T������6�/�H)SA��G����R_B�,���;������[�|�vqU��RM�K� �3W�A����%/�t�/)�/n[���]�$T4���tѐe��D���+��yI�e3���A-ar���#��x ԉ̾6��J���x�!�&Y,�.�S��F/� ?[{�/#<�}L��:XB���Nq�Io��jb�pn�Ϲ�f���=.U܏�푡���Wy�q�o�}dt&�P2�T/��4m�S�/鍪G��J���`��J�����������N���q���F@{��>ȅ�rK� Ӿؙ�|0tB��5�G5��Kt���~�5�f�✉�u��{��j�o���?��b�2X�Z���2��|���x��U6ygB3�o��*wN�&� s�
k���f��ļ�P����)���9�z��7O�`��Bڀݗ�v������l�vM`9h�`A�B߇ \g|i�!)L8�	�!���K��(��8��!$7�Prc�����b��ˠ�_��R��i_��z������l�e1�EM�v7	;~F�ڵ�M����m�Wᶛ^ɸb�R14�72b���H��
���!� ����'��"=��>�lF�1S�	��?�m�*h�E+�2��&�,h���?��w�s7ƭ+��8��m����l��MB��z�]��>'x����-�kq��T�����B��&\�ѐ���g{�),e0.���毛�����,`�%h��!�Ue/�4g��k�
(�fb��� n����f�;yw��޺Ξ�*�%ǋ5�)C�U����n2�ȸ%�)�?��j��>�0�X��Bc�i����2�dL�@�a<YAƣ��
�ڟa�ȡ�%�
l��J�aV�A����3�Lz	�}R�i�� Ub�Nǧ�ax/]���<��1�e�[�	�I��Q��S���2��"IF,L}����e�����
��x���M����=Ԡ��sעX�W1h���Ӭ�9��q,u�)�U"�X�P���\=9�~~�K7Rb����tfp�v��eZ�P��צ�hWY��Q�e�[!�q�2Ͻ�a,G��Q	�S���ב�FE�	 >��7E�/�3�,W���-�$<�\dl�_��'�=XZ�5�\���,@�C��<��e��>:^a����[#q�������kf�c�q�i�S7��	:�����[�|�?~��FvO���:k����i6�M�a]�0a���l�ك%W�A�<�K�����X/S�k��&��R�,�[V�\�p�"
d��dGeӔfU��Lx	^�k�Q��B72�u���CN����qg�_jvN�h����z�@ ��ޜ`��z� ����ROp���V?�l/�X���q�e���:z����VUPI^s������KcS�C��`:9�Ib��P���J� !�$V4���<ڛ���|�K�h � �L#D�]�
� �ˡ��M V}��|n����x�ޡP�������6��2,m��2Ч\u+��~�{ ?��+�*FGw����dW��?�$Cp*_�͕5����+�����L� ,�"I��yT�"]���Xt��/�kqy.�S���s6�b�����}�b8�I��;,K2> ������.f���4\�~�O?q�ۮ`P�eg�cB�-0R���5�V��T��<A��S�e��Ǩa��K��&�qe�߭.��Ȟ����+5w�񂔩N��<@8����� &�}�J�i3���+����Y���S�d^��3���j�/��C�bg��<D3�'��^��p�v�E���㔱#�T���h�Tg5�76��r��ag�Xc�S�$�Q�.JX?Ҷ�r?~�2�O�8�\qO�_?H�D�E6]|���+�c�^3x^4��@�w���ͯ�nDk�q�|��*�z'��`���=}�v��fJ�Ï���5I��E/�Nq�����I���8��Z!���kw����LQS�q���,B����˥:F�p�&wg���#Q�������ߪ���%Ұl��JD	EB?i���e{u���/A�A��B������f_\��2�z�n���t>-�=b�R@�������Vk��������vF'�w|�vG8FhX�~��3Z]@�V���(���q��$�\y���aʫ�0��Q/������~�ܹ?OI��!	���2�ךS�6��8�m�I"i�}�
Ş�\߰�u9ssz���l�Ac��ZLVK�m<��� ���{8�����+�ga�Qq+'
?�>�%��e�S0 �e�\��N4�;dO���J���8�]�ӳ��_�AU�����ML�bKfbX����60�y�ҙsCK P�w4F�tvxo�)P���hg���70[�q���$��QX���H�Q�T%xB7�YYT���m��������S�;�J�3�_�`>���PD���=,#&A�u>\wۭ�к$n<�i^0{�k��d�5,����)p%�6ՅED�`�"�YI̧��&b��?��BM�h�����~���z��S�_4e/���3��rM�'����.���q�f��}�kZ2��\� ��oG����C�D���PR���!޹�E
o*�g���`:4��֚�؉(PK��Q]������oGּn�'�e��h�eʋb8�~���2�>�df�D�B�Y�3���e�?��$�EYc���$e;@�;��<J�O̾S�.8L��xj8�Y�
����B?
��1=x2���Kz|�j� .�O� ��