��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>%��}w�K���ē��fu�}vi��U�㶘�ㄍb���XT�$���sݜ1�=�5ޓż �+ןp����,��K�D�׺[��3�m�9N~�H�&\��D��>�԰vf���֘N��s����7�{�Wy0��}er�-D(,MH��)�ˣ%߲9j���qH�4%�MK&Jj� {^�|&��^��iV��(z�E$�Y)2��%�b�܏�(��K��⑆ 9ж�������1��c=�(�e���$Z�Xè�j���8�,M�>y�s9��vc�n�sm�^��т�������"�V��8���'��(%ٸ�:�����w�4�>��Ѭ�I6r���[�����=��b0�E-k\�NMn��[���Ő��lͭ�i6�I��}�!�` ۏ��{���T�L��F���~B�����ZY�t���ھ��;����U<D�P�z&�%FAɸZq��dR�.<]���GH�c���|_�F��������Rv�+?+��_�:e��Mv@�#���hoi]���,�x<�}�`��ati�"�־��к9>�(&�����"���R]�Ei|PE�����Н���6KA�7(2��h��n5܏��)��#<s9�U��"P������n�7S��ow8G1�+»��EAw]�C��#�y1��J�0�)�o�=֎��K{�D�S�z����/D�jGڏ�BC�A���N�@*�"�۶��_A�`R�R�텙7�9��LƩ���R��<k� �c�FmH���fT��QA04�'b���c@���Gu� �����A�"
m$r����/�r�O#ԍ&�7�z�s]� �Z�Gם��F4�6�����X��6��t-"X�~fc#�h����(����=j�R�g���A!4x��]��j\W�/���`�s�>�T3%�  ��	�Zol%�����2ʮ� ����xM�o��yVw +�)9�k����3o���T{�'{������+G�r�k��4��,if�6'w������	X��Z�5�q��8��[�Pgy����;,��J �|��}7y��qP/��-��zQ����	�Y9<�-{��>s*{��nR��p��8�D��oDy�̟����C��*Bu��)����������I���8�Q�D����)sD�'![q懶iUfjV�������e5l��rM!�i*xmZ�Шם�1�+X��R����x8G-}:�))�E|Z�g�ļ�n����,�(�X�H[�:������U: ����2L>���f֠�f���f�,=��N�
UȚ�������Y%��yW�!U���rh��� �H�������Y�I+pW�<ߤpO �@!.9���ީr�\�$F�
4��4c�Z����P��K1� i#yk*���z0�@-��/� m�)i�*a��	K���^�0��U����%�����Pe�������F�"���X���Q�y�v��p�H��"����^>��;e|�>�l�i�~�݅("��1���=�U�C���B�����6�u�S���7p�R*u4VX��/���?S��e^��l�h*�`�B�Ʃ:Qt��X�V6Fo��|�H�V�.�NPzjҵ��zW[��a��\&�h�2?�ߺ���	x���&�?�|��BG}[��49�5xli�_o����!�4N`��	=���Q4BO!Zfh̝~�m�%͕�RgS�Ą;U�A�l�2 e�|1j�W��ػNs�蔜ԯe;<$%�I~zzOF�dǆ�3�����<Co�"*Q�`���z��� '��>Dl�~��vי��r,`�����l�~���ŘϞy�q�oڰ���;���PP�]b@y�s��p'���A�`�D�B�+��?t�i� lz�eF���6WU�*a�brzI���Zp�ڴxT�բ���o�$8mh��\��L����l��%���:��"�G�9�1�%�����~pb��,�]�{�� ���隹��*�ִGa�B,j�$1�zڑ��P�<Jd#}�g�2���6��R�>m����,|��>F:�)�KL~��BO�W������h���"F?>!M]@<y7�����$���FZ:���:2`��:Ӛ���9B��a���_=�wB>p~�7��<�6�t𡅌S��B�̦�&�5�+�*�����(���4&��d���{��j45��\u(h�xK��Se��hP�3���pO^p��P�m����I)8�5X�٪��w��ː�������c�_sT��E>�ǎ�^^����h�Q����h,�ň@���y,#?
��ZY<�F����$pD�E'��.7�G��H��st%��c�P�U��R?�����݌u��6������H��(O>�E�ʑ��̹���{���l��^����(n�"���d�m�''��/j�uޱ{^*���U4e�j�f���`n�4�7�.C���a)m8F�*�0%l�b��|��dB6t3%�8��虘w� ��!3Ǹ�k	�&�:���o��+�0ނ1�e�/%9����V�辧��[+��d�D������8��{�^�l�Q�+��2׿v�c�}>hL�`ّ|��Ez	�|���ϵ�ݛ\���?���Q�g�pnW��1$X"���UHh�M���z��ɜ��l��]4��$;+t��U�Ld��p���B¼*�*lr�=^�dU����5�����!�X_3A����姏����F�a�6x=@��+�0��!w�
(��y�%0��	¹����V6�yx8Ǉn����Cj�A X�JQ��u�T[U��2٨�[->I�I����A�u���(2�q~��s`��E�������M+SO��p���D�\�h<���*xrt�1Bnu���ٔ�����
N�p6WU3C�Ay@9l�j	�YPu��^����_b���H�}���8��Wg�n�?��+�����>���n-�6�S�_PTgI�@�ʕ��OL��:E LI�f�
w4��x"��� d�L�H���q�Fe{7>�7��T��m�����Od �3.,�!z^�fh���=4E�S7(��i+��h)���Y�Դ���;����V"^7��'�������1r���~lԪ?��$�n�����j�������]��cZx2�����Js�o]�{����!���е�?F_����:�ҧ�����OQþ�k�������Ώ���p6��Ƶ0�l�C��Ln������y�J�.��z�U|�k �����]Rz�(��6���7�$�������i$��RRe	��^����5}"*�����~��`�]ÏnЗ�+��������#lS�D����A�*Ŭ[i3�:��s�|��o�:��੣R���	���ա��w��`AD{�N��Ԭ�!|(�.�h�~�N�j��I��$�{��Fw%�v���M�,.0c+:�F/�����M��٧�Ș���h�I�.Nr���$�[�+���6;\�Y�"t7�}�<�w&��j��D��} ����)��'FA��A���-&�vaA�~͒�_;D�:使~e�����ܛ�,�8��q�x҉Ֆ�������ys�bH�=|۸����"��,�U���9����� �.�7�����ŞG�W�� ���Xߺzw�?'�ΔF
`Ӕyo�����x���S��G�Nl`}�V�����6OLU=λ=�S#��_���׬�z�'W*��N[舸��c�7^o��ĵ'�6�"������Us��%�6��=uh�����Q#���xE��=>���D8^gF��B�}��'�\G�)o.��R;�����(���I��������넬 {��B��c�FW7��Nm
Z�q�M��#a�Ao_���|އn��%G���������׵Wc|�A�G�(`f"�e�+Sw�����ׁ�7�Gp�>Ȝ����2�O��;�`ę�ԟ�5��z��E����Cw�$M�R���x��ld.�B�?�'��[Ri6TY����:n�`L8$DË���(��!��#F�?9�-��[��G�u�<7y^C��<Y����|�q2^�j�&�t��:���EY0�����H����7R`�mBG�"�X��_�6���*3��;��ա��Qpl��+���>��rA?Q8B� S�$'����J/��V�Z���1W�
JL��f�*����~�cz�x�:��]��ē�j�\[���l�����e{�ݰ41���_f��F���h�{,W�YKGU��̶�1�����8 B����ow4�ƑX���`�����8�#-=QEL�̧ ���j�F͇�����kK��i+A��&
��( 1��'����w+1,,s��z��p5�W*�S�{W�+�+Ź�[��2�$6
�Р�������(tr��Bͻ�7�qjX�*v���:�
�֖D�>^�l��<I9pvz�v_Qh�s����������(`TCT�{(��0o�gs	wN��>NEF��!�ν-�n
]j}
-��W���U^��5*�S�^Ƌ��U ���#1ґ�NL��@������=�l��K,���ʈ����<�JA9Fr��R��;M!i�֋�{���Aʵ�'YS��:K��ba����l�.�I�9`z����z����tL�Γ�=�l���t�2�ZO
�b�%��P�w�����e�h	.�7��$�iڳ�*�k�x���UWY_�bpȩT��ă�Й"�. <x�*�V_e�M�W6�����]N(#�+�DT���p(��;}����hk��eE�ˈ�i4Zw��y�BU��7oP��i�_ؙ���{_1��{F)�����>�w@L��^F�kݗN�W���#f�����1$4���4���A��ѕ;��� �:F6��V�z�PMZ��_��.e.�O�G-%6��<ԍ"�=	˽2���"�
:	�����Y�gV�=���h�Г�,~*�E?��9�M��5�ta*T�O�!)R¡e��شI���$�x�j�ya��IMtZ�_�v�2̆=�s��#o��KXot�_�������H�:t�a�[�o�� �0��-ZQ<�槽FB��n���(��� :���ň}J��K8�p���ݕ?g5��Vw&qR�?�&ٚ[
C�дM�>$6}�N_�����/�Ƃ)�i��ԗ�u�#?���l��.��GQSprEvg�VEv�y�H�}J2q�J����v�0���O<�2�k��}�5�Ӽx�Gl��@����+^^�J	 2�?��ʾ�#$;��K��g��)������0��t1@���Er����wK����o�OY�ގL+��s �;��Sd�jX�̀H _!��r��X�2�Q��6�DG�Ⱦ�s�`C�x�U��{�L	1�S�0��:�
S�5th�?y���'�w�����,;[��遛EÛ7��{����s1�s�����X2q:�Yt7�J~b��z;T?�!*uA��U������9��jvo~��*͒����i�wr~b��_^��J�D����{�
g5+t����ɖ+A��G�w��l:0F��/ny7�.�s{~e+�ݿ�%`=] t���e�)yk1.=�$taz�+�"l�d1��K��P��ۨ��>M���v`�gX֚�Êٔ~@�����v�<�[~p+�Ѝ�<�5J�o���u��bg3h�2#�*wr�;��-�-&�5u�(4���bz�x�y}�+�Sc԰�V�Z�����2B�Ejb�h��ܼ<��*-S�02P0��zZ�)%�f\�z��е,󿖔�[��&�7�o��������U�RSe^ Ֆ'��� #|��bm�T�}�bu�Cwq��r�r�>���^��L��/xg95Y��b�������Lċ��J3��=+��2d��QF]�vR]?��D���).�]�@ ���շ85k�K;Inwswjw���7�e��$� ��6hl
�ӈ�������\�B��/�$F��-�႐Vk�f��*!�Yv&�M�Y�ag�$�&<��10�M�b9!��T�uM�{���W����.8���U�ȹ�p��>���Ϲq�����v=O��R)%lu�F������{+Y���ix�éW7Վ�2@0>��O&�+ֈ�3��|z�3wd�`�a;чL�
2�g!�'"�V�Ūk`����9���PC~�b���3�Vf)i��]R��@���E*��%����Q�~�l$�f�5�z��
����?i<����y�pVC�B������Py �Z�6L�N��������2��'eIf!!�Ώ���F�����1NOL�,Bk��������=Ζ ��H{������m���:���Ǘ�L�8�ٽ��"v��j��{>��n�0��8��M����"�]�׻8���������+�vƶ�귴����5���Pf�J\C@rj&�1wۆ��¨u�;�gLH�&������0�o�@:f<:X62q�o�@ה�O�[��{�����;\��۫�[��3�q�Cqt�}wٮ�����C��<Z���9pŁ4VP|��$`�Q#�� Y �Ѥ�==��ZA��Syα��tB��1��y��3���N+���]�҅�/�Ř�;B���I��� (�f?��]kP���zU���z��z���(��)�nL�1yQ\��$��K�d�L�xPCY�/v`�O�g�J;�Kr��2%�T������ϟ�:>�Δ�������w
��!E����YX����Jn(G��Y�|���`�f��
�y�;7;$L��z�-��]�8S-�9	�ߡ��rd�c����aF��|�P/0��륈��.o*$*�pw�$�.�����k�3U\t��������2��X��Y2 ��Y��(�h��Cg{.,�
n�W�eW��n>�t:	E�8�[��N��Q�ͷ�-�z�F:��l��|a�2k��TU4�B�5�6���]s�ػ?)Iͩ��%m��4�<���]�=s���f,hj��M���$��Mˌ�]�����Fq�Qi����z�<0�r�����2��<	��=���������Qwΰ*��y��ȯ0��%H#,����O�77�������@5�c���Q�ݻ���8,P~��)������%�ZѬ�6�R�4m�q�|"����f�ɈXV0/���sA'�6n A(����/��w$�4j�Cu�c\#f8q���Ϝ�~���y�<��%!�aO�� ��?F�0d�A�z��n���h^e��.3f��n��{d9����f�r:�iOFl�
F*�y}�ݺ#Jn@������L�\z)�M��A#ۺ	�7�Fz������9yhI��j�����~����@l�����j���ҧ�ᾉ��1��y`r�ܛ/B�?t�䓡�g�L�R���x�uƌ Ɏ�hm���`]_+ZX�y@���؍1�i�RurC�Ԯu c,낟��W
�<��9o�c`}y'5�?x�V���&��J`v�Z]	2gUᣬ�i5�/�L�/��^J���4W͉��Rt�=�<ݦ:���D�M�����_���UnJ��[� 
ޭq#u��^��L��Q�M~���\E*�nkE�y�Ə�R��d|��0*ޱ�03j�(�ܷ7��
����2��h�����V��l5�Vs��.���w�O1�q��}��}��F��a~b7��Wx���`�~���y(��� i�(v݉�I���PP	�n	���)�&}\���]��/ʓ�%��A�0&���ѡdw6�A�z��\��1��� 9�|~Jr���;�`����T�Mc�7<U\Ė����t�2$ņ�AR��:���Ɓ�l�F��Z�췪9�.��A.��7	j�d�S3kpo�#pf�J#.�ۋ�
Qo����j��)Es�%;��fy�z]��/��['/ߏ�K}��H4���u��^}��jyle	�ւ�x�ݝT�{N�%Hwl�9�y#���%�Qu;�����E����X��sj�*b{�2ɗ��(����t��õB/��J�2�+rW"v,"��(�11���Ҏ��E}4}�S�k�&.vbC˚�R.' ��,��;nM�R���j
أrIw��:[����`>�OG�ᶍ�K�N�?U?aR�d��9nRō*��i\�$��rF��F��N��܄۹�I]���J��"��'͂�r�t�C�&+�l*+�<�I(E�fb�r�MK��߮�^���Ő4�w��o�E�(OkY���W�Pa��ؑLl�b��\��+��ni}ε>�6���mIǵjᲲ��8|��-i�!���[��#8� ���I�5���a\W�s�[ФKo��Y��ݙG�k#� �
�ު�a �|G���A�-GOJ�`m��mՒbX��*�$Ӎ�+5*���צ"Zx-���]��eM~x+S���C䁩����\XƯ$i1?�[�}"�O����G������)?uh˰�&:_�pv�C�f1����,�n��g%�c ��ԏ�:]>z��vo����	��C÷��U7�VՍ�D�n��`�X�˱�\C,D��[n)~�ޓ�����ꋬe�MS�b�4)J.��Q�}ꖹ2�x��!�׳3w|r/��TV�@�uC(v�?@X����k�R�*�?��:���eE�w9A����FY�n���qИ!���]8��1i4�Z���'�qm\g�9�$�$�eXK�����J�v'���J�~������~��qh���Q����S([OzeQZ1>U!Qeĝ�~'�����f�Ș���U��w��Z�2+Bc&5J�3�x콌1��x��������"��h�F[��A���*�0_�6+M�E�
��(�h~�C��M������Yry����#ecy$H��4�\��6�G�T��e��x�i����[�}#��ӛ�)������O�̑Q�m:e��
Ί���ʴfD��5A�]a�B��A�$����B%�߁��Jf1�!>�S!e&!u�_sm�� �mfC��6��6���Z�q�&<�n���7X�Y�/<3�'�,�6��^>���t�}�f5-Ԡ�]^��.�',@����$GC=�͕��PZ���"����ʳ��D]|NȊ�\�h�޴%���WĹh�j�qNZ�wacF�����)ÇA���q�����u�@������zn�{K.�{kŪ�N����>�j�I 03��e6�T�Ewx�04~���樂�6�":��Gm�(CI�N���PA��x٘�k��?ٌYZ�xۚ�3P�Ytu��s]��7�:]I���V�҈;����X%o/0C٣ނ�DƤ��\������ʤ�lEX���!�]�����8N0��,4h2��^f�/R��ͼ�)|���Ϥm��L�r���_�N���8շ��%�Q��@S�5	�]������'1�O+�x�B���꼌§�-�Vޫ���R;��݈!N����޼cB*���:oR��E��&�]ق%��ϒ�:ib��*x,p�y�t���={�Y\�*Оe0�l��M�B�P=��^��Na�6�n�0�>g��tc�e*e-X���9���ݖB�PhP�2�/�5&6�1��6Ry�-���b�ma(���$��Ͽ��M|0��Iy���G��&0�K�f��z�Z�M��uR�H��KӺ,��&���I����)���������n�k�-�c$Xxa�ks]W�� D���$?��ءGj�F��kZHz�(Ԭ� k�ޙǝei�J���;o��(+�ӹO�H-��f��c'�A�}���d#4hh�?�=����d8��)"�����w�b-w�	'����/ػ���+�%�V�:F�~m'Ƴ5x3C�ଛ%� 6'*3��j��L�Z&Y���mfM:���`.�?�������͍�!��M����O��·<U�H5N�.�'g"1�������ʿ/ �T�R����dJoj�h>�#��>򛰧N�v�u�W�;���d`1f�n�n��=\�J�9>�_�(��e���4��.`"^^Y-�6� _x��-�7��\n�E��I�j�Q|>�䕼�GHIIh:��3��P�B�r8����s�����P^%�Z��7E��W����KU�`O*�27g�����N��HM�i|���/����PJ��AF��%���o.��~o�Ts�~L~�f�< �'���h	���ye��j�-~��XM;Wv��W{0n(�Q!�.��?�G��E��Gr�#9��6[g
)\�̬��V[�U��n魷h�>�a�ۿ�G��������y��~�7�J�����`O��|q��Q��r�flg~�{nț
��R��dh��m�0�g�	 T�7i� N�\b#�DB�H��4�0[���)4ɧ ��CM�w�8�Ly\}zG\o�� ?������|�86���
^�O_�CQf��R��>�Xx�>W�XC��<b���V�h ���஍��7����d�>��嫐��h��'�z>_��C�v���a��'��v��^���]�#�q�)ԥ3}g�9;黄Gho˿ ���U$������pdą����,���(��ɓ�;e��rL�;�������-�}7��r��ȇ;�n��<�?注���+�
t>���T`��W�c��g`-DZ\�F8��P�-Z�fR
5L)ɚ��u�Rf0z��Su^�_��j��LgiY ��5bm��z�(Y|˩��e~gs5;�+�/�8d����N�E��';p>|'w���#)���+��i�	�Zh��Py���%�� �	�ԍ�y,�M�#��inu�L�",��M�M�C-7_�'3�C�=�y`+�8�V��R������.v2e��[A��`��[�ͳ=��P������}�FC_c��R���Ƴ��_����r�}1��V �v��=��g�<��]���3׻��H�pxR�|:��ν�ùpW�i��:t�PI����(��hzD����gB	�-�CMwm�J�'B�B5��d;p*�$M��ڀe��'�Ʌ1 �84&�����W�!�8]�������9,�"�%��'!�a��Pl�q�>�ŏ̍'�M~]�P�ϳyΣ�Vi*�A���ĮD|���7äU�t�p�r>��B~���#E2�"okl��ަ�Պ΁P��~X�?���0X��Q��K�8�84Smai`7�Q��w�W�tW`2a�iq��]�"[��m�!ҕ�D)�Z���qp3�3`��xB]�n9Ü�Z"������cq'/��e��nLIkN���8KB�*�W(���i!����@H%m�IR����8�{X)Kz