��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P��v�"<ߞ��&'��k%P碶�R�ӣ�sĞ������FY&;k��e�cO%���B�0��Djo�9l�Y���z�m�&S�[�� �|`�kK���XD4��_x����r�O1��Q4� !��ޑ��g@��U�.�Q5o�o������7�"6�(m+�<%�٘��]zuo#�g/���lB"2�����$)�Ң���r]%�� L`���Y'�,��$�6���\��0nG}�)�`GmH
+јv�:.v(�L�q���6�r*b~��M��	Q�����)Q��{�U�,K�]��VXԘ1i���tI��J�9QZ�	e7m7j�V~&iF�#1թϣ��gELj�TN��7)� �su�����*�r��H�z��{곇�9�&ܘ��0�v������MX[���H�$�,������2�C0�xH �'���ˉˢ��{\M��m�/��l�jz��C~ۧ�F	27w�װ��D|�����O/3�e%e��t���V`�U��5%ef�ѸI9��=�fOE��&��$+jj�\ѠW���,5w$��]��",d=�wni��)�|�L�c2H֛O�N٪�bD�:�����ݟ@[4�&?R�������g
�6p=����-�C{G"�_��?�N�"s�J��\ڈ,��Fg�"1�k<��a�ۨ2c����
vl*�ZR⋸H�80N���T��L.=P.Lpl�4qr���rG>
2/�;�)d���������"�gUͪAy�T^��|YE�S�Q��[����_�K�%{�_G�g�LbNB&���^rQI��ب�aR�bD�Q���̖ƅx������l���f9�Lz��K��3n�}i�o��f����Q���,�5��U�=j�5kL���[�~mup�eZU��{w�Mĺ��)�i�����I�h�4�� 	RN[�g��������G��vϭR�L�{��joΟ�u�K0�-�T���]H��n2�a��Ϻ���:�\Cm�w.$�+��X�QB���Q��-�*�;���� �`e'.3- �R�ߐ�x��"�
��D6`6h���z��u�y�!�9EK��.JsZ:%���c86�Wu���5�Z��}�T��$����w��NY���s<F����l�n�C��f�����DQɲ�C��~���2THm�d�z�׋p0\�o����	l�͘j�Ŋ��&��0M����ڜӟ�?4t�	������+5�*�#M�&<�͉�{��8	�ܺ����Fɼ��S|؛�Z[� �-l���z����#���	Xb)<`xቹ�s��T{��xn�g%N���g"y���l���٥g'�6��g�]��������[fD����;>Q6CM7$*Wأb�"cոs����ɫq�C��8���vѓ�
���#\Ӧ���ղ����m _~�J�jcG$eUd�YBxR��"��ؠjkx���ʞ�� ��${<�2�)��9�L�b�Ƙ�h+wx7���$��5�5<_0�4uBc�pw6@ż�
� ))ة�W�+��B�j+r������e�B����)�&uӞEF��+�<A�&���L�9��a�G\���|���wAh!`�ǝ�`���H�i���5lq1>��2�&BM2��9�O��T�5�
���c$0��qyn�6�G��g�#=�/u�B�,d�\�����̍��>��CG�|4�sWUp��i�jj4 ��e*��o¢V�~z�A��������a��fq� �"L�~���\�%]�3���A�ef��W�04 ���郜�s�f���
hT�V �F�$���>�3��=	�7.����X����\��nݪ����e��y�&����Q��
*��F�OHY|7�c�4���&=��8MLwֈ 23�J��D���D��ʲxB\��,�>W�2~ګ2��YS)������L�� �����f �ވ������>Lj&vr���M�����>���*��\>m��1����Z�x(@ݧz���������x`ş�?w�ͫx:5���%���dJ4��*��\,�$Oq��\��d|a��I��x����Ϲ���TeH49i�&�
W{���zX��6��?��_zY&W9�є����B��2}�#q����C^��zDծ�f�^i�I���p�Zy�$�.�>6Y�[�)�s�:!�q.�X��r��W��{�lM,�[x�2P<3~��C��jJ�p;���C)�!��Q�H�R������͌�itH��/��[�sD���(�u\�c�d�B�����0Bx����\rT��ն� �0v�v4�)��җ1eS}�P)���:�}  ��s)kv�gD�z���ik��dY�;��<�ȷ�q�2t�>5����(��1�����k�и�O���@E(���}? �W8�֐i��Fb�v6궙	�{өb���f%a�gS6m�$)�X�k��c�Rg�&꣢T����u6��n��eY����>i�!��GmL�6���@Q�բ�LL�Qq�)��f��wt��O?�H��3��\{�A�zJY���F��զή>{�q~Vh;��^M��2CD�u����$��	r_������&Ǚ^�`�r�J]3�{D9X��no�GV���6-}N�ѷ�9Cx�����a� ���k�ϝ҇�ۄ��[�{�JP����*�Ow?t����Wqon<�?IMSʛ�$��D�0��v�?��K��Dіap���P!�A#FnX{�`�^[¦x��=y��+��{ɱ�L�z�\ӄ0at��1��T+�}V�N٫z�YGL&�o��t�m�Eeu}�r�m�#L6'��z�) �&m�t;�3��:�D�ߚ�����I�,7/�\S2S�����>R���W?�y��;�1-趶���6A�@�ȥD�#/�W�B��:;?���
ys�9�D�E��E�h�rbX:Z�XK�w�+�H�h8��c��5�ͬʞ����1W�*�F��.��ք��'Z�@�Gk�i���Ҥ���sM�J����&\?�;�x�e��iq��B��X=qp�s���N�fy`��0��wWy[�b�VK�[�������C�2��$Ŗbڣr����u�]>9�u�����~��6�ؕ8
�`ڔG����<�^#�̌�K�v��E9׍����:F� >�a~�Ѳp(�(]��t�#]+�۳"����G󷃟�Xh_�\����d�x>�sm�����w�}t��"mg V������I�QE�/h��K�ۺ�؛����P����L@��PCY���Uj�N��x�z�L�wƬ�$YϽ�ndvBο��ȭ̦kI-Hu�ܒ�S�8�#��C���T^��&R�-�o��_m̆+����������Zu�8�	�OB�Zқ�c�Y����@��i,rqԻ�����=õ�
�,��Q�"�a�t�A"g��|�Q���01�E7�E-N*�K�s��簹)Z�&W&>
9?N��?g��/��`�pN_��lGh2N���{\���@�F�R��j�A����h���
:��.�����ɓF����$-n��jT�p]qc�f�I�|�FMߎ�O���g �.x�Ts�n��it���@�m��f;:R���Ym��$j�t�D/Д�Sk:�5٠P��>����h#�g�W��΋��q��܊�2z�+�80��)T9L�R��W��$z>��W�|:�G���c�����/�q�(�2�����&��͉��g�"�Nano��T{� �0x}�y�&&�I=�W��t!����"O��X�.���X�H7в-�ҝ�/p��p�M\D���[�u�>�M�[���t��c��Q������X��8����-9��`�䪪��"��`���K�ʥB�Z�K���rԳ������>�+s�����7+�8��z�r���V)
*p4r�|�MH8R�>�#����q�!X���}%.� h�\�Â�q���Fc'9d�ڑh�=[�¤�Z��c��d��k��i���b�RJMw��H5�h��SЅf/�����Ѹ�ٜ�E��ZϺ����y*u�3ݜne����g��4j����7����%�C����Ox�а����v�����:P�o���_�8?����A��\ƨ�]5w���ʯyq���K�[gC)>��z��~3)����9�U���R﫤�O�ռ�2�s>�7k��6r��z��M
��'���bG����� ��";b�^���t����ͳDyPNl�6�[Õ��`�3{���@	�x_h����YJ��\;R�j��>�2��K�p_qG,�������du4/$ԪV����sd������Y\�a���Ͳw�#�|,Gia'8��k�)�~JLHns�>I��4t�����{2�X��F�dL�����Sq�'21��2m�im!����^[%���S�p�{o7W ��qᑞ����|7�ѿ0���������Ժ�s��`*"a��p�X�Q"�S����*�߯y�
���a�v�+���k1G)�n��W�Qz3L�G���@[��|/�u|��K��������
,���ݍ�[̘;��Դ�����(�S@�Ȓ �Ɵ��{R�j�}�[���d�3 x�iKL�=+�_�����m_�ҟ�	j��@%�S���l������0� �L,i��C���Ӎ?�r����Eܺyd����J��cޯ���oh�^A���
�~��u��������}+W�3j���jr�����_�E�k0�ܺ�U�8h:&C	t�`���F�Ű�����řkpDʹ�y�r@�s�W����P}n� *�eL��C7���"9#�������D�3�H����*�W�<?����>1l�K�h������Y�R%��*PžB�|���7�]�@�}�ޱ����� �j�ӍAZ�F�<�+��.ʳU�c���0��p��(���y�U1��1n��g�&�J�	�Jf0��z��w�؏�$���II��*)�J��N+�����4��e��� 4���>;�O�=�I�A�[ @ka���q&�
��	1��X��G����m#���-�os�]���
H�[�Hv]�Q�S�9p�6����'ԵaT�1z5�X�������蜵�tlۉQB�4���l��A7��cԝ��h� �+�����51�X�)`��$ʨF��8�r����7�_�r�$�Q=z�i��L��6�ނ�Dw����y"Q���&�!m��W���ۚn�!߫ �>��K^���F��Z�P��ώ���ÙWn�� �i�'��J��Dx&�h`���-0���9���'�N�V�W�X�c!~����7[��nm<��^(��&�������p�&H&*	<�<*[�)���+��'@�6]AM��3wͪV��x��a� �ұ���$� �]�A�bX��|[յ�ڌo7T}ѝ��Yޢ@xI1�oh�w�ؔh���"R���g���s�V-i�`�j�p�eL�����5��)%x�AOc	�IbY+HRSc�R��J�0}/�ٽl�����Su+�o3����4������}\̛m���,>8���$y�܇p嘁;8�eǶRī�$v��9���hz��<�
U,F��71)!�-�#)���<�ED.������C]�5��n�f��pO���h�u*9 R.���i�;u.�E�!y��f����Gh+	��e��SFG=*	aʀ�T#h�a��6��E���,o�(��JO�r��*�$���;oʛrZrB�*��F/&�99 ���s+�Z�NP��C��S+�U���gϨ��V����-������g)#g�����%!H�(/nP��oڮ5��b�,�h� U���#_�Q���-�0׬R�T�>�b`%��ٻ��ۏU?��
�т���Z!��Z���7X;��T��G�5��j�{�]��+.`�W���g�:�,�cx���t- ��|$���Ν��N�F�'��J9ۥ3�j#��ux;�tp/ݒjk{S���(��|�蕪�?�����\��X�T���,p`��+KU.�̸m��U���/��0���V�}��ÃmI�d�B�NtR��]�G?M���?9%�?����˰�Ջ<�>GvE�H?̑�(1���G�t۬6��Q?�
�� k_	�TF�y�����'��Y�,\ŷ�T'�Kv�<K�h��͡�?E�J����o*0����GV�R��z����o�D;���й�q���X�,ME�S�n5&����Ѧ�<2Qjr�J����Q����O�h�]Wz�s}�7rf�d��;�Gooy�G��
{"�����9d�C�tP]ev����¦M�7?����
��N&����7�x�-���a>P
�lmzF�gF�P,=	�LPrI$f4�Lୠ�c��Z}^ �i�Iw��ťB�P��a��fnB��J���l�װ�< Ycv�_,�<�v����t�gO$��h(�@*��oJ!1y��A�����C$ע�|:4���`i���e؛�qӐ9�?���ZۜK+��1�?�d71H]�>��P�9$�+���b;��K���L<���]5�B)S�K#2�}�J��(����/n�M��A<��~�X�`g���%z
��e�����F�jc,E1�� W�p-^���Q�xzc|&�������`߅I��pm-��22��,QA.S[r�@2���`�7F��d0���@�}5����d��j�Z?2L< ���)��
jQ5��e%��*��Aa�:��لSpm�$L1;R-�����:4�z~z����"~�6��}PK+R)�ncaw��[8��f(�y������]U�:�y����z�r_}׹�ww�1��z���"���w e[���'\�g^S�u"۟�T�d�~��K��(V ��@�Y�I�۲V��"�CL5��
����)tz�E ����!�����m [΂n�J-�<[?�x"��[��az�L(R�g���"����-dH���6SF�|*��( 9Ţ,Z3,����E�����/������;�M@QP��Y����B���%�3t�W
�u��G��=}�P�U�9�Uq���3tz�QS��E�W=��%10�6N�D���؃9lKM`r�&f�I�l���/��u���݁�c��gl�S���}�u�-BE�0)Ѻr��q�}�7�%���,��m��ĥ������蟴 �����w��NTZV�c_/8Շa�s���h���&�K�5���h�@��L�	L����O�#��C�~b�G֤���O�l�t������3�����F�s;�{��f$��l¾2Z��`D�m����D����RKH����&ax1Țu���!�
6K�b?T۱�	ow�,�7���j}�$[�L���m�����R'��̬V�0�}U�6�R�O(�a�섐"]��.�m)`�VF삶AÊ���S��ة����mF/�����{��~`Gp�kO����<(Єe�1��hui��G\�c������1������[�:Cu�y8���r9���+W`�h���fwW��ؕy#��tx���:-������в8ۘ6}}���`�{�4��v~�2�g�b��Xk(ƉW��K�֞y 	'd�C6���<�!y�۠���e�}J�D�XTt�j c��?Chj�ϓ�^8H"KdH��aG����K�bxZ�+��j���J}_�Ŝ����T&����Z�aZ�
���iɇ�N��p�qf�-�M%;4�]R2vȊ���Z-�c9�uW��D�'ʦ�sN�1��76��'w낒�\ .�����O��ɇ��X���WG �#o��\`'GKۿH|�� �T����0���W�^֤�M�q寫[�)�[1�*پ��W�Ϛ�?xn�]�^L��_�Q��ӆk��o/&�_L*m$Q%���;[A%o��?1ɪ!�.ld��^mi/�v}��d S�%d�Ӂ�D��U����L�掦$���_q��"0nrG.C؃X^�M���t��,=�n(G ƊҭʭeE�|�6Ĳ���viNS-�6)"ߟ/Ú?�&�9H�%�
�U�e��xTv��߫�h�.�kJ��F6�/�WL;+�Tx�D�/��8{����,\�B��@�n�K��L;�u9��h]��� �%�H�)�Ĩ7b�Bb+-�)�	s%N�8Kn'��0��G|�x����cR�"D�ۚ
j�]�ܪ9�k�Q��m,b���gw���|���)%���.a3!CoE_����;Jh�c
 _h�8��?^MQ�vì�?�g�q2�._d5�������R�>���lO��M���p�3����ab%^p�ʓ����zk��m$�;�mb{�~C�N+�v�r���,.���V�J���u�׾��C����bҎ����5^W Jğ��N1������K�3_��|��s�f������Qk��W�P+��Ͳ��ag��=����>݇P�ǭV��3}��'७Q��_R��Ns�Ԅrv���Y�J�=�&��z֪�� ���,ف�P�?+3��;�5Ưw�#�eJ�uH��*;f��t�b�_}�#�a�'�ZO�~˂� �5��SV����X?�����F�wvt�]�iZs��$���l�l)�.�>�.��_K鯞G��Q4ny�U��P���lW�E��ܣ`�qڐƢh�Ѷ�&饮G���H��yT경�[w�ڸ*�wpa�yy��}�=TL��:�%x5�R�����G�YH�����%~�	o��F���B#�!N��o?���<�K�ۄ3�������s��:66�ZF�UQ�|}�"�0��G7
���wh��ɂ�G��㠙r���6�,GH��T�AmOFȟ1o�5C�+�~o¥E^�#���Ck�i�>�FQn��C�*|Sx��P�M�zu��:�骤��y�o��J����Af̦+�����F|�W�џ^i�Z�(�[E�k��;t����4�T���U"9����������p�~oa%��َ��������t�9`n��C��k=����5~#�5db��'.\����Ng�8�̓��} ���)$��q M��TG1�h�x �v�lO����f �\�W�����khF,�&��Yc���I�O�J���ڋ���B�.�;�Z �+I+���yj�erQ���x�^��k	�3���~c�=?��W�=��Y�K�pj�T��t���������-QJfǩ� �?�2�I� E�(V&D����ڦY�2�1XEl��ƃo�a�����X>�i��ga4,=7���c�ȸ|~?�}��f�����G����Q��Z�r�ު"C��#6p������������V�ʨy�Xmp��ћe-�Y���`��g[�Ĥ{�h��Њ!�Z� ��]�G��/>"�$�ϥ��/��g�|�d�����_�j�稊�/Rx���8?�r>9O�@݃�X�N�;2��pK%� �8��r��?���a�P]_f���������y�ɠ(��`�萰�M��p�d֯���GM�AVtߊ��N�#�L��	wT���2���,E)�����d��%��ǴU�϶HT瓟�"�q�.�~Zt|>��,���Ҧ|u���#�� ��F��j�hx����[��ĳFW.��N{��UÇ��_.�:�K�$`X����6�
/��Բ�Z� ?��AR�ϗ#���s
�1�b6�+1��
�wLbo�Z+FK�Y���%6�7J�,zMg,�I��Q���*��������+�����v2f>�N�n1�.�RT�@N
<
`��C`�ɋ�̘/�3y�y���W�.�e�p���{OX[�\�n)�tf�?���5�"@��%��[�3����֡��g�{D�`3�pJ�J��B6��L���
a��O ��,� ,��1pC����'H��L@��ټ���+�짘���0���n��5l�W`�
>�K��ܓ�*屹���$���y:�ƹTR�v�{���E�[�+)� B&�Mv�F����EҍGX�	����Ӫ0��a����
#ȫ&J�ֽ�ݺ�k�ls��S�p_�C�CΪ`��qu��X��y-u�5K�foN��=��q�5���*Ӄw�ԋ�)�ƕ�����S���4�7�e�����bt�q�$Ɨ�fS���%E������Վ��?��#O���?�/^K������p=yŹ�)y�E߬���.V��r�[�������m�{ڥ5�.;�^��M/�\x�^��h���t+_�(Fbi�F%�j�O���|z���I�Dq�,U�"�g;ǉ�[S'}]2��>�]�?�y-�B������d��A�����b�Ϊڈ_�F ��%��eV�(��RЯ;��T��l��#f���+��|�a���%m�,���^�c ��� s����,�B��ޟ*T-�5h�@�
����ň
�L,ғ���T�O[ϳ�\?�sjr�N��E��?�Ơ~�� b�#����?����Դ����>t���eJxM�$�بq*yX4�e ���\�W=����3���҉�dZq�	�3y���i�����%���A�ၩ������슜�R�.��C+Tv>;�@�2�|�Y$'d�:�"�.�ڛ9QX��m3�DZ�c�8@0X��&۽���/�rs�R6����@ja��St��@я�L���w����3��0eȴ��48fܾZ��XV�>.�	������.H�����5Q)���E#���K��eZ��� N��%�j��(�ǯHM�ÞJ@�m�bS9�HW��ej����<��o6��s*n���mT��:���f<m�Z�w"+ؐ[U#������5�Æ�'ۛ5<Na6z�qf���x��M���z��D�o�֎L�[��פ��hQBLnZf��̊z����|v�ǁ.^���Ck�����6���Q򦔊wS� �
-tgElY}�Bg���0�xnϦ�w��m��:��~�W�9����V�9,syXhF$?�)N_[�Rj\ w����|'�|TVD���I	{��8@U���ڻT�HY���o��ޑ�����ϐǯA��IB��n-�N��엍Ξ�:��5?�i�ժ�oC��1��Yʩ�*�
I�V}s��$�z��/0Hm�P��6�3�j갪�X2�4J��`!�4̍f���X��U�N�L3�R���f/#(�*b������p>���`$&
���26n�
g�^ z����u_4�yz�ؤlLn��-��I(�:�HB/!Z������	C�Ԉ��By�W��h���χ�Ci.B`�h�m�&�Â?ѧ���e'h�m*ODi�057��4�ĸ6V]q��= �LlYi��Ў05fH���9�l���t��[/�8<b�����,ӟ����yؠg�/ ����ES<��#���&1Jn�\j����F3,�������ZR4���C����-��%�TPI�"ݿz����y�v��A���-<���z�<��5Q5*~~���Jߑ%��M�T_�Ҳn�z��X�S������n��}�r���������������!ؓ��[�X���<�>�)�Y�$y�x`��w�.r�������7����9	��[��0����УG�y�������CmSڳ��Z�G���߿�p)&�q�����Q�����J�/z;W[K��Զ1BK�PT�\��͔nT]�Ch�1=�Nk;�@�|M�a,c̟╳��S��r�c$�2Z�d>��r�s�V&���
ZU6Dn��^��=fg�ur΂� W���r	���ܽH؄3tCђ4�i��PϨ,W��H��P�u䁂Ǐ,�)��V��8��`��ZLK��]�#�4�$��� R��X��`��3x2^:�+vʂ�e���LW+-d&���H(�M�)7*���9tA4�;��[و��j��!��B%�;���D����Y�+e���sPs�,���U��ӭ�*Ko�n�ڋ����)�K���N7��c=&����Q5�}�Y�v���W5�lο	�@F�j�Sσ����I~���ͬe#�g�2a]N�Fb��]��X���rb/��R��j���#��ނ4�(kM���&�l�D��{�L�$ɜ�����S~{�d�C�=DK}��iQ3"�����CMU����%�;���e�s��
E��Z\�1n����ߤz9����(�]앤����Ϗ�T��]���M���q\%�B36,�t��2�qw�-�a�k gJ��֔�C�f������ܐ�L'��x�|�t�����G���29t� �%���H�oJ�OO��]L���(
N��qH2���J����sl<�65G�NK#h���g�0+O``:�k�5��`4���K�,�h�NR�����3��Z.a��E�֗�Z��d�Ű�J�W���5R'�:����Ӌ)��J��\_��,%QW�[��:���B�'l��_؂;����
=�4�H\��C�1�$�>�fF/D��ց�D7,R�m*��2�e�.jm�:��s{�Y1o%���(��T���gT��"]Д�)�i�+��3����s�<�q00�~�W��Y�56��p����A,&���?��QOV�<����@�<Q����0JĖ0p��D�yj1$�V�����RDUW=�ˇ�ע��{4
��	A�Pv
i3L�J�D����$ɨ�'A^f)��E�'͂�8�`]�ӧ��d�'���H�i�!��Ѹݲ>`q��o����߽�����TS+��X�	E�5�d�UWXesF�%�*�M��)=�7�ݘ�����췓�=����odx��~���(:7�:FV��vW��1I.ߑ�E����7r�����;���&���h�q�d�l����Yʮ�Ą�Z�E�0�l�UȢ��e�M����J��ɞ��ʺ���2:
����/t��3�r�ӑ*l0�U�'sRy�ȩ7A�EXz�I����ܤ����I��p�[-��Y:ߢvp�X����~;�q�t�:��S����@7�b^�L�؏߉K��PZk
CC�+��4�uNs��t�^9��;`�V.�T7T�h�LE�\��`,������j q�q��4	���݋cp��d44R���~zw?B�*j��}��������ou͸dd��j��<=D:?�Fɾ���	�s�o�VD=�ۛ�����	E��; ��� K~�E!�9��\~��2k�;7=�l�IUp ����oW
�:�2�}�^�<��Jz�!�R���.&)>���uh�F
�2X �s�Ƀ���M�E�VT��JIq	�߬�n�� b���\{�.��b�T�_#*}����$��7$䬭W���Fg�7�,�ʠf���!�B6$_�Z�xSV�]�ΰ�;����vO0����O��~<�Ҁ�5B�Jk[���Z��J��t5ȧ������n�X�W,I�����r���2�9Ʀ"�E�����������)R�PD1��#}�i�4�Q�G2Gp��P�)"2X���&�;��!��ʼA�~FDE���!7dʅ����.�s2ɘ�F��J��'A��X��'�9�M��!Y�r�}��'>꾄���4b4��}	�w���Ө(�*&�JwE��L�N9��\R�η���gd8�b��%1�gtp�"zC\?Q�	�!eߴ��(+�h�M�����8��vtOa��V����1�	U�z��
������9�5�8����� �-���}��bQO�S0l�q���L�g=b�(��t�$�JK��4Vs�o�����M�����F�(���扏���|��XV�ׯ�F�k?����/����n��?��*F �\�"A}]b�9���y�ѣ��6;L��b��|��U8ѳ��{��@�Xf<����zB���?!|-S���e�_�Q���E/!u��9�c�ߘ �j_'<�op��[�x2�k����ua{շ�^8.�<��2H ��'�Q:��j�.T7tx�6Ǽcf=T�X}��%�*'?-��;ʙ�y�`��Bu�:o�	�o�8~e�W$֒n���V|�9�a��)�g?`���D�Y�c��@wȒ���O,��1pH����6����ez���{�C�ژ%�����}�A�д��Y �vN�*<����g�v�&�4ּ�X�4�	����!�����ױ0)�"��*����\��H�S�6�f��A��Mu�5�qP�1�	F��E���s&�gkM-�iU���]-�Q��6�i*ۥD<���\\T^�'����$���&�����9��.��x>�2k����	�|�/�7��(�^0Cm�e��3�:J�;G��!��.t�C%Ӏi!�M"h��|E��z����̐﨡%T(�������.]x�y���&\ƿ���r�Hb� u��.�]F ��_'�6+���s\	ꀠ;�~s5J|��x 84qp�Y����tUk$���6�Q	�Z��;U��D�����بZ;a��`�\GJ�Q�XL�iGBV�F���Y��B>�C+��2E��p�m�����f�V��2�s'?Y�>�a�A��ׄ�٠�i7�hx�� $e�:����9ȡе��FP�I�fL������y�P�xY�=����!4�3k���0�<�Gd��u(����*�IS��{��ő]�"o��H�.P�{mHx2�����:�������ŔŠ�D��@�W�ެ�IU��6�d�P�U� A�	>Q��c�%�UE��϶�K2I�����	20G���Tey�n��e�^~+cW�bf{��)��O�<�ԩS7m�d��=
�kz��Ҷ�z&�볡G��.	�6���F���I(���:w��.^�dG�Q?��A�� �t��*��׍�/��&�S�ą����v�6D�GE�U�A�_V9��	`�u<������ojGa��ނ1o�L�Q7��bt{��vK�j0�Ll�q�3=+8�Ψ�Ie�2vN	���nh�������q��CYhią74����O3P:f�N��+r��qXS����=�\�5GG��4����h�mԨ'u%��'�^�xX~3"	?q 	Yu7�h�/G�u����f�QR�b�k����{��zR��\���� �����&f,�nk:3ic*>\!���W�w >��٩S�;�\���,~Q�8P5�D�4bIUGCho����	��*�A�^�������(�u(�~�Iw��X���`Qtĳ��m����N��|�ns��Փ�p���#utqD�ԍ�#�N��^�v"�^y��&����G��K"�����R��=��$����s�9�U��j���A�M�b\�`&2��՚��oR�- �,ԟ��5�� �k92�#��Zԧi��U@�<�(���R��$�SL�/tN���{���5���mR��G��lj�:�i���[]O�m�Aq�蚧��І�'�c�9!�3�++ZP��!���ށ!��*���܌��?�Y��9K��7���#�%r���ú�ZZA�禹oU��5�͸o�����N�`wa+�Р���<_��\�}�M������Ɓ����ҧubX��{?ͨu�<�����MnV\@�zqDlߩ`!����d��n�7j��C���'1�����~�N}��s�m��Cb�Ѯ�Go�����5�5M'�w��Q������QV͇�z�s���㚴����E��y�ln����y�۰�43�ZH4p� �GNa�;��Q3���D6�N��j���)L�sJM���c���D��\#��`� lZ����m�5%�j0�����69��U�"�z�=|bXd��J�:7�Ȋ�>�����ɘB7���qi{���A�H�i�V)-F���{w9I�p�}�$��\����(�|��7N��ʓh��-�2�4�࿄\������s�Xf��g�ٶ���d�#��ռ�R����Ԉ���6?%�{����<lKTE��&^'�}G ƓJ-+"k��E5ثK>�n���� ��mhu^�d�Ŵ��;k��FHc[�8U"J�Tk�3��X�qJ?�6V��B�p�[������-Ř��NS:\W��S�3��4ŊD���4����T& ���_O-�6�S��5����h�J^`�^���d3+v���E���x^�m��3�%)�h8�����c��P��4�=�s�b)�W]v�n��Ձ��T��F�R\��/Ƣ<�3��4El���[��eU7U�,���'aB������d:�q{ݍ�=cּ�܈�4
0L�1az�1H�ɍT�qNӲy������-a�˄i�[�5�����K1��=�>D%��9}
�2�eU&g�P&
�W`o�����x�x����.:�d/HT��;�Cr�#*�v��[��m��l��8�C�� s� ��>˄oє�<B�EN�Q�	�GY>;��.�4D�O�m�8�����R�%�W�9q�"l�lf�EvcZ��#��V��W��P�h~��p鎂�.F����!�^��E�f�$��h,���01��)_hi���e����S�V�F[z�]�U��3Ƞ5g&�FuXG���w�8+vE��1Q×�|TrF�r^	iN����ߛ����W8��c.�As�K��4 s�m��_�FU�����M3#}�����lڅ���S��G/��&�Tg��
�^�#:¿{� ����aw*t���ڪ{u�ӌ�JPb����}�=�#URN=�=׈���=�� jr�َ@�o�9P�-�*v����'�I�Mh���c�j+�����\�|z���:,��[��u�iM.-y�dl�x��C�6<���jw�uU��[��gbC_#����t��
۰�S�i�p����]��j07@���CL�5�4�W�,�C�_��W4��hk4N��:�j~/|x7;��7_2�4�9Ȼ�5/��'er�AX�e�jP6.{��L8�n��l��L)<��!g�^�z+_y�`hS��4�^}�h�]$O�6�����vIl�+�pH��������NpnԿ�3/�oH}��k&��=��������X���y���|��"�	u��� ��G�N�84>b��8&����o���o�|���F/kHڰ�K�X�_b�A��B��>�v#]���S_3+�ݟ{c�[X.�O�y��q�aX�JZ�6Gцd�Y|Ě�w}c៰6���㟮F͋&��ai3��`�U�4�+0��?Tܠ-��s�Up|m8�����g�&������$��n��+^��DQ�n͗�zp�����l�p��Uŀt��z�pS�Na��W/l��x�����/�	+��Y�/�(�hp������0�^�&BVB�a#���R�0��*�A���o��H��~� ��9��k0�<P	�:�DGa�,nA�́qUȎS�}���~�q~��^�uG�A������j�`�j/zx�Y��-���[��m8�ea<@�IV��="��z�� {�)�J�d��5��fN�"�}NgA�l2 "��c���Vp�[q��3E���O�'�6q�.��G�/z���K�eU������Qf�,�Ӗ��쭳%ɢ
N�?�ۘ��ׇ�W���r��㓩��(S�D�'/H��t(wOP�0 ����WT�9W!g��}�[���
��u$>�F�3��.eE��gA�����������I ��JqO�H[���R���R��J�ї@E�o<�$��<�r����J`�ґ�3�Q:�� ��O棶}jMÔ��-T������D_-���E�H��)��뀴��!��I���Q����ׁ��b�5�N&�M]B�P������Waަ��݀��}��o���>�xw�2�\�%}��Se�8�,*Q�|����8KJ�l��l�h�d���M
��gs�l��s���."�h�ռh�W]�mv���v�����] ��cڳ5\j���4��`.��p�@�Z���G��T���X4�*uǽ�N��V�)�5���؝&�7#��y��ZT���7D��N0�*��XS���5@P"�S`��T6NC��X���� H���,1R7�.�w3���MI7��v=v�F��67�a�>K���$6�/7�G�)��Q9����BA��h�+���q��u���9V�No��5a(��B
���XR�(}�H�D� � �2I%u����G�3�߆�,$e;7�x���^��l�_vp���_��Xp���r1LQ��S�x���I�����XcJq����ڷ�
�]��v�U8f��E���k�i��:�ꤴ$�'�>��D�dr.(�x������	t����~��Y�uBHR{}�t�Vi!^)M/�U|_��je�]��_����m2KX�8!��H�_�D5�٠�E��#��g�T��N6S�i��N�_��=QYR֖Fq�Ne��!�c聏�� ��F��Qu�����B3�<��O�3���:��N
M��4����"��5�������
��WM"���#��0Y����~^�>E�5�c�O�Ђ���b©��Gƫ�9݄��Xh1R/}4��.yl���"uY��U Y��d�th�?Y���GH}򍦋x�� Q!��(|�?��'�z�<9k')��[NB�͔
���P�)���v%���m�A�ՌX~�)�*J��iQ�yy
��j����Y�l���&t�1k����ؤT��� �`Cgc��|�CO�v/2:[�@����dr�3����������4�[}V�y��ۧY[w����ȳ�ý�6�e�n��x�SJ���U�h'"�q}�gJm�������I�F�q�p:�h/΋.�k��U�N�>�4I�ވ�?B���@��b�Z��A�^�Sz����.iҒ�р�3l�"�;Cܓ�;<.��OsW���_v�OB��Y�NE�B�L����6�M/;�V��i��X���ٌ��W�Ŏf�����$�aK�o��Lۙm)T��`�k�ᒯh� Ӈ�j.�j�Q�
<��P�5��g���6#ﲧ�V?�7���{�U�{��91�R��\�}��Nb�Pq-��jͣi?td*`n�3�E��#^��t�������� K^��|�����ֻV��i�b���r�vqEH�n��
�������C/�=�T}g����e����=�ҙ<f�B�9`E��3�;g#�����Î ����ѐ|�Q
d���1�� ����L��^��wV��?��e	r	mO����Elѳ0`Lʃi��MS�1��R�Lf��}6���hFO`v�qW�;G��Hj�Q��M��	�Fq�9w�w�g2У5��}���(�\i��7_ͷv�e�\�ktZ ���N*�5��U�l���&P�R0�e���H��z���|���I��@�=zm�FUK�|2�E�
 _,�1�Q�� ��Rhj {��A�r�Ts���D\� ��L	YJ���&t�������<ad�׵ׄW��`fm�
���ޠ�7�(Z��S�v���w���O��yC�xMB�z����Y*by]C�P����� ��3���B�����,�<�)�=lh��ξ��π��\ݰ|>w�E�o�,}m'Վ<tȅz��]\�Xlr�$g_v�aZ�� ��������?Sd�-jptק�������p7������-�d�<Maop�Fʛ�!��;ׁ獯�B;+ٲ�?�W�@�y�ޮ��A�ބp�:cB���ψ���±���%b7�ʹ�ʨU^�%�(%쟟 �Pu����rR��Z�#1K�r�I��#�y�W��+�o���r�sl�)X?w�X�J��~�Z�>���v����Gz>凂�J#�oT3�l����$,��2k0h{���Ħa�T�s��ބ	'�����L#�<���q{lQ�bY�g.Z<���i>�j:�z�h��W�o�TK֔���Ǘ�';Z������XL��)Ni�ø����#6�J뉚b�6�_W�_�T�M4��X��_�c�G6�v�(!�x�^後�����d��s��t��<�t��h9ȩa)�3ˀ�?��g�U�lM*�Ь��2*��$�c��4 ���%(�H9�lU����g� kiw�έק6�}���&��	�	�����J����C�j�:�Z��ò��-����^�a&T܂��'���xT"��m�=�py�ݧ7��[Al/���>ʼB9�a�1�E�����r^�<�n��$�n2��פּp$na��V����pX���U�FJh�N�C��;�C�"^���L(����PD���� �Ρ���-�>�(!4"�ԊW����>���U�u�1`-Z�5Q���Uߠ�	�������=��o]y?E\	C^��/c��zP�#^�ùj���n_VD5�u����xv�<�0�*�v=(���έ�>p�һ��l��J:������F�ht����6J�ɜ�,�Y��eVx�Q�[��Ϻ�L���A��r�|���$�a)�oR��	AZb���\}�m��y���-��iz����06�a�eUL�Nu��þo%�˷y�at� dxT��!*������#��Į�X%ϻ�h�]�Y��<V���A�5���o����))ۀ �슪�uf#3�XF	_�^;Q����#D���餷j'�S����S��^Y��N:������-d,�,�AN���|'ڴQ���C���3(rػ�e�J&���A�[s��k�M��+��kw�Q���A�1k^9)�7=�3<�!���z��f�f��M�X�����8x��鄵�����Z��!>�9��<������֍�٦�m��O�.m�ANm�,f����'��h�n����%�D*2������7���~c
R�h;�'.~(9ކZ�#4ׅ�?�h�9u�z+�R_ȧ"�:tU%s;P�CSXOa?����V,��fm�����~\��.��t�s�C1jm;di#	�6&Y����Z�Y5�>�Ks��ߌ�@��K��J	<�(��j����s{�.��mEI ;(&�b.�����4�3��G8!��������'��R���v�!�/'����G�p	p�ilJ���]��X�^]ѷKhf����;�{�&��4�������o�,`�5��l��u�;q��#H�チMSɯi�wy��|��v��S�w�	���x	��o??Gn�u�m�l���_����۽��P�V�g��$�;̠�`�p�&྆����8�M��~��=��X��G�ﲘ�?A�$iWxm�`�O�6q#x�<a�G�$<�T����j����>RF9r7~� `/�ɓ�	�\Y��K)�r;r���UF�UZ0|A��_[�3@R��t��`�M��.h�b;nl�\���~�h%��R�;"g�EC�^�,_�H��JFGٛ���=#Os\���Ӹr�P��/�F���ң#��kF�Y���G��6��|���6��?��+��#t.�M�;��]e����\�J���!�ֽ1���"���mƀ ������5�gT~�Cӝ0�p�՛~��$�\sf��j���E�b�!���u��I�q��)i��P�J�������q����hҠ��H�n�!rQ|��v�ܵ��[Fŀ�J#� �$�=X�"�|���x���r,�{�G��P�l]t�]��l�%jO�}<Y�z�\-M������$e,_�W�/5��J�=����N�B��M���,�N���
�]Z��5O�~_�i۠��}��Kp��#Р@GF}I��܊���=�de�.^`p��Ec�?ї
U����5�
n��J�"/fZ�oJ�^%.ô�?Zy��,jM�H�@�+�-/,��&��6z���mFiCנ�"}l�px��A�L�

��`TG1HI�;�?�S�C��=F�a2Q�Q�T�#��io��o2}��M}���^��tC� ���q�	v����<z�NƸ��9߉}��T�|���#�J�6x�Q�-x���@��:�Ō�j�*�!̽t%�7�>�N[�-P��=��i�I�G��b�� ���J�`�U&�I
0B��V��8[���0�	~��D�'���8�.bשF	� �[>��tpuI!p�O��̨�d�m8/�G�u��z��_�)�&n����>����a�lT��=/C4 �$VV�q��a/x����N恌�i�����e�>�5(�,Y�֧N��i��0�-p��P��l���$@b0�B8l��]��ٞ�4���g{ۜ��1�Ф���zX���U�o�.4���u��D�q�g�_�!s����jд��kPr�����14O�tu<t9.���c��8��2rk��@�jYkfR(��o6�$J `�f�z����AW(=�\�|Cb���zо�S���ۏ+���a�;���C@?(%js 3������N_��p��#�=J"!B�����|�>�/.�۵�rl�H��d��A6��,�P���e�TL�܌�^�j��?U˚�? m���X����N`��U��籉8��D���ؘq5o�Θ��
&���Ƽ�4�W���9�C�(?Þ�d�[f�y�Np���t�sV�g �F�WgS�+#�#�򆈎��΍�Xf�,�8SIU[H������n<_Rfe�1ز��hۅt$�
�0{!/(%�����}��R=Y�̙��ƉK�ܥ���*rR�s�:�i�"*UYL~���)�,�
/	����x����( �S(B��6$�|�:[R�H
Ff�3��TRa�=���)ޖ!Dfm8�hm{ڡ(I�ppҷ����AR�[>�L�	h��0䉜���!U]f	!F� �a��->�Q��G[�7��c���6�) =X+� "UM�8��)�-%;0�����K�l���'��\�~�� A�&B�у�cYMU��s|��?�(���n��q�*U;�x�	P( �	���_��щ��d;��Cot=?8@�aCT;T G1�gZ�a�����I٭d�Nu�y�'3>��l��\Wj_�~�8�E���$��QWɴ�}g  s)2?�?��"��d����z�VZ�;���:�) �]P&�[kx�2�m��,�q�{W֎f�i��oJ��F���GΞ��Q&�tN���DؿV0�T��&̈���F�jo�£)'�(����zX*xs�/��:L9}];4ڡ�l�+��,Z ¯�=�KR.E��X��,���d� ])Y��������%��Z%yƭM�J�� UƛW�������R�'_U*����G%W.��B�w���Қ!�(�Lc,�Hli9C�C�(~�FI�ѝ�����-1b��0��>M�YSsSv�gZ;�v���"��5�B��Q�ԪN�C�b���]�趙�J�������A�ڂ����I��c�� 8����]��s�Rc;xҽ�2�X�*-�IC�a��|r��0j��1d<�tuJX����H�
��B�rx����i�],J=��\���V�KJ5ȳB�0X�D�m�537��=��ʡO>���<ii�k�k�ޣ�B��3	��F��j�̯����#�����՜���$�UZ�|� �C�m�3@ӓ���і�$8�%�ʯ{B�T2�[����;N�yԂ]��Mv��VS݆����Uh�M8WWs?�EΌg�Vu�����9�S?_\׆��S��<������s���[� 8��m�7��E9N��ۚ�2:�e��jH�Q��Z����8�7�'}��,9�-o���`;|Qh_[��-�s�+,u�XO���o^��Jޜ�$F�ab����
��?��^�?x�����ֱ��m�:�D�wO���SZ�мf:��mW��6A!�5+f��w$���s���{:�B{�����7N.������Q��i����:�`(j�f]���T|5�&Fe�bKT���a�����yũ�������Y����_s'^�y�tb�:y8�~%MjAq���6�,�-G.c �2��XU��(��jU�Y?O���{����uF��s��N1{G�LQfjN�1N5!�>�>E��W�>gw��R��.��B��(�rC~/=��i()�	�Y	�s�k^�����k��骔w��Y9 5����`PPF�$��kt0G��/�F���A�w��Zq�#�,�ך	(��n1	4�#�y
R��]�j$&��X�
N�%��.�
�s~ׂ;d��!�Q����#�D�	w��|��u���3e [���v;�{�����\tT"^��Hhe��u��B�+&&���\<�G���O{����Z���ț�MݘM���ykL�^�.4�M	8n�z8J=g	w4�J��2� cU�~�{ޗ�`�8�b	 �ڿ2�{��M�2��l iP��e�SM(�x�^�T�p�B_.���)d@gʕƦ��Jr 1rZ����� a���q�%(��3 +D�D�+��h����r��D`�q���d���v="
r-mT����)��(дŊ,����>J�9GV�_�l?�J<7��A��u����y�MQ�~�1(�[)��ninn�
<$��{BO�Л���&@c���
(�o�c�-D�.i���� X�Tt�y9�=6�A){?����U���B��X�^sR�0�1o,%�v����:^��e�	>��@�΃\�KF�3?�>��l�\`J� =�=ը`_uc���aZ9������E�`I���/J�jN\P��A�5�{�]	(���;�bu���XS��q���X�%$�����5]	f��k��b*_�{�ex��bP)��EF�&�c5�4�~e�N�/�T�3^c�;ʸ�E����V��T��p�1V�;k*��G�t��Y1��+��8uR	��,q��x���,/�� ieF�ql���)�8���3(}ω�c���S�+���g2��f�P�H���-�|F��	��ϒL�~N��a����+� ]<\�N��L�o�Jԥ�VhJ�Ӻ#�~��U�k�l�[A���'0mW`��ߘyN�_9#4��\����#dsSY���Wd͐e�'�U�a����r$��۷JC>�t
�p���ǣ�����'y�	�H7F����i� 8�7;��ă���ټ���� �HgDq��3{4�_b�N��g�,����YC�f�U�p@2��\b������A#���M��O]�T��'}>��%��A��4��H i��b<��������3Fd�N��rs{��S-jp�w�����C(�2Y��g��'D<�r�~ 9+YJuL��)��g^A*9�mu*�$�ϸ !d�'�+찭6�U�$�N��l�>JP��H���ݭ˺9,&۔$�ySܸ-�Y����y*�F���s�2�"`�O�L�ʄJI��B^�6l�誦����;���kH:�8#�0�Y�3�H��9 TH��iw�p�!
 ��Q����
�d�8MHK�D�"b�%�{je<ux/ХH��n��!���b���_}}RV灐0�(k�Iw�d ԠM1�Ʋ�n���;Ũ2���)�rj�����9[��%wv�z��,lWnU��qxl�x/J��Y������dL���jgd���牝��� �۩B���.����.�A��S���׿�r�4|e�������f����K�Cl�0u�|d�P1Z�͢ʼ��T����|����VKl��e�6@�U��vW��k��RE9���.sޡ�s��'�ã��iAӂ�:�uGc�S��6$Y��{�/��f��g��F/˚$��gHw�dQ�<���&D�9Ŝ�)�����w�g��2�W��҆��us����55eI�Zn��J����D.�ڒ��HI
0���n���pY&�ٵ���{���#��ч��C:�BB�8O�|��n:���z<�}o>zaE+����Dm5�5���e�=�w��+-?��h��[^�iyR�nN+����J
\+O��P궞�^Rdɶ�|�7��X�[�,x�*�-!�:��%ۭEf�2Fۥx�4�aMaN�<v2!�.���1$�]6��Q|��}�wJ�>��x���d-2~նIJ&�B����_�s�h��M� �9�f9��󁚤޼�
���"n�xwPB����g��Q��9V��qA� ��A�$REw�b~t�Fٲ��K�j�%7Q��}bk�6�i����zK�䠦��Q��y�L���
>�$[��TK��9��eCPp��}��b�Y�i��[�`���b2�ob"�B#%q��l0Q����=�ʱ��|�hc�W2t�:.x�-7A�^��2���)~�Viee��^����s��G9��:<Y�_o�SJ��p�Y�������\(���*ѫD�-܌�{s"�%�B�V]T��2��wSY��/3{H���[�젓p;AbxȺ���i�����v�W�,��;Γ��e�1ؓ��[�F���%Q�u�+�!g�/A����~���c�
��&qf�¼T�|������eǵ�z}�)���HJ��r�	�;Ғ
T�m%"�-nDt��L"�J���ͥ��c�[Z	s�����w�#��֢�'䍟��<
�p�����Z_u����������F?��%#pk{&�T�Y�gp�_kt6h��o�_�O��j�V\G-*U#�,��Z����?�ei}� .�������9���xuH�"�N��C~<�&��ԋN8�,��R���%:���y�ݻ�g�Go�t�%�����p�w�j���:�NE���ԭ�V�/�n� �9��;m^������h��`�4%���6R �m3!�+�<��� �PdL)CVC��1�ҁ!��L�g��[$E�ZdKn�E���[�ϲm֧� 3w-T|&�M�U�v�ʸ�!D��:���L�l^k<��ӴW_��9&�z`�9l�J�\U�*����^l��é���lY�S%��G�*�Ithy%=��8��vgzz�F�g*��P~VF�栦��w�+SH��HQ���r����d�����2��rSn*{��F���Koԅ���N4(־�шG3�ߠ�Ҷ $�cJ�����[B"_���+h8��4Tt���*2��oA�������ɀrKD{AbC��� w|�J���@�;���r�A6��k?x���_�f
��/6^F�'�h���_.�#G���`Xk#��zi��Մ[���/#�  �	rT��)��+;�(��RH<�m�)v(|C�
;��S�AԜ�wQ�LsM���D�����cd�O�p�.Q,F���̌�����<q��r�+���45ݠ�����G@
��EM�U�KP��N��5<�f $�0��I��ǡJ���h-/�(S�>���M��!�f���W�Rn������2 �o��D.�4UA�`������)%�p�\���Z��U�A<����<R����ᴌUT�b���<pL$֨F$�1�^Рw8�U9j<�!jKє�7ZF�� 	��B�b/䵛���$��o[�fe��?⬂n8M�+ӀL�6�bD�zo����\*�K�fAޠ>�Jn���
&d�@ݐ,���������(�f�=�n��\#�S�jOM�*�G㔅���� �/5�K��\0�P��M>O��R�&�$�,w�j���e��e�H_%Lr@ ��a�]W�S��8�ֆj�"=�`�Zۉ���,<�o�!��w�֘-��H� �Z��1����-I������
��D�_�7F�:���X�9V�
�Z�l�O�\}/�*ʘp:gV(��m7l���m��*�GL4��
y,/WZ��m�Hߕ`ּ%s��7�4� ��[�,�K�S�����m�b[�m{| v���.��]ӄ�Eu ����j=�Jw����U�;{w�6S=��U$���L� 5��+��F���cׯ���f�
�ƀBo�a�����ߺ���~�i�d���x+
�)C��w	���I�����Q��#`�<aL}��xɌ�^��O�&ּ��]�զ�T,/ۺd�uB=��(�o=��?�O��%X#joj�s�!OF�*�S�����o7�Ι#툧@���?�6N-R��G���{��oz��i2,ֱ (����տ/�ys3�e>�������	�H��TݛSE7�'�ot�o%��@�O}���jmI{9Ƨ����ٔ�RX��}_n���(s�һ�hA���[���ZR!�� b�k΍��T`�r���sϊ>|"˂�l���:p���܀
F��+�Bkv����L`�G�en64Y�b�O��B�M��!뤢��s�;�K��| �Յ����|ܜ�c�p���=��d�c��W��{�{��n��ՖA@��ƪ����wK���SR��t���/�);-��_�;PO.p���VuWEĘ<��k"]sm���F
lF��DHH M7+O$�rv�僒��]�D�rE �&;ưC[X�&�r�=�^Yc�|ak�;��������?��bx���8N�G���5�r;s�w����pF������()��q�����gO �~UF3Rn� ���	 NDVP�5X���;�GJ8D�����u.��$��k�d�Lw��{�qaojK%(ͧP�]���0��;�5'8k��Hr�7�Qˁ����I�M׉W���A��eS��~w؂��bI���:Fcm�w$pe*p_�jg�y�鬳�pn�z� ۼ����k� KE��$�2m�<EGM���';�s ����j>㚠�b�}}�qָ.7~��y���G��f�2֌M��r�r��z'7D(l���s�V.�c6�n_N��;3�)�����Qt=m��e6	/��]뼊����g-����gB�ȴ�d�]��y�/""`�U�Wl�X�u���6e��l��uO�7o���]G�#�p��-b�DS�Ln��u��17!��O'$�j�is
NG2�qF��S0N��V���)"ʛa� ��k��e��"��8*�s�<(� �xz�5f3���~qnd/�PE��T���"g�^��	�P��T��v�n�l���<�oh���%uĠˆ�&�2Ox2#祲�(��I�7<>����L ���v�4�L�k�����U]���E�>Wa�-a淗3#��`n�)`O��WGEM�I1C���Ԍ�h�%,��b}C��65n�#d�W����u	b�oåk�d\��E^��j�紌�.J�jc�p�������QU�/1��xp����x!oGoi��pD�o�|6�G�Fcc,罬Gf��pT��QP�Z�V��s�'#'�ʢ���Fy�w�)��3#&��-$U�2�Q�(��{�_$����1��ۑ�A'(n��%�im[�� �����i�v�+��o� � #S��n���J	�dW�D!5A���\,(�����m��w�g�y�(C�:�d��O�/i�k끄D	ɦ4k��A^����]m�
`k��Jt�w�򭩠i��4�A�v�vi����z�[�m�ث+�<�j-��C�1�Dd3O�@����2�13w�@�$`Q׻7����"��jJ�BE���+�*��A����%��Fh�[lN�W���F}��g�2'�n�pK���S�h�����v-���,J�/[�m����h5�Mwd�>\�5g7񢍩��L�U��I'HmԘ:Sy>��8�
���K{g#x]�5��������u����t�`EPW+�2ܢMZX�Y�h݌s�Ǔ�d1���)��(h���R�&�Ѫ�m�b�#�P�_��.P:Y}˜�P��7q��r����$��Q&�PW#�V
�)-MY�;5}����f9O;p4);~g��}k��+|��?�ՠ�$�HZ�PV���8"�ί)�6	�3L;TO�6�ܱ��cD~J,��y����K4��f��u�0o�"���.�{a�6p���!�&��W�]����&���2ei�D�^��M1����^�Xu*i��h�W�!�9qV;�p�]9�<�KC�}��Y���ry켞rFZ`�y��(�+��9�.���Y���H��$�|<��3�iV�	J&�uB��a&�^�{vv�"��)w�>q0�-�b�v��,/l1e%��W��j�C��s{ur���=k�S�����83 �Z�&�5O�˸��"7�`���Q�^KD��襓�A _��HJ���K&�Z̚,6�sl�E�i� vP@OgY^l�[Y��\�w�wsd)�����z��T N�n>N�D#� {�`�7Ⱦ@Ӿ�V@s����k(җ+�C-���n�#J#�/�*` �/ݜTW2�� ���_�,�.��QV��㪳c���_�Y�[�����4.ԋ��=�@%C�X񖖓�i���M��ƧG�<�_Lh ����_����kИ�h�P�Pٺ���\��F��`��g_u9�_msD}��vM^b5�V�-9���Me	@K��u���I
��JT��V��X&����ި�_5��"�;��qN��\2��F��V�N��<�V��0�F��}�^���,��H�s܃h���L���B��G�e�!U����OR���c#�{D(��[��xH�u�O��;���{JT��e.�@��4����	vt����`>�Xv�Pdu�V����� J1��0��u@��)� ���]�}��J�㷛���z�oy�.z6���ZL�0}&�%7�Q�N/��O������v,?@�v�&/ಶ�Q����xߦ�`������c��I1��/KH���n��(�����Kː���d�M�q��9�V5:d|J<`�H�F#[E�*j���P7��d���[����lUy���O�g,g���w8w{v�&Z�󾪥Y)Du�v�&ps�4n�v�f�P7ƕ��L����4�iץ6�T�EgZAϹ�7����=1���ĚP�v)�R����4��j�,�9oh��wPʼ�_�P��]@��Ro�ǭ��Z��� f)���t�_�wʹ�bc|�
i��[� �S�5��^0�1��Jp����f��4쥺L{{�n�����O�~8� >K�#�����fx�g�\7����m����p-��i�1y?�᢮ �-H#C��+��)��)�8-n|{@C%���aV�n"�;&5ZK�
v�W�xY�<�[�<��Cm��s���:�W��\�L�e�Ո]�.���0�sg�qv`,�;���%�
)�_b�K�"���/���}5ط�XZk�w������$ 4\���	�,�[��]�>XtYա���Q�� �e�^��7�[i�s tP��������p.X�����}�L�g�l�`��OPD+��V�\�~G��Z=�B�Q4ܪFV�������?�W
�&/ZI�����qs�Y ����z:,Uʢ�AM �Pr��*
������*��vT�->aЛ�/�(v�Dc L9(s9���Ku5��^�6�� 9۲ݣ��T��~��R"?���(͍QQ[QxRŴ��bp;��F*TW&��r�]�`I��hPG�(D�r%4��:�4�|�޼fc�{ᩬ~����w�(��S�f�C�	)`�#3)�uvʁ龷�.vV�9�sve�?{CL@���(�kJ^�����.�kz�v��f��(q����9Qg��������oh����iL>�}��N��5��Wq<�������9��)�d�0�7�+#���\>N�
L57K�GB=�G�"�5�C0�2a�� [:?���62������JVY�&2�!�6SB�J�G�qk�Y�Yr@8iq<����pÖ��{���8�hA�G��f��8���kgt���VĲܫYqn~�Y��+4O�X-kD��w2�Ϻ��b���D/��_^�</i[��U���g/�5qǉX��1E�fcj�ļ�5�Cb�,�	Mb]p�
����
�
���7��n��kUU1��Cöb;"���qAk�����n�L�In�ǅ�-�W�H~,����h�3i�99�o���<Y��7�;ک�R�N��ǫw�¡�jr�q/O�K/J��ߛ�Am6��Q3�u������]�
���p��]ۺN���e�}��3V $� ���ҙ�'�r��(��:"����ge�ސ�,ʝ�%���+�V���?���ZyE��� /�{� ^0.���� �P�G�LNj���Y^�ܰ�K�RG��Vfg��OJ��K�1��G��pܺ���fN�g�UD0�b�2�A��7Jf_�������T�"E���/ ��fp�K{}�3���T�4�c���+a�߾��r*ې��l��Z�?���Xd��2P�����Ȉ���Mq&=�{�����3l�]3��\﬚4�-�W6�GB�p�7e-�68�����uPR ��l�pBV۝l�߾�JӑW}����D	 ��%_��"2���PP�W����Too)��;{o{��Y� t#��h��gQ�{i4�wB��A/��\+$�����;P=�J��`F�4��]ǫJ�7pa�r2�)[mT��P@ �)�KE3���}�`C�q&�9-���Dc�H�����q���sGŠlU*������#�Ŀ#���k���23`�тR�:m)���wz����8�q�V�E,N�������s���0������C�P�T���.h�:
�ʦu��`���FT�j"I,�� c��!�+�hL�J���oa*�n������<�[�f^gq� ��� �Y���
eV��e���=���C�7���5�,�pS�2�@�&���s��y3����4�%� ^=�N���Ī�Is�3%��4��2<���f���:XO�'��X61	�8O��p�j�"K�t�eD[�����:��U@W��P���g�A��x�f U��B��&�n�}�����H사(�{�Z��;�n�9cEk��6���ZU�t��j��w��=�_�Qd&��O%��*Z��`�(��=Iѩ>�ҰǬ|?�M�F��T�7%�+|��V	���f��G�2�����?�sS��C?\�+�PA������n5���"]Ҳ�Iv���G���&y]y��܂�'���l�q�s��� �i��pR�:m����z��V9zrؽY�S��G�#���&�D:�Og.�����
�Lŷ�&�e�pO{9Y>�~�SaX�ô4�z�׾&��V�!��]I�����J��d���}0��f�}u�P�q�jn����m�4�K����?�*�xհ<�MQj�67*J@�3?ɫ�4��pH�a{�Y�wWWL����@yvr��lv;�yy�b�J/�s̿�Ǳ�VH����)�i�qZw�9Nep߼\�E���7�)�t�#��Ou }�8@� �W��)I�gc�e���.��v �j�R��w�����v8#1fL)��vTŇ{u�b���4�R�@�ht������U3-�<�wiv�p�GB�Z	U�/#D�k�<D���%x�cpH>	�f��:�%��J-��,���(8X�q�b�$�~
� ���?FHX��)���T �ERG���!�p���������[�+�����,RfZ7��q=$+Oh��d,|z*��0S�J���lB!q1����}9z!��(]R0j
gݞړ�&�����
�g5�e\�p��^�E"!�.	Q@�m>]����{g\?IT��p��vuN�oK�GH��Piuv��#v/�Q�WI�p!��E�ֵ ua�������J�/oI�Wv0�\ZF'H����/.	����`ѭ�3#�>��t��Ə�ĩ
89�|LHj�TC�ǜ&� +��a�Ƀ�Nǈqa;7�^�㰃�:�h�`��ړ����^Y��eƌ��	�=��ÈB_���ɀ��
&��R�R+��z)R!* D,h�}6�d���I�@PYtke��}?@{ߚr�-�jE.+ O���W*�B����S�r�8����'V~��č!02pF[�f�<l�>� ���ysط��eЁ��i�A�ōӾeO�sg�?ʯ�a5�~���9.�M� ��w���F��_Z
�u3���>�Բ@z����������1�5�ut�>��O��n�q1�;=
���?�WD�r�J�i>MI~���WW��2I&�� �T�ޛ����Q7�d1���).{5$w)�f��F��'��'s�C�2m�nnKs�LW���=�q�F�B�Vp��@��*40��(�Ў��q����/}6�7%os��`�&����2�Km��˺�4����Z�x����#4+�2G���9SB���Ȋ�#�zrP��̲�;$)\�gg����e�M�������ҧͅC�I�Ơ63{lAsI:M�2C3�b�Wp7���O�G	P��i��S�̄E�#���Tv�*����1i�2�Be���0��R�Q��_�*4�ˈ���������4o��ĳD��v^��W/�=���y���wcĠ�������E��3�d�N�dt)<�O[��u�n��N��g"�E�;?X�;l�o�d������EO//E�$��w��$��7�.�?�	oE�{��k
˓���-|c���	�_ۧB �|�o}��sS������N���̵�v�E���ԃ�K��=�����<,ޚ1�Fƚ֪`nyt��>�໮)��;_�{�7IM�*�y�:d�DE��D����	�V{B{��5��:�����R���=ʻzr]	����,����q�BH����ѧ�Q��c}�twX�v�})`طa(0����"���j�g�~3�GKy/]>@m`��p�8%�`w:\ �"�fe:��U�S�
�o���{OB���4Y_ȓ����b��q�ŋu�9�����W("x���ȇv�U�/��x@����t���*6��%w��ߐ�*��SF�B��D��`G��<�_��v�J4�?q6�����̙�g���z�}xsx�?��WT�g���M:�+��D���R���e6)��øVԲ�eTp+#����6@��䗌r��:2a�����X|��Zv �F���f��]r�li���
���'�k�ֲ��j>��cq�VEk���0�<��A��!�f�"��*%�?�]=����1�э��׊�'�Ό�4�lG��/WXf���C����FH��y��(喁�I�D��
�`�s'}"\3�ֽ��{�_�C��"��P[ʊ�n�-.o����B�[��p�6���℉kG*Λ)"l�M���i������1��x�ˏ�|b�'����4F��R�j*�w��Ò��>ד����%0�v��(dGј��?�̳��ܞ��0x��Ni���̦��%��Mh��
�Q�d�h$cSj�9j���_`��-g���`2u�� ������"����$��z�2��{��D���ؤش�^έ�#8��if�����5�B�;�Is �A�%���G8n�� �ey�E�R�j�d���>��x��F��;X��ר���GP��T�_�V���Q4. �~���l�ީG�ے����'ǥ�ٮ`�'
^�u��IFn�h����6�S6RE��6a�ú�uZ�؉��oJ�n��&����d��Ռ��	F�3:Z���uXs�/wוL���6�h�y; �aN̤l��#��'�����Ũ`���Z�!�����R�D
���T��o�x���"Y���@��}�LL�^�7���UD��i�sat�ik�Rs�ݫ(�������b��.h�D���"p\m�!޻s6��2L�i��-R
%BA%*�3?���f�|�.��1�kc-��_i����E�<qn�p�Y+@���4�c�qE@nE��ߝ��g�N�4~�|�DoBx %M�f'�'�[K3z?�p�VaŊ��F�V
��B������}tIQ�l>�Iw�P�������ԑ�//��$�"o��]��P&��h(�������� �{c�g���j������X������+���>���V>�.R�T#x�������ވC���#-�Lo���d������qzA�O�?cs�j����. Z���i�s��&u5j'D���<$�]�Ғ�T�vfw_U�4��@j���wOv�ak-���Lw~ �J�����4�t��\R/�_)�	��4�ӧ�=c��h�ѱR�x�.6z���Gό�>�$��?A������F�]E[�8�£�z��y����¿N����x��r����GP�`d�������i�I�i�EE�L-�MG�1���s�|Lzũv ��4��"�<T� #���?_�g����	�آ��}}o�h%D.
1t�>�L>�Z��N�LS��i��ƪX�d��%��?~� ]���B<�FR�ڢS�r��������+������u��1��Y.�0gzƟ����S�G ��z�Q52�����Z���!�d���X�<|�u���[��͑�
�8/"j�3}*U<�Ϸj;����0�X��ؤ���W�m�+j�ĭP�*��4 9f�6�A���nr
�H�O��h[��;�}$���� N(\b)�1t���D��n���c�u�/����=�s�r�
s���5����l��Qc�3B����b����l�_���Θ����"�f�
����g �8ldnC���Eu������騫l.V3�9���1Z+3���5�4o��lr2��v���x߼r�ޝ�E�S�*x����>��X���po$�*ނ�n�RD8���q�pQ�I�.D���Z3���.\�_ّri�TA�h��T�`𷯨6�y�j&�	ٝ	���.��.�X��,�\6;�U1���8�XHt�l}��R�!8p ]4��몆Z��ێ �J���Am[����w��]���S'�(�y�"#sUM�mst daj��������6���E���:���p4�����)[����Tɝ]�j���F"`�ۢ����O2��em��މRHs�pX�xG�4��S�aV"m��e	���Q��bo[�0�֍��apy�ra�ǚ�)�[?�y��ۜ�;�E�@ǃ�R���`����E�z� ����_���Q��3����ؽ6g��=_��Tr����F �\cM�*�]�-���ɓ5G��Pc$Ͱ^km� �ZQ�<�A��EPM�K�p��q���v,�Q\�Y!1��Z&�Br��L��ʪ��ʉZ�)�� �G+N�bn�x4m���i=�����l���^S�vE
����~>�=���5�N�����d�p�����K��4d�'�1�āܶT�=�X�%���P�oGSj�ӲC�ӓ�hS,�{�W_d<��[����4���0Y4��X�IW#q3M#�ٳ�
�h�N,�9���h�v���s�Ү���SΜؽ��[
�W���#�-ސ'�yU9=�5����#���|q a�ߢ�ǽ%���/�{�����Xg�G��H����%>K�]_Ŭ�D��H\���K�(g�&��|9K��.I�-5��@O�	w�:�ף���q�V��P������ނ��} �vj/,��l}@����x�:����;�/�����+�*%S��	NL�BM�V��/%T�P����/)ru���YD���U�JA�=5��xɺr ���:r�4�_,�VP�:�`���i�8�ȋ7���v�.�<�q��������@��\�3��t��I��[��[�j��J�U�Ȣ	�\�B	�����HD��,c��~���MоԅJ�O�ߎ���Jt�:��G4"!���x��ܼC�-�wӦd��$���I%���f�x�#���}6���e��I��`�<m�^�N�2�E���p`D������M!��)^YV'��<���sӰ�'p
���?�e q��4�������&��m��=�����j4JYg�����S���W[J*���Z����z${�
x�T4ӳ�_w�9��ϓ�()�}	3��SA/��üZ\�GCN���Xk��F$���6D'd�7Nq������F����2��+q�t�]���>�7A�IW��J?G�%�T�R�z�@��#���6����A��q���E'x�Qjs��R�M:�ڭg�ca8�mk�D��,�t�ǞG�kD��_D��u╘x����X<�kG��(���'�����
)c�g,[)Du�L.������l6~Wp�o)�"=��j�R��C��2�([�w����F�A�}��{I�'yj��מ=�[�9���P=N��x������L��]@p!(��`�y&�����SB�=e�ix������$N�Jz�§"t6��ՠs����/�����vV^�� D[�b��>�.�4g�B����Bv�l�L��O���(�9;��G���5�ϰ���`��k�X�s�y~Q��d�8Ƞ��*d8�s��^x� S�E�R�����EXyC�a�a�}����;:��. ���3��+�p����w���jf�Q�ۨNJ�
%��/#��Y��.���A����T�!U2��옄��,b�5@��S���IaݝܮsW�B�|l�`3�O�lT+�* OS�j��Ue���"Sev�����h���Ѷ�+#h� ��.���2�[�Q��J�l!h�.�ӷ�yhN}�n�[<L1/?��P�ӽ�N��:Q��0��=W�ι����|ą��MV#�(<u��CXi��Լ+ş���5&@�cUU>t�ؿ�1�	�7��M~k�����;EV��rЛ��%{R������Fs37���5�c�B9iƍ�����ԑ�A ��%L�JVl̹]o��I�'C���V���}��;�ihP�'�]#��C��"k�i���D�i��n�;aZZZg�f=�y(�~�S�,q�r1�#�)��9���❮����-��٧r�@F7�p�*�H�L�E���W]����"�9��)M�c
�ʊq�z�UʯZ�,�u֋�VZ�[������P�Pag��o���}��6���{�5E��Lx���m�6��k`d�P���k�9��h�g'o}VJ��e��ǣJ�2�-�isך�T釣
��::Ӻ#�i���Ħa��yl�B��/������7���N��->Zε�(
B�z�f���; W�D����$M���7;B�S'�dp��H����� B�t|�~[�yEJn���1�)��M���I0�>�Ũ4�9�eiexcz��+�����	���7�?@���[��\P�}`���7XD��L+WA~z+��������>F��b>��V��X��Ki܃=��}u_�4p�o����C�%!؈�!�C׹��5�O���V�l�;�����Qũ�St��ȑ�:��\6aE�d}�h9^���d��e&ح���c�ە�[��$<��j���3�[Ֆ`�.�8��T�<����]�@���]�G�?M�i���~)/|������}v+��r?<\э%��TI��fY���s�cCꋘ=��M�'���ﱺD?��"���s���q�͏��Oʓ��[����"�Zv�S��պd�Z�l��-
��R&B$R�^"���5����c@-��[���SA�!�u5(�#�`%c�zr._JĞP&�&w��]�5�Hĩ#dvt$	�WG��G��D��p O�m��tpO���5�v#�q��Ma�$o�rS���<��iO6O�7�i��9�P�XQo(����ߍ �E�v7Tz_~����/H���)�bD%��^�:U/Pt���b-C����	Sy
3=���8��S$.�ǁ�0��P���cDen
�b��r�|����x��f���䯰~��ʿHM)�V��1�P�=��d2��r*�Qń�B<�0��|:d�O�/9¿s2=�,����'��f��X�#�H��n9��sX�u�".ل�u��$#m���o��+���D޸�$]U�A����eaB^;,�2f�����Hՠ�i�R�ͮgQ�"�����b���j�2�U�Z����R�8�N�H���V,ck�l��������WE3����`���gb����|nz�|�z"��w�K���(�.H�JK�7����1%C�O��<��Ʊ�>J�!`����B9�UՔ��@�7;0�Qݞ�/O�:XJ�F^b�9�����+����EնH˧�-$���F�,&5���k�������0��$g4�����!=�}a{��:�	��e!��!w��HS�ZV�4��+ԯ�'p�!\R�="Q�?�������@�\��j�*읏�{{^�Ǎ��]��%��z��.��J�Op�z��CʉSPU�4�t�K)i���޺<�������l1�W���:���`�5g�\A����'��CIK<T�o'�o� �G�>O�ms� ��w�q���V�8{�i^E>!�w����
	Y�D�"���7�-+t�q�6�3|ů7ݎ�yM�r���i�ub����BLN�zM��$vޕ�!1E�ndn@�m-<^,q��8��q�Y�z>[��؄Mvm�R�I|-��L��W�O�}OߍN������>~�K�2�nH:�TfE�S�]����M�(3w-W;�ǁ���8��6O Yp;�,��g��<$��d�%�<1v��>��]!�kP ��;��t�`�2l�;&Q����lgr��iGw�T����� ������>�h���Yfi�����,�~�&gv\�vT� Ŧ~-'c�^b�)��炠�{c����GI�c����P�Aq�/��'��TyZ���|L]E ���G�6q����i���0$Oym�W����]��/�01چ�Fk�h,=Ea)�ٯc�bm�8����S]���
�속p�f ���Ւܠ��6U9<~t�c_rWO����Ӽ@�b���$k�!���^|��e����I���G�8<"	[�.ݍ𢿐�R��L@Hj�Co$��S�ڛb��!�h�:�8��m����ʷ���C���Aq�ù��_L���&�!��kW�v���Zf��ܼI��n��nN˖���@d��5�#JΎa��1�J6/S��U�������Nw��A��h�i�c�6�|P@��W��;|�� c�Tx�K�W�JE�)�6�@�Ҹf��f2d�I�2)9���>M|1����h�6�_.����f�4�����#S�j70��&��$��n�:+�w�<W�[�w�[�d����QH!�ZG]b �y�#�%_+Ӊ� ���G�J����vE���_�JL��Dg��Ň��#�5Fr�!B͕���M�Ѵ���f����Lwk5ګ�{a��5�>i�Nyש�vP�Ii�Đ?� R���;%�=8�)�p�6���3[[G���ʤ���2����@$h�j8�4dB����rY��Al������^'�O��pv23�+E �O%w�BF �k���.̍-�0�0�F��i�8T���p��Q#�o�
���\�М�:��9V1 �@˦���F��cv��Nr������W���7��͵Hˢ��*�2���:�v���hjט2�"E����&J� �'
��O�zm�'�V����� ܟ���5^�y7л��? �j͌s�@�c�9�)h�O��!��obe��Pb����y��Bh��0�︌�"u|ŵT�IS�-@ 	o*���'횜��|#�*Z�����T�������xV ��s�e�	'd�́�Wx�-�N |/Ox��/pS.	G��a�p�bC��(>u�����\�#�l��_����p[�_6��Bwټ�
��ژ�9�R����K1��E�^�7n�c5-��)a_ B,���Vک�FVX�����#�PΤ��Y�L�����Py�RP��5YYd��E.�/���`��?e:��:�i�t���R��Ʊ�m��43��u�.ٔ"}���?��T���~��������9���>�z��y��D8�*vI�_US�q8�!.�BZ�?�b�]��޵N��}4���:��޾<��g '[A�z}��4�J�Ƈ�W��å��
�Ѹ�����rQ�B�VoAP۴.� ��1g��L�z[a�O,]#�K��j��SN=�ps晅O��B��''8���<\,����)8���䏲p�9z&��]F�H �-ݟ��j?w�em��X��F�^ߜL�Ψd�%��ޘZ
v���\bL+�_ �[n�'g���9�Y܎��F(K�|�!�o���� �P�eDwȂw���d!+�A��7<\o���m��b����I/P�yBF�5}ɻ0�D���iqz�cU�(��h��(P�DV�D	�򄐋{�Je��R)�����74?D�u��� ��]�������ڿt�!�Eb����2G��$�Z]4Nފ�r2�2�1#��^�$
�� ����;����$R���;kVGڢz�¯�@�R�Krn�����#�򸠿y��)��v�c�3��Jg>�x���t�)j8_6R]Β
ygi��`��,���s�`z��9�L�/�3K��h^C�鹊�!g��c]��t��a 3�6�L�2"���[ e�\8K0n3m�oN���4�8�R�"v�2O�!�f:��I�n�E�q,gb�7:�X�H�r�:�ѩ���b����p��݈8��]��+/.�ﮕ[�4+:��A'������FI�W�$��_�׭zN�����Ѧ@�ɑ^� 7���f��y��a��}��t�(�>s6����>�+_�k��h5�LÑ���.�c�dm���Z.N�"8�U�֝Ζ��}�1ʂ{��q:�[�A���*��V�q����|
��k��J*�wۻP�L'ə��xo����R��
<'+�Lc&�Y)r�kVR������{UM��=�[Ϫ@҂���\�����a�#�`j�Bx�<AA�?&��L��,N�`��C��Z�
N�Ȑ�m	���W�5��?��y�Qp����Bj�/�5���%@ɥ�Ir�^}Z����.�ļ���h?��0py����K��T��o�F��E"ҙ���g���E�n�\���DB��Of�}�I�!��4�EE���~�a#�.�4��Ze2h��J4�	m^�LAv�uy�����c�).*�s�b�C���(�m˝C;Xu��@���Rі���am,<T.�:�9-���vɹ\xĐ�\a���\��&�;�/��c	h(�W����U2���3��8z�a��?�t�A�i��'�� �獊�Z[Q�SW?�Z��P�X-�g��M�C�^����������J����7���ܞ`�VL',��Y#S���/D����e�˷��8H��z�~���
~ ��'�Ȋ�Jdc���������R��-U���r�D��S�1�����	bZ=\ �7�H#����_q��!��Y�n����	�ؽ.������[,���U�`E���B�𣶕�m�Z>�d�p�`�n}��.�	oj����<o�{0�̆�J4x�� �son�'aɒj�F����S$�4[n�������X��	9�p�BR\e�H��g���m�]0#=mi�HM��]��$�N�}%��[�V�i��3v�`顤w�Z�R��٥J�I5j�|={7Ϳ��ѝw��w�v\�'r��$����~�l��@vVRu��0 �NG!�ny*UР�f�lb�.f�
[���ty�S���<Ȩo�#_�&~�<�B�'�",�X�r��m\4��Б���&+yH@�|��RZ�8�M���$>�5�B�W@õ&U�)�j�:�V���b��c�02?�}��e�u��>�^)�9�鱷)M{0k���I,��p��L/wP.�b���Ը�0+3i�V�K;�¾O��f��|Q�c��L�/y�Q&F�%Y��>ml�t*4F9����(��!�Ǳi?�߅�p'�����TKi�M��Į��[�����h���hlg��z��}��^I���ި׾1c���ь��cݩ$��y']{đ?��U�WE<y2�oqd�B���{��L���/Bu��#�	�R��M@I�����낟�8*d��1�z��f�v��$,y��΍}Cq�̾P���8λb��@�:uR:��J���.'��T�����w^���À�*?�.@�\Tƪ��s;���qy2���7Ym��N�r����Qg@ҹ7����U��3���"^r?��qWܽ�O�&��-��ޑ�+(%�?~����S���	I}�����T��H���t�홳| �q ���*3k�Nh�w9�/���l���L�=�PV��6l��G�eǆV�G������̎K1�y���8`�e���&��8rz]Ad*x�\�c�}*�����P�(�Up]�� ��	X;Cx�V�iY��*�V�� ��h�8�8'3����QR�y��.��4�7P��v��/���b4ɑ���~
�O:n�hߛ������o�Hk�3�Tį��C'y��r�酕��UE!Fs��cVڳ��?]Y��ԧ���P�$���xQ��$m��\6��/���4Y��"��C[��Ј�{�y�bcxSA*�p��x�?ԣ��,OC$T"4��)�7:c����2zq�;<�;�� )�bᾁ�,�uW��I�N��$��P�сD�gtȋ�;0>[�yQ�迺�k�#�����;���kXǣ�A�ޠ������L��?#���L���+�5����م�p����e�D��E��/�[$V��&�����}�_�=�UQ�ZT��y����*�X�g�z,1;��T)�\�W���m"f���0�,#�1T{FƉ]$�3>�;������TyBAQ�ahy	��	�%-����d15)���|[_��"h��e�W�e���=�$�ZM�f�]�
��;<��(���w�6�`�2)���N�Y�,��vf������刡2�l�I��ȅQ��Q.Z ��	Nv��l-zv��FH;�ؕ�RR����"x�kGk�/z�}�J�݇[>a
������:B�Eq�3�Ϧ��ztv���Lg����Rz�J,��.!��G���GT
a�M�3Vz�P�:����OnρW�g�,'z ����	�𦘡��J.뵍���au�~+�TBʑ�?&������a/�+)���c��("��6j�f�Μ��:kj���J
]r�ȼRm3�Y*�qI�O~!����P%⻈O�;�b`�P:i�}��4��������p�k,K���8��vZ%<�?J�~����|�{��k`*�O&O��,Ώ�+��E�uV�c_CE�nZ��XZ���^���4D�,�%��sTsb3�b��T��Dl���d�S� �Sd����Y�g_��d�.���K��s0���vū�Z�w��q�Q	4�����"���=�0�[�9���~F�dִ�{��iW" ߯1ѕ�UK�吴�=7���B�y��C ]Z��eN 3 p�RA�^��w	/����}�ڮ_�O��rc��I� ��?L{�#��m�dw8�W@.4�ό�zn�_��\�~qC���`o�֜��<��?�/6�ҳ�#
İ��[e���E��*���q�EK���W�J#B�c�{I�>ikg�|��|`���X��;`%W)RG��pv|��g��mT��lc#:3�ou���Ü�����G��Weu(`��m�g��oW"<~J];��
���Ȅj���>��^q:M�V�2D65ŷٻL'���xPt��]JbI:@Yٛ�2����t��D #���������������;���sm7��^��>�I�j�a��uw��5�[E���aҤ����_&�`y2Jz�j��i�����w�XOYo�H!��?�X�3�P1`T�+��_�S��R$kG��>�.�^���b���y uh#Ԁ�:����n^B�3����_`��i�.�Uԥo�:Y;�I8z�A�s��MZ�l��I����'�c�_=�`���i�bǕ���cu��n��Ê��71��+�<��5��r�3]Ϲ��f���2��x7���>7g,�*��vw���( Z�=���8~��
i��GQ )0P8()B"H�S!>���
���A�0!�eW�u~t����eY]^��#�q7�P=���wy7�{c`�0�k� ��Y}Ju�h�γ����C,zwaz�j������<���U�^��F���W!�pܫ�\�	o1�m�6�(b/�����ʡUrXi�g6����/��%�z���T�Ho^l����hK:�;^6�=���+�P��\k��	�J_AQ_?���u��H�ז�8��5u���)���ҋYB�8K���9M�٤��wB�4�!�Ġ"�c2�Em�4�%�+��`8���r��gR�m:�-��c��~SkX��/�SW��dT����4b������ݺ����������ӕ����q�K�ߢ2�v��m� ���ǫq�*��ᕳ	��a ������D��o���He�r�ۖ^oG�`�Ƴ��r]��*u�`"�7����XǛ�@��ͻ4�>���mD�����R%�����'�LDD}^���Lf+�Ԧ:J�k`��
���;��jiB�{8W?�ƝZ�K�� 
k��U�O�z����̑j\,�U����}(�l�5(S��a*����T�P�4mr�+\+�uu����0��_�cׇ�a���!ܧ�+�J����W���BGVksh|22��z�\��)z��OI�@��ٵ�M������6Y�I�x�r�u�&�h��QB�ٸ"�B�%���̨jꔪq����Ms�i��WM��6@�]b������N���v@�0]~�r��������j.ȶ{����P��l���}��$������j���;�*���%ql�!�=6j�����P�O9�Y;ڃq&,��e�Yp��r�S>;G�C=�\X(�x(��O��C�T�P����)������"ɉ��>��:?��Ď���1��){�hT�$w�����I1�'��-C��`%�ߣ��n�>���Ʈy�`���t�m1@��v2�H���>��B�
�;��?����{�P�R���-{�t�7.�3�]��'"��*L�P���Vq+,ɀcIIM�1j�pj�Y^�+�z DĠ������җ*8�XK8��2dx�Ԅ���UuJ>��6�6��9����⓾�c�w�!=��l��9�f4����2Ǎ4g���8o��Z"�N.W!����t��b���P����-�]5��- ��nW�f<6�"�S$����u?�%60����	mF��������'�h {��ă	�
�����Ը1��ͮ���;ӑd��:^�+ł��v'o�%WC���
k�<�u��n��Z_=]"����"[�g\�M~�oo���2d���	�H{Iԫ�\�1������plZ�o���9�ĥ~���9��4���b׎�0>-�i�bp�>�H��+H�]~���q�2�����pxM�4R�@j�8�Օ�W�D0g���yDA��%�����Z٫̞�*����������B_l�f��9�\QiF&����o߄#O�=�B��F����@yn�2��QU$������?S>>+Û��
b�O���,Z���ETu�y�Կ�3*�+<�1�6�5�|�ݎ���-u��QK��1��T�.7K�#��S��׏>6�x1W+���
>L-��o�󂓠_RO��6�L!;��'h*R��*�8%�[����*,�ユ���T]P!���1�L0�ſ�N�����pb� ׯ)��15��C���Q`�M�g�<KϘp�Ya���ccf\+*D�������8��7pL�?�ۣ����:m�y_/�;�'�&�Wh� �2��d;&Ў�}=���]Ը�*����3�t�)��r���J4�e���_���cy �۱o�W�NV.�=9�ӌ�������4�S��_�gC���fT]�?� �>�̜��2�����q�ׯ>�Վ���`��a�����2DSv:��tf��>,@�� ���o�����5z ^��кB�a�t�"+ˢ�4DSZ�5}��\H>��""�S>��7��
��\g
��Ҝ���*���u0���PZr)��:�TuW�Ԉ���=��K��w����e�{�Ke�ߡ@��m
~���}��Y���X��9���h��W�.����D��"֫���W��pӠF���Sx>۸�t�7L��Qf��O���ٴ�OzO	��u� ��{��*���BN�����~�{ٕE���Q̻`h	��dX-"�V������#�ƫ�	=��D�-K�w(/bZ�
L�Z�v�Au�����*Nl����` ����z-�Z�R�M"�I!j\W#[q1s�bO����\�|Oe����;6E]�������4M^�#��\-��tys��2l�߅���}p�#��j��R"�*?�ESQ7�����-�7X��Go��ߪ��c9�����+}����|���ޝ�0�G�r�Q�i�'g�=�GM����te���C�i��gvX�bc?��)s4A9�% �w��P0�z�՞j�������} wgٗq�����@-�E�Uf�KO*d�P
�ye�ݬ�l@c#���Xq��^9���i&�E��8�����vv�Њ�w�S4�[��EVj��eU�S�AN��i�h2ý��͇��%�6�np9p�R.�<49�x�f�[��3�#k.x0�o����CF�5\�wX��y��n�Ty�I�JhƉ��/��҅��M0��)�ӖfbH	# d�ӓП{��[m����^5����<ӤY��/�4��k�1Yjl�q5���U�m�H���Tu���Y��p��Y_����=��`ԳP���ǒ�GM5�H�I�n�4�}UX���WU�	�s���Vr���~K{(�z<�M�S�Ŀ��_�B]���CA�@�>_VQϯ�A��W�,].��G�;qa>���>��>� �G�1�{��)O��bt�"��Kޘ�L,ߕ�3��h�i�fWpNGN��G���r�l�"����r�o��B+�"���d���{�	��q�����#��&g�췘������poӜ@0�A�6N$N]R<H*m�q�I��cN/���eV,����$u˸h4���h[��d,7f��hM>n����b	Qm<�ġB@ґ�+�g0#p�H�8Y5�jy߁6��{��<������PXlG�����P����G,�Uػ�m:��H��M�Q��`Ht��b���/�SL�c��:U>��I����56�:3!��G��Hw��|5���k7�Ø������S[m�$h�5��=T�٢YO[��4��F2	�����xe��'�G+λMS�����+Қ'�r7��LB�nN��I9C���
i���mD� �Z�"�R0�L!�B�*U9���'A���,z�p����4��Ims���c�ۄ�a]�f���qV1/�X@�K0cCx�xz���ieY_�� ��c��Δ" {�b!��z����w���$D��,1m�+Mv9����B�z����U�����b��=����3�:�
�G�#�	��ԟV�Qt|1�T}.��}��-,���UB�n��\�܊�䜔OoOW��#��Z�g�
(�&��FK��V)d�Q����J���⫞9�U�+���������m=EclykP�RvAή�-#9�f�>oM�.0Ҳ�+u?40amۦ?��ș�p��R�b��|&0b����}Gw��(���PVϕ�
�_{Z�Fu�D0�<{Ou6-�������۹o�(��SK-�xj�Y1�Ï�`J�v�@�[�`᧚����6��_؆�#��.���\�TeN|Uʣ������2��9�O�&BK{�o�+���R����?��Nɽ���n3��AS�<�i��^9!�X9P�ę��.X,�I]��PU����tρe&J�R㘸�j���:l.��,��4�%�����Wc#�����+��	Lү���-V�ul��c���X-8;G���UgN��$,_�8�Z�����V�E�N����HBN���1���{������>�+�A�h���qZ�.��XvgL�����3,�^��T�*��q�1�V��T2;I�N.�F�0�����H�̟ë�ӊ�S��I;�'�"�b�>}8+���*�9��M�&�y%9��d��K�ae�w�����Ч��v��sb(�0q�Z ���~s�9���U�6W�Yr���e<�4�# �w�m�hwت�9m/��~A_����o�6XҊ[��Jt�x	�L~iB:5i�ޏ��afD��*Fo�p�@��z|�J&[����4xi��K`�B|jxrk�� ����`pM����T�`5[m�o�WT������w���9��3��"l���Cω��Q-�z���[v����Rh�&��&z�=�4�Fk��=�e�r�W����G��|�~.	�LawH�xC����p7Q� ݩ�AX����ش*��h8w�ȷ����Rflٱ��ԵrMxݯ�D���p�6�#�zs���A����Ia�"���x?�:U�;���k�]>E7g�L�es�^�z� þ�d���Bkg���U 1#ag1���[�
gڋWV�8��t9.�
��Re�S�x�,�����s�^���{�e�y�?Y�����1us�h�w��þ���^�7e�����~�1�z��?��D��Y�4O�:�.S��=��iͬ8�ud����#7�q�����}	b/y&�˄��'��+ZjX=Z��}��W.~��Gⳣ�H,��hI��kXFz�*ȷ�[dP�U+�5��Aqm���ˤ���X{F��+���*b�DSr����RTm��7>t��GB�A[�i��e"s�^�yxM���+@ڐL�$E@�	�X�6+.�*~���M�%^�x8��c�u���bt準/��S)h�3o��rz��HRF�[�6���]?����qo]�ۿӬi, ��H>R4����{Q�|��;������t�����\�D��|����2�x�_Ch~��Jӓ��oE(p��yU$�Q��xV�����z�1ܮ�,�C~dYƅ��ժ��[�蕅�+�B�ll������bn�eE$X]S� q�d+��"��$���a.9�{sy�=�::̪wh��D��<��t閹��1���ӗS��; 1��.*�4,��|��sN���?�~��o7b�$��@x�2�I�����<A��d,�����V!t]2wx�ER��o���_4���e�/X��R�d_��Ė�]:γ]���n�5�Z?��_�Q�#��;9kǿ[p�1���|js��^���,>�i��.�ؘ�/��Q^��Φ�JNH��GϕԒ:�8aJ�K��V��4�-�F٘9�&�RA��B[�L��0��*7��>Q��mH�U�g�=Z=Px�=��@�!i4�/D�eI,PU8�����!y�#����b�u�Ӌd}�+ç���S�sgɟe�3ɡ�q��$=�uF�Ȇ�.3�A{$#�^'��A��@�D���B�5uQ�?��XI$�ȉ��I���C��Y �i7���|�����
0���a�AN�� �l��Vk^ŸP��M�D��Zq�,�'��l�$��`��7�<oC����1k�ϴH(�4?�B 1x����Z�=~��^����=\l;����A#qm�U1rtU�~>��u{�^�f��.@%U�|���o�c���h�3�St�1Ayc�b9 ,e#��2Cu��䩔����9 &�̤!��z8����||���P˞7,t0��ٻ�&{Yz��}��nw�;����7��P�ډHҨ>�9N>�������l����H���Iɧ��J�ה�]�0�%�&�K�ζ�o�2��С�6R�:H�>&�PB���@)ziF� �FN���@����M9i�Ϻ��f�:�mu�^J�3
f�4�9���ԫ�%��&�D��i�2����t_$,�T׳I��?�﫠�0��}�%��B͔9�?�f�Lꔆg`Q����n�R�b�u&L�����c���q޽J��Շ� �?Uu�_���z�g���(���k�͛���턮E�j�den�x�N�n�CZ�c��0@eX��Q-B5��~@�?m�B����Q�]ᛅ�
�_�X������E���(�!Җ3�8(R������$C)�4��#°���-��ԄH�JW��C�F.z4Y�;��p����h cH�!�;9ei;����5Y���U�Y�'��誆��d�2>���۞�c!����O���:�>ёT�G"�$�����m�#u���?C�q~% 'B��/����:�^eO�v0��׏o�	�dӃv��Z�S��o����x����= 6|�hi�����jY��� �	��/�ф�y_Ꙑ�>/�����|1@Ҝt	��pb'\���"�)�L�K���&,����cT�)�LKx�X»Ff�]8�NS����9K�ŕ%��\Z̙���t����Y,�j7�R9\dxv��`�fYƄ;D h,���c���ݿkT �m52rʨ
��_�xu}^_!��3G)��ŏ��ĬZ|�#'��:,,=�1����Wi����mYQ�z�����q��p.f��a���PQ�e6,����l8������#ų��������%�)���g�UuBG��I�]���r�&'t@9Pg%A��3ى��~��3�,�0ߎ�k�
���vY��qixx������ʘC3�;A\��{$����}�.U�=.>�)�]���R�I2�D��7�1o�� ����n �Қ����[;�}Q�"�0��L	���WFe�����eT��R���\�)��9D�!��;�NުxӞa��c_8��U�̉�&]�1�E,���`�b{I�0���l���Ƌ�1�i�@�8~��b�����i�N�ܹe�<�4�|� �<kn�y��@j��W�oTQ���l��3�^U�D#�ۏ�s��O|�9���}�>N:j��v�u;�@����S��yiҡV���=W�L�0#�*`ߴ�j��HJ��n�2�U
���0UI<24Ʈ1��z6�g����R�5��L�R-�DdK�ػo��|&��]<���+e*�Y��?6�l�F���S|�^�9~�=+��2�{o�1�
�J^?1�ɺ��2j��kFtR�D��Հ���pߴ6���xvv���2�����L�Hl8��S})N.3RV����������E�D��{���N����2[�
I��I �Ts�'ƠЖ9x�¢&&P|��j���ia���m�I�l�>��&]Z�?9Ŝ�>�������"���w�a��D%�!	H}Iad�J�؏V�q8�}�W��mc4��#�k/�E3y��������d�M�u�9*o�UO1#'��{��>t���T��*����y�f*g�|'��4]7�X?�]RQ}=�6H�wt��&:'�G�8[�(�e�Q(x};��ƂL��0�(���W���qt�����Xf���V[KF�Ϥ ��w2�M,��a*� YU����q�j��Ō5t��x��u����MO�ZC�����W3a4.+��Ia��a��h���ǟL'�8Q�PK�������{	]p�?(*��^��b�~,��=!CH ��a�㲴���+C���(�4|a�9�#R����o�Uz�~�y�Wd��7k#AFܾ=Q_�>g6��q��+�eKHԡGz����]6����qõ��Gn��?�?���z��3��aԯ��]ˠ�'��pL�jү$�~VҽhbeBق��-TX�&�:��)k,�4��w��QBVoʨ�4=pa6z�	k���V9�Nv
�~�ö���J|�����B|�Ǌ.��
�p��d�W��㡋�YR�y�����^���F��O:��B%&���1h�M[:UA�kz�Mc����v>�����U|T�( i�1\�6�Y���jcC�uT�\y5�N�HX��*0�;L2�5į=�	�fb��29���Q�A��u|}�"��=LzW!ιò����/�8xp�9'��|^��:���Kx�ЯvP���-ɽ�߆ ��%�M{K��V%�t�v�ON�|�Л|*�]AE��)� ny �/�>Z'A@�İdln�c�[#j�V2�O�;�M�� �2�(��&/w����	� 7E��\��D5o�ȸ�����^�j<��
�4��Ӧ����(_���"�\����!1����p�f���V�l�HA͹��WZ���4K9g��أϿ�;��q#7ɟX��"3���i���� ��P�D
��x�7ؚJ�Ĥ��Vӟ��	"��{V�t�6M�3�� w�YM��4_;��oU9�����9�?BAN!����j��������I4n����:��vJ_��f7�v�lQ�.5����2o���B|C�7�U��[u:5R��� O�j�{���I0��^��a��5�V��%(cs��{�P�
���WW�����&nS);=�X�&���p��.��ܷ�J�m߽- :1	�틚�"`sl���������{�һ��.��,DQ_�^���qVq=1P�W"�4F�8�S��,��H�U;��Kf����[���C%m�˶��q�MqG�=%�˻k���ߔ�l
̿�lIb��[��zj/�;����ﭭ_��Y��՞t�;��h)[�4&r���քO2e%p*ˏm��~a�i\|�����̳n*�qԁ�̀I�s��:�O!"�J/v�i@��E	ˏ��(}����J߯N�e&�e0s�|�����wf�}��C��C`���"R���I�x���@M�(-2��a!���S[�m(oEw�'��^�|�̴�?4$��b^�y��7�yi��L�U� -����3?�y��b�m�G*�.����d(���$���|=6_E�nR־RI�}e�J�)�A���.�$,���&��+9�1��ݗs'~x��ս(��2�/z�t����I)I��.���B�6ȣW�!�rg^�*ZN����c/G)�+}���t��s�����A�rЅ;h<l�>��" "������w���ǖA�~2{=����6���u�/ES�U�)�2�n��x��m�u=2�E8Ԑ�z�,k��5���s�����4*n���=������y���mӃ���9���*!t�fHg*�' ���L���nk��>Q����}�N
��Z�P4H��ى�-ݤ���$��[#�����辗Q�@�]�4'�(=q�Y5����әx����s-��h:�
qq� ��
��U}o�QM��rW���B����z�M��RyyסhZ*�P���ƺt�x�=�e��K���di 4\6͢����c�A��U�(�Y^�]�=����s�	,���߁�E\�9S-pL��ט��eg`�.1m����o����@f�i2C�=4�+0�`r�0}��x�|��{q9Nś�߃6D�N� ��b��91[���/?�7��R
�7�R�)AY>M���p���@ �aLnZS}��5�Çw���J܄��7l���	���r$v(�?L�woC\�����''�	�#,t>��W������{$� �vc1������]rG Gu�U�p7����eפ��g�b�(�@ʢ�?�aU�y�U"�� �|��!0��ve�W$D�F�1�l� [8�����{��A����L���_ŦM<�ܩ�6�H<aD,	��T��!a50a���#�?��B}��fD>v����w�>\u(���]�n����0s��˵IK���a�<>@�@��L��zK�r0�j�����o�� ��H%/�ח��I��& (^-'�w���{ ����ON��BI�F}��O˗�]�<:��Z���m}A� >K�#���J�$;Dqqv��!o�X@Us�� N9*�@D�̑���\���������D�����n�^��%pFZT灛��e�9��r�	��ړ#��K���h`�tML��:���.+��D2;8��r7vX^ �'�C��+ٝ���T�0l-:�r�"6&2(Z�]�u`�D��o�f6��wg�Ni����,��xڛQ:�@|�b�4 *�w3�'�}}'6#s8��Gy�1��h|<�Pl#K<F�u||N��M	(�b�\dd�O�0w0"5ј�6�";a�v=K�f��O>�&	c1�H��j}D|!�3�OB�ٓd�#�S���x�8�T��;C�Ꙙ�pכ�����?l���k�.��Rd<��t�ظV0���u1Iᖞ�L��"	�,r`H~I����C�!�u�Z�����I��;P�亱]�o���F3<�v>���`,�`�M��Q�(�Grbt
O��h�pc3��J'$�u���b�8�4"�dٌ��:��=\<�$³��|�c���4�WG�?�T�-��{���ϋ���q-)!�9K���|��D �k�ק�xZ�ӲM9YEs)g��#@I����������1�iքE���I��BL؂���mb�%��F��ѭ��nh��d�/�{�|���b3u�n���j㍖��J:�=H�2_����87;J]NӒ� A���~y��?C�hJE�{��w�Iw��Q���Wgk�xp��;������7c�z^�/�2R$�q⌓�B�#ܞ�E�@ո���o���_���ۆ�4S/_h͊An,�O��K3%��<��_0��>J SUvD� }�kW���R�3�`.��^��0�M�Z�OYT��@�v)�a8[aA�;�`C`RO�����j]�@�6~��c�Q�����
g6-gD3��_�zj�f"�a��5�ϭW�v)$4�q��P-O�*y�s�g��P�杂Q��9]tG V�HJsP_�hЩ�Z�e7{��M�x��I�&Ӷ_�%T Q�I�&����}^��ȽQ�FUs��j߶��mN
{Y 8��Z�i?�D 
�:���bs�B���F�Z$�z�'� �N2�\�r������u�yf�72s��t�e%P0-���06�3Ť0KN:�,P�*07��t�v�s�8��HK���o�37.
��t�υ����'��-��_;'���׍G8q���#�CP�Raʖ� ��T��}3��D9wDk�5�MN�ؔ�9�5�iY�'�%�`������.<3����XȤE����O����$�{I�T]�(�ɟ�O����Qy?f���Iq��"��t�	t�.ޫ�D�fR�{t��P��\��� x�5����a��9��-�Уu� �T�q�� :��*I���	ϱ�RWt�K��ޕ���&Z`Z��λ���a���üx�x�K6����!�V`!m�5nO����Y�H���;n|�����e\�}.���Br]���+�۳K*K� c�Z����:0E�E�g��)&doR���N�����KS���¸�m��C���m�hm֤��_!'p��܁���$�rb����]B\�cm���|L�`A�h�om��ne
�m����&��<����d�;�]� ��	E�xN���L��o�y��n?)�I�oR@�'�4LwC��e�z�3�۔E�����^���i%�xj�K_|F�EK/�4�[�yՊ���H@���AϠ;�a���`?�o��"����fZ�ďH.1 89a��h��gl�Emc.B�d�ۗ�M4�ou���&w3}+/���Y��&nv�3Չ,�m��߫�J��d���h�+�fm��mC^&��yF߽�TWΛ�=�v;j�<�r��O��x .,d��Yt��|���Y*��[����[��`�k,��`L�#D݆��E�i�`.c��i������љ:~�Mc�R	P����3�?���c�aX��6���z	D�R��'�2�K��Q���n@�rڈ�
�{$����W�����`f�5jȼq�$RE�/,BoT�99f����H�i��7� ��KޞU�L�e�2Ɲ���գ�]���.Gs�ŏK�|\�x�+!U�O�����]�z=�u|�JjL�07�X�O�$�wҏ�\jV"���nM{V�&sV�;�n��`</��
�2<HX�w#=M��.AjΏ�@`HT�uF�ͦ
�)ݫĂK<�!�Z��r��W�@�{3���Rʶ6(qa�e�>�+I��l�j�D;�2����MDr���H\0��J�O���q�ƶ��Q�[r��������aFm���ϒ��$�����Þ�f�ʈB�|hfK�����&�t	�ț�c���� ���淏@�Z󃈝�'��ΊU_B�q7��3����Tj��g�.d1ط')8Uo�7�R��NI�����%����"0�c��=a�P<d�5���s��R�P���-�ZV�����˚<\?�(�v����*�N�l'!Ƣf���VU�izYӇLX��k �O@�/�7�(�Q����GR��~����P� �RP1�
�|�I	Pzԝ�yy#�����tW	��:�@�7��w��� ���?�*j2��!V��AN�H�xy�'��"�YҐ��)(�:�	O+�i���m��BVoa^�����Sԗ7K���� �)(R���bC�ɹ	Jg_��D����v��g��k�F� ��l�`��+ב4�����J<�Lq_o1H�OI��[�ڌT�>ث����!�sV(:1D^��п�j 7�iݕ��>Gt��Ak!m�V>�����E�jt���~D9%cC�A��r�m�a�
N{��g��aBuE�(���rh����!?��u�D�������K��X��Q���c7.Vy��& \ $�#�S{�{��u0e�V�/}�A��C�'6��W���f�S��ǿA�i�ԭ��Ǝ�e�gJ�$F�+[VifЯHN��@�����9�c��9�w�|>dR��ko���Xi;u&r#8Z��7�JE�ڴʼ����*
\Q]<�#�"jH�,�&�{el���i���g�Uv��R�xP]���0��..b����i�\�����&%"����%f�D4Bb��}1�&���׎僐����"��I:���B-��=\�!��+J�Ή� V�ş�K�B�Ԗ�����*p�YANuȁ���?A	��:�����:�{$C�Ԯ.GhI_#�{b^'��:�h��uIr��M>�%�C~�C�r����oHY�J��:���~���q׶(��&y'IS�A��s�l��k�V�5��/���V�v�%���[
��b�MKO������s�s�����:=�@=I����X�1�݋���X�|� p�u宇r�%��׽��	<�Ȑ�>1I��FZfF�����.�yy9&�H�N%�qf
KH���'�0��U,���`f;dz�Hӓ#5[j��q�EA���([��/�)�T��+r��Mj�-6Sg�"QMO]���d䨯�A�I�Ľ�%�o�!��J��\���x[�c��E��Z$݂�����pol�^�vRQ4c'�[����;�0_l�^?���T�熭͸�W�����9k4g����d���>��,(�,���{ȹ��#�3�әԘbW��J}����*�M�����T�U|e9F�K �Gف+�W1�NB�p��w�H��lպ%>��0{o��)�&��v�b��f�x�&
�i�F�Q���p4R�i=;ŇЗ<b�����͹gy�K�L���!�+&�P@x�x�&�Nm�ȅ�s�>��R܏A�:7/.4�4=e>�Ek��«��WO�
��.h�Qi/�Y�<��TI����*����b��s;�ج#�Δ�kJ�����ɇzH��sA��I�6��&\Id^m8����<uCyy?�%G��{�V��c3Ʋ�P�(��������x�9MqS%����c �&8�X:��v*���̪L�^�:.�*��Gxle���~{O��N]~W_752�s���S9F�����\���U=k����^�M���qe��a�%���Wr�7��u� ���Ӈ<����e4K�UV������@�y��ތ��=�xi�0�h>�S��?H��d����j���N�[ީ�n�mtY���!I��lk���v��N6��|�!hH�x���mS�t��YS�a��1��st)�qU�2Iu�/�z{������yؙm=���Vd��<�<����YO�H�`)��^_�?���٥mm-��;V��<B�VVá��VnN�=~w浯�F$�m�'����1�:&>�_�c��q��� �7�	Ǯ�BHV�XKC+��g/k\o��v޽0Y�*�:�X��l��s�K?C6�E;��lsyA*W=:CS�y�3�Y��=������~Jr�b���_оGM���~B�K�\CQ�S	�_��#�eI\��S;��n�"�*F�?H�qR� m���fi&9�j]g���k��x�� &�kB�y�@���[ep����kb�����>I�#@��0\S�NKJ��Yc�O���sA�.����~u��z����g����,Oiq�	Pޛ\��|���n~�J��<J5XjU���p��B��#��ڡ��M��72�����X'ݰ�4��3�Ɩ�7��ב�[�1[׋#�v�=z������jc���DT��X���t�L��+c��U�<K�c*���}ܧ�����x�;�SiS��cY�,>��{�/]H:>��'�̯օ��WVᨁ�Г<�+l.hw����jx%�a�.r��CPb! ]8xd�jM1@s�׀4�n�(5��4n�g:�ak�T�{���E�&�`@zU3�+�4�j�ѳxz�D�o�Ʈ`;h�r0�O,ѕ�f0���B�~��9��%Tٓ6@�N��b- ��%���ZA�l�W!�v�)4��^*Y�n6�h��ri���#��^���('�:��]�DN���h��&,.��r�<�o�:�h� �s*5�%��' ��Ru���5-�Cd �$"�JtG����Wc�P�/�;A8�r���^g3�g��x����5�/��S�?�=�5}��I�8�(���O,l�Q�W��X)�M�H��M��B�C>��h�9��R�8҃O�JhB�7���G`7 �PJ�Ձ�����:.4�{;J�{��9�� �$<^��ׁ��y�+�O����Dnw��Z���x�S�Neɢ`zY�94Xۭ�ڔ�\��U�*��9F���� �x��Zݶ��=h@�v��^'�MY���a��n��.jn�⺼��9�# �6f�'H�+�7�k��/)��*m1
ǁ7`�)Ke��!UK�7T��n+l�����&c|��@�EʠW�$��,�-ěg�>^8���n%������p�}�>��e��PƯNvz�l~ņ�&-�tQ���oB���%�)��r�*��&O� U�E����J�؈3>L^U ���m� GCfm�z}����簷�#�X-�s�/�I��YǴ��h4j��Q�B�H^�4�7ڭ!(&���v#!��4�11�	��O�!���44�ca�����o�Nk��e�`�-bI�V����u�w[�b��7VjG�<�fBb[T�k/qѰ�Ӭ#��u ��n��㢜�b��[�ٌ�{�.!�`�-�U5%�{�f����"��K��[����AZg��r��+���+��:��h�ZR�C�����Vφ����^3�wt
R':�����ڜ�3ᖸ��(�w[A?ojh��:n]����v����#faRl�XS���K2�D"��oW��j�px�����A���+�cc��-f�:
�x�J�32��2���jb�R�%ą���^�`��5�C����W#�H��>B�!J�K밿��2D�P�h���'e����R��j4�X?�F. ����F���|ҍƽb ��� ���<�Hjj7ʸv�G&�ma?(/r(v�*�@�k>����������C.$�cCX�wE�U?���)�q�<8K=�>b_��l:@�X���M��:��8�����NӇ��iXO����l�q������	\��,���>�a2*=��p��t!m9�i�P�T����o1�� ���)~�rh5o¦�V�Ko!0�{���n�|�ޖ�Ť���y~]���2��y@����M���i2��;�+��?nGx�VYp��rX�t%o|��lE0�?�~� ���n�x�0 ؟	,�#�\�%�����@,b]�^�A�7��Ѧ;<B3�,Pw݊�&
�׾��c9�!kkZ�XV]��0c�����5L)V�Ή���{u�l�,Y��8�)�����,w����kq�!RJ
��l1�ɒ;&�<@b �ꕗ���������5����٫�	�jgPg�����$��+l��]�$Uxa���tĖ�+a�J&�|8�і���Y�}H�����w ����(��fg��}�+��H�^޵�����R]3��(F��_����'����W����,�nV�X1R�-i��j|-�5��>��\W�a����9��p�i�o�pƢ��NrQ�'�g1$�Jx.]@�O���d�(�̘l��̉�>��'�I�)� `��R���J{qzr�󇉣�5��l`'f���޶����HiaF��ͨ�z�q�!ϖU+�-�/��2���1�KKŬ��ֆ�T�nx�����d��Ϛ�9/vOl H��rH�M�j�\����/jb[��p���V�\�#�s��Da�f�1�����Ċk��7�ʾ����C�k]�%jK�sd|(�%uO��4�B�����>��r����O�7#��d~���B���0TJSv5��%^�`\vD��#4Q/��;��`����
=G�&��'}���Z�!�ܺ���D�~�5���+K� �����WX�=K\µ7//qC]���A[��ub��4��f��TY�V�$�Q��Tڡ�w�"��P�������v����i_˛���(L&��F��Ei�D�L<.O�^����!UUx.ȩ��� ͱ첢���,p��0��53������h�p:��f�����|d����V��k}�����+�~�[�]zs�#�s�0$h�hgJ�yC1�W���>�����r�!��"Ҳ�O�_B1��z���\&s��8Y�>��:��秊=�4�N���eَ����V2ez��+�#�Q���;�;���Q2��YMN���ύj�c��z���_�z���|�KPwǔ��*�Z��l��Vy����]1�Mᑥ�k�69���V�9�9��%�Nc*v���]���z;��H��_�8\��ȲYj*��L�<������_�^<\8|;9%DGn����r&蚜�E�o��<�pYv�n��93|��y��P��Tf��Q:�����4���V��/"�ka�>�cA�v�y��h\�����_\3qz02�o�'�b(8R�Mc�
�6{B���uv���ۧ��h�	�l�kNO�YK�������o��3��[��K���[;4+��+O�de��Ib.��N�}�,U%�P�[Q�Q��@�o���T�S�m��ɕ�O��H2p��Ѥ0 �j�qI�-��R�����P�:���ۯ��ih��e�q�Uz>�p�;M�?�h�<��$�9&>E~d
�/�Zw�#�o�|��Q�d߯�(zr�gQ[���}����q�Å���"�=ᄑ�(�����e��|*�<�LM�gֳ��7��al�&��[�k��	��]z��He{o�$�E^����}�IZ�.��X|yQa3���げ>�}pZ�@L3ߚ �lXg���%j�Sy+��V]N���O�\�cx�T��##$��=����IQ*���x)�Y���JJ������	��;IH�SЋ���f�0��lv�;H��(�C���X7�3��Ry�95�U���Q��/=��\��߀���6���#���^٧�o�O1(�|�m.0�!{��OT���(EW�wN�js+�Ó*}�ɜu/R���s��ٚ^�İ��9�#����ڬ��=��g����ޛ��fF@@�������
��S2��i*����`Pϱ<�1Z��?��Ç+\4�i_+L�#E-$~�X[��.��9D�6�(�(*�ڟC	B�z�Ct+F�X�ϳ�?����h�m���C�#�� ΆU�O,:'�_���M3����_�ỹ�����ׇ��
��7��}�:wm����Ƹ|��sɭצd�x*V^C���
�4b�ƿ���W�t���D���13A�ȳD!X�y��Mc!��iAPS|<�N[e���z��{��c�'pЫ��!��"��)�0�ؑ�/(�O_� JE#;Zw.E[�Ɏ6�Wr��A�cQDZ��6��}�����G�*��� �Y��t����6�;U���z��� ?����o>0��F��YQ|+sc��%0n��U���5^v�ar�HTIW<��6�yW�hk.�<-B(�ɘ=�'"�Q����^�v�����%�r�C��X�U�S����Z��nF���9�r+г+0=W0������]0W�Z�_ڕ�m�MA�*W'��ӠY��|N���"��<n'�-��_)�I� �&�<��n�_Ϳ��kySy��ҳ�2�p�t�>6Į����^�����D��x�Ks$���I7�hF��u���&�1��@��Q�tǐz-���C�����n̄ۅ����6�Z*T��͇p�7}�=#G4F5��R#�x�v�mמ{Pv����TÞN42��_Dŋ���J�.�Wk��3�n�(զ�w����bC#�9g��߅֙�:�>�z�����+]j�ѯP���We�*�`�旴"��i��/c>�"���?\��'e�/���di��H� ��K�i}�ѩG<::�1�$9G���gI����
+
r��S�يk��veK���K�$Y��<֔����m����f��2s�2>%ЁN�q�ܪ�1�&�K��[C��^d�-����P�p%�i���&�f��*��N]&�=B�����U �ύ��=w1��&]��:��,}�e�g�?�5X2�/�n�Ik]���>[���g_=��u$Yi��}M��k8 Ѵ�����{-��d�s���:���9@x���!Qӎ:	ˬ�{G�A��E:��?.{x1>i��5�;���3��^<��i�aU<V���n��y�}@�0� +
��^��0���^b��e����梵����\ʰVd�;�:Ոt~���I�@��{#���ky�/�(���Pɷ8�u(�?v3�˕������)G��������kH�n&��։�ߪ�tj۹uH�#�/HV~/q��լ�m�y��/+dF���b���(:1X�����C�����c,ubw�E �E��ī����s�|iJ�/����J�Fn�Q��N��!S��Z��ܠ�W$���3v�Q�-0��1������"~[����Ʌ1׭�.��l5�?�,b��t+�5g�s��O�����4�N),ߙ���8�׌��{㼯�֫���N3��	�
,�P����5i&�J3=a�X�E|�cb,��2�z,�ǣb���'Cpl3A�I`>p �ehG��������V�7�E���8�"d�n�T�-�;�8�M�嘝D��"&?�( 
�!GG�4T5|�A���h�����,�Q�e���Y���^)ڱ_���y�`n�Z�[EGǕ��6������#Gez2�U'�;�ã����2 b{Ge3���L?Jݡ���<��tg7.f�|��=�J�_�^��?�F����������&�k�Us|k��� �N5r\��E
���()�^Q)���~c��h�X��}�!ҳ���w_�I�G*�@�x��f&1���3M��D�Ԥ�Gѓ5ΫY�������
 鰧�)C|��R
)eG���\�Y�p����|zo���ub0�L�c�
Y<-	�ꮤ�H��_>ܷ�̙v��	Ҭ���A2�����<�<�H����S�3��������5�����v��L�4gE��׌0e�*��Hy�%���ִ�~mت���3ȞZ+d;V4���f���Z�Q�a�t����jH�tAk���n�����3$%㗢.�\�)��]g���Ra٦(�b�͡�N�����^�i�њes����o���ǅ�1��O^��LƵ����C!_r&��Q��%ԍ� �Og�=����$�5���3��'��Z��b1PÞ����^pT�?���X��W�6s�Mf�梖��/&�&XRg�N��%�tba������L���l�\�ixwZ��k#��z��,;x�l�a|U��A�J�:ɜ)���4t�;5���W0�wA20m��-fB�����s��v��]�v�!t�t3�L�����/, 7��Au�������_���	�T"��Џ�Z+v�z7�Pr��z��q���iKC0��AsH��%0u�淗�;2Fa��wY�*�������NMs�:�����V�\��`O�}W(;�|�́��}���-�c6�	�-G�h�J]�k���ZJP�uȺ��qG��u�.�g)bM�(i��d�[{����%�����C������+��Qq�Jfr]�$I�p~��B)���)-e�n<����A��Mf[����N+g�[����iQ�g*��s���36�%5��J�n�a6�Q�P,��ٷ�]�k9=0^8	��S�Ձ���t�i����ς��
-4`�r\�\������<o[�U��~)�ѩ*�_@^}|���ٷ�Z��q�aԀ�7���&VJ~n�AF�u@�E��J��fKap�A�#@t6@	��Br^Ѽ�|1m�<A��z0)��E�|��+�6�g=�X���鍆�}oP�u.b�?��R%�q^哜{i�)�o�ou�i�<x-����ֳ�X&XWXG=�t�d�.���fm�7���S�
���x	�琖��!	2jAv���%V�q���"ȤY	1J
S�@�%�[*���CN�;X�����_�fkPEx�3�^��ʆt!Ӽ�![����j5B����AE�F5�������Ž�O�үˈJ0~��}J�.�v�3A�+=�N2��
���o�m���i{r|@pM�Z#��l��g2�9[��a��I?1a��ngk�VY��E���E/���.�Odw8Mk��� c�>	���r�R��~��Z�s���#�%d��(����?��[�2�H�2�Ŝ�������/*s�CTi;��[�@ۚmE���S�P��k�;�D|fEMk��&&��Z�C���!OF�նjL��0��ڗ�?e�Ep����ӪE`��S���W�K_X�]^n'��=*��wD	[�v	)�;��0�Ix0=�~U��PoH`�E'�M����J��dv�81�<Ќ��7W�7����"H��Lt�v��7Ah�gᾸ��x�#i�y�.\P@�����o��C�י��T��7ʊ�6X�S���ZC>�F�V'I�<�71���R=���Y�Fx�Aso/��.��MN�(3^I�Nup��?
�;��P\D�a��Ӛ�.�_k��A�S��Y)��("7�x?��DZt���O�(�
8��сP�d����Q�&�A!ک���d��'��S/���L�f�a�����rd�*
�J��_�ɐA����]^|�%�N7EW)������<ߨ��:�~`���܋�}�+�:R]��2�T/>[O��S��6��@�9�>�d��#B��
b�,d��@:d��B6|�3�Ic <�:!�A��>tl�P^�6��}	��O�\��FD���	��(��y���IV��i"���;�r�ù�{�Sz���-j���R��5i�B�=�f0���l�����'c|�I(I�Cla ~\�(�p�4qJ�߾TĿ��n����zK�5��+��:Y�B?(��-3"�c��<�'��'oBbM�O��I/Fe2l9�(���Zmڬ��ًX���ڥ�{9W���y�����`)��F���Ț�NN�σ�r�+��\�h�T.o�f�46�Ţ�e�-���QOR��2s�V�y�y�U�Mל,k�5d�aN��a�i���nEu�|��٭��x�)[~dA�[�'K�T�&ΡS�LI�Rv�ʦk�~��ӈ&�Aet����a�5W.hfWg�'�����Z�	�zK=(��~`�o	fj�Uv�lR\�@8��M��x�/��4�T(��"TlT��a���c�1�ͧ�0�M�dl��J�j�>�o��Ȧ�m	wuC�J����C��'�C����Ch3��LT�6$�ث|g�kn����u�
�8{ېiǃ�CU�@�Vfi�'XhC$�(��N4G�����ǈ5BZ�JkW ��<1
��'�-�wL �k��=6�&(m9J��Aɞm���������a��i)w�|��)ac�o��POD���uÛ���dV5�2���h��͎��2?�`1�m�9b�J�k�X�kX�7k-}9=��/�kGʶ�>���0�n�_[ �� �|��SJ���U���5L���Q�,�;b��� �ǁ��,�`��ƣ4�hj!xiO�WNQ��Τ8n���Kx�� �}B�yc���)ߔ�w�s<l�.�v<��I� L�JR��	3i���Hu��)_9����x��֙W����~%��n�,.��d�G,�����p�