��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P��v�"<ߞ��&'��k%P碶�R�ӣ�sĞ������FY&Ś���#����,h&��[����W��Ⱦs첽t��w��]��rLT��z%?E �Y�](�r�n�(�bIaCJTƢ�i!�73�n.����0)�i�Y/�\�Hqk֭�p�#��+�����Ԧ��6棍��#}#J������Wc�2lh
��*�� �5]8�_�9���r��v䍁��@�#d4�_Hz�0������K�ݽO��Ѧ�+�ݺ������nI/�	��@��!�
��,џ��.��3c��K�v�룎�"�3���|�p��u���9��{�ol2����ZB2�(��x�T^Դ�� e]���>4i7�M"y}H�P�Zs�O�j+�c�JC��Ll���i���I�z>'���˪��.�ys��n©r��|y�A��	�/8,��z%d[}�f<��MA(���P�*���aM^Q��L�.zy�a!o��\k�l��V9[�(�rSL1�����̻nB�s_h��]��c��iqb4�V �"��ir5VH���:���C�Z���4�:�R�K���RN��p�u^�仮���%�l?���L�Q�Z����^��ST^|8W�T�<ӧ���]�����c�������'.����`�����I���d�,�,ߗ�����LЏ;Xxhk�hk��'G����������(��!8ا^J�ե=hv�u�oO�h��L���LEv��Ծ(�cj��"+��A��r>�DU�6oX���K����0��GV5�l7sȦw̭�N��F��;���D�����ܧ�t��'�\��-�j��
 �Tq�������>p��W5��EPhWu?���-�d��iKf���.��3��If���+�8M"?�]�葈�K [��-	����Ipr��X�cP�J�E��^��J ���P���2
nIk:e�Hw�eh��,*��i3�F�du����
������I�a���(]�cM0�x�=$<��ﶆ��ؼ��M�R�_�D���E��}e��-���A}���)�B�ֿ���x� ��-U�� ���� b��Aۥ��6.@*o���֓
�C� 
������b,�~p�l5ȆN��7R)w-3���J���&�}���-)��`>��x���ǭ�@
��\���x[y�6ц���B�}���P�b�3cS���"���U1�±w���BI�y�s��C|#���kP���{�(@L<޵Z(�p�9qT���d����S�為u���F�v�]F�)�m�6G�t�C��-o��Zf���l1�3�*���̅��u�{e�Ă�G�~�i�NW�Z����9���[�W��"��! 7�؜cr�ynv~`$�|i��ᤧb�D>��(A��po�9D�:U������݋�X[�K�mf�2���_b�$K|�����="ȋh���(t�R��Z�Z����w�o�����=��n�]�pRzdp�H�[@�$;��moǉ��X��)�s�P���*��h�
�	��{)�(��r�w *1�9��9є����1Ж�"���N�h�b��%�(��9dH>��4�=��^ r�J�nmo{��z�G��������ڮ@\N)k\<-�-��˶���^S�/��$�P�����8�6��ǄXz�7��1T����*;tӜ���ѻ���{���ٳv���D;d��.�D.��Tze�,�b+�j��%���&H��8i��5$gE�\��N? �`�(�W7�:GNn1rs���^�p�aM5>��S+(�տ54���&,Z�2KH��Ǔ��Y����y:�ΰ�x�	�?nm8��bb�<e(��v�s�&�^
��1a��IQ<c*D[>�:4p1�r`�m��*�À���`�G� �`�����l`�v-c%EJ�ֶ!έ�W�f�5)��;C�)S(��I��%�w�?��T�Y��R�Y3��%�㮲�E���x��LN�ߝXQz7T�f���Kِ�M�^ge5C)����X��Q�;�v&t������+�V�H϶	�g�hh���y&V_��w�j�1���Gf�D!*����������J��Ŗ�7�n:�-+ey>�;�)�FhP��䏋��d뺦Vv�C1���~�#�����`=Ky�ΛG��[�i�cc�5T��~����ӽ�d�#�&�[���]�5�Q"�.�u<j!r�Y[�@�nV�+��%u��L��z�7_ĵi��C�$���.�d�B��w�O�l aB3Kj{ܣ��BOūzτiı�����g�
�9$Ut��Nf^�[z}���/���TxP�pW�#�ȩ�v���D����P�,�n+F����#_Te\M�'�WnS���R���bP���ms�5Y�Fzc�D�)���`����9R7�+1&GE�%m7�q����`C���U8@P[����ܑ�W����Cذ��������pdBW��k�.'�:�����<ﳄ�+lM{��o�M�#&JέI���'aLs�uQ����5�n�	aUP��پ��٥|��Q�̮l���*��	��KVc�E�ɤoE�^��<�_����X/���
2����¥ <HNCy���Dx;7�����	�j�ȶ��W�ٺ�����ǒe��@yC��t?�~�pq[	�Z�N�2i1����A���E�)Mi�H(�ÀH����p�q��|�g0TV� TLJݞ��7�H�u�b�k��E/e�O�r2J�U<`��r8���/C������.�5���כa�t�Wc��g�$0�a0`J�{0+z��*������F��z֯�!���ӻ=�z�R2����;&!�^�X���+1w}TV#��\��f���B~s0�#�~-���v�拦�T���鯹�[a��4r���՝��k���Z�W4&Z4�/#I�а@������1��(����AarۢıJ�ʙ	z�D� mY�p�1�+�;����bR��b���v*a�}Gi�ԻԤN�q��IB �4�O�h�P�yWh�mX���@�R)�]���Dl��뒯֞ +�yF(&�hm���������7��vA_�����]*�s��Ed�d��
}�K�`n �}�9�����݋	�R��#����S�`cם���hN��4V��0�
tQĉ���+�/|�g
u+6�L�b�I_��'�
�#�j��E�;���G���xo��!I5�0O$�<\|u�i�  �;;���Ϧ f�^CE�����/H��(��Aw�;OG蘡���ec�E�p�|�e@�h�G�
�@�"�D�i����62G���h� ���J�Ө.�GX	͏�_�L�"���De"�
�*�{�m������zI��n�<�WK��M߂�Y��� c���zi�at�2dʳ$y�����S�mߧ[u�T���l�#�/��P�ޫ8+%5&��>����[���Qu>�0��`�[jƅ{-9C(�]���o-���'���g�:��/f`1`If�QV�caX�t�
u�vJ��I ��P#�V��O��qH�$�N{r��6X�n�N����s�~8ԷF������r%?4��v]W=����'����i!qbP=��9j՟*�&N'�/�|�n��jР6�NM~vW���q�Πj����)Vf��	��.�G�#z鲝i��s� ��SS�w<U3֪3���/7�_����[XMB����[�߾峈]�(|�%��'�.똀U��"#��7u(�>K.a�h٫w�RW�W��o��יL,@K>ͷ��* 7�+�x�ac)Q��[n*!2�I�7�Nr5���
`�o��e�]»�A��v�#7O���B�=5��]��+=mNέ��A1Rw�R��>NV6������t���Qf��T�3���L�s���su&�}���9�!�7���C�5gT��ecϼ�fQ�,��1�6�~�p�M� ��^�������ŕ��`נ��$�q��9���W�<`;�l~m�,(5�\4�>ޕ�Vp�=��0���ٞz�?-Cщe�j<޻9f۪�	��DN�	��I�M������]ܘ�?w�HF<�52%���������p����#o�}���:�,\zc;��
%��oG���͉UB��Q憟���9~j���"�E=�n�7���Y��2��@��m�/c�A5���I�GH6?Х���ln.�C�~
d��I' Aq���j�ɔ>6�R�H|�C�	�G�C& lu�������l;���<U��<zl����OÏ�ré�F3��1�c���N��ZI�V$A�EÊm>�.T�[qo�h�\�Y.���z��쪊uA�/��4c/����o�[sZ.w'�6p�Ч�,:hZ��u�R�mj�	'�__Sb���Q�內���۹��aj��"@�[�t):���	]޶���S(, Q�Β���ś=��J[p���G'��Zq}���>)�F�w���ya	�A�F�+B����Ğa�Rx9�!W���wK�q@$z��>,^Y�?6p������$u�u#��Rv�S�вj�j�/�wXx�T@<a�֢�g�p�MJ�b�33���k+�M�$k�pGd���~Υ����8��͙��\����P:�w�|�l;5�+�0��yc��f�#O��&r;T}Z���f�B��Hu,s��wߒ�R�wh��|1 ����=�S6�Se1���ڣ��)xR�\^�"����
\�����/��D�]�qtz!�e��a�*b���U�ep3
�,7ƍ�$OM#�ju+Po�K�q�n������e�X�Y=���!RZe܊��� �S�e~qV���[H�=����O��R���~�-��̒������!���%ހ������Fn�ۮ�2�f�t/��+�W���P���\����\��Rr��\8���V ���#AI�/�}E�	����Xa'�	~����l�f"L4��l>�"��(��i.PtAtY=$t��2z��j�0�ܵz�&�����p��	w[�ri^ȓ���7I��t�o�Q��l�0�	���yY�w`���.N��� 2aj���/8�8�i��_ˌ|�0܀�(�oc'.����%P�zr��#c6	�r=l�b�ѕ7g|�ἂ�cޢA�**,+����~��.�lY��۰���]��2x�9�]�t\T���G�m�E蚫b݄���+-"_&�pj NMC���x�t�R���t���_�������UA��$����UIi�{�!n��1�g>���{��XV8�ᔤq}��l)XA��CLFɱ��'*���l���3��H�ŮyYci1���؇���@�������p=�~3��(���c�.6y��W�Y��T�g�2��p��S.��;�WL��������n�� F�1�A��6M�
E۫3�#k�;#�F4��0l��'��%�T�P?e"/�����Z�wʮ�YC�@�{�r]=��%xG+�o���`�h�9YIr��>���b��v�H��2�n�zn��El�[�Zw�1��VteqG4p�����I�ʮ�io���͠�=�	�Xe����b�\ƱS��'fy�0�����{�Q�m5l;E��mtD>��n�R�^NS��󳱠r�
�o�ϝ��ӏ1��G��I����V�3��Εs8��VE�U��� 1�����r�[���M:���P�!s��O�Oє�g�rI�a rV�!�)r���0��0�8k		C�P���<���$�Q	�j��Z#����b)
��r~�D<�����Vs&J$�I�>j⥳	���������#���j�`�s�����u��eÉ����m�礿ܫ5�Q�'2��t��Y=��vJ�S5'A>ٮ`���~�_z�BLk��ށ���k!�b�II#���"�{ø�@�hs����WG�/L�^�{-T�{؀Ԏ��"��BD�w�C����Õd�z[<)Z��҄����E�u=A�}����A��5�1��m�����l��8�!~��q��i5����R�=�\<���
��o˷��b�U���3A���7���p�té#�!�D�	����l�L׭�ښ�G,�� E+����gg�cd��^����IT��Q��FBԎ�^����ǵ|V]
F3�������D5]��GK�BJ��@�3we��4+t�9���/G�zB9^t�2[�|9	�Q�w��*�����Z�87�T|�S�Ü�vk�2��2%u�����Ux�i��j����&`'8+'o���Bs&q��k�,�}CF�\�[��6;��v*�|oQr��mKI�M6����ϝև�D�K�i�U;j�ˍ��H�Ȣ��*�$eka�w^$�1��!io���i6я=�J��2�!�^����G|*��ڦ��9p��(x>�{J��r���w�}�ц���Kq���Tu�P� ���9B~z���7~�ӀfX�?�'����ItP�*ˊm�^z �ˌ��ΊW[�{R�<�}~���>f�Q��s{�.Z��R�1�nݮl�x�m?��sdNc��Ę�{���^�pdl�b9�{E=�:��[�g���_���ma�e?�M;OM �L�8`�&:�����е��8�k��]���\$Z�2�����&���6Oܦ��3��%�= �r�5NGӔ�N���F��N�a�����4Ҏ֦"��Q
Ӗ���n��j�f�G��3��dț��,���Åd�dԄG��F� ��'��9�D*10�����m�e�)�=MjR3d��8�c9$sNU���1�Y��L#��@i����X��g��;�X��HI�X��z;`�7*,�i���iH�l2v��)L�?�~�(g*s�/w�J�@���ח�����{������qhGsFO�Jz{�[��S[4��÷���#�]+߅��t��r�d�UB�Y�i��Ƶ�?��7�6�,q�d8�f	'm����R�|���x?��yT�9o��J����/T��j��)�C��ƕ��E-�l���6�ӆ34ǒ���������F����TK�SJ�� Rћ�ۡ��`/�w�������������_���" �����3gJ�1��>9st����ydVeڵ_t���r�o����{������#���q;��|'�M���H�k�c��e��k������"%H�Gm��ܔ��p s�X��Q3��@n��s�'�y�
(%X��8�9�n��z�)
6����9]��l����	��wހͿX;8�1Å��}]V���V�U���\�"q���*FH�쎲d3̄�tfj,b+-C�#��,T�w�u�1�
v��8��ȲnF��=�xr@�Ň��,��G�qA.���<�9j���؜T�!1#^����C�) � ��\{�%�d���E������V�k���E�(���5��Wh$2):v����֑�f&]��KD�І��Yx<����e��@S�j���%���u	˺����!8�����5HBa_��-x�v�&�3A� P�m��y�n���)ȴ4[5�JDWV���� ��^8�s�z��._y(��dt����;ڙ��-�~t�XwB�&ʹ����r����V���8N�����Xh'��?����[�Ͳ����ڝ���BA �:W����s� ?�aL���|�۱��8O�fq�l��ۥ���Y�<�����M���2"T(�u��r���S�'��2���PΞ#�����$�`��b' $��Q�������lk�yC��E�f��V�r���o��SM���� �}�1s Ýv����<i�s�s��Vb���y�k�Kv������8+'�̰>3�ER}n	הO
p"	;�
Q<��[	����ڑr��g��9��N�\�X%�d�^�*�'����]����^};���
����I��e���o��^ r�U���V��Mr�M�)���7M�JLVb�)@?c+�$�J�*�Q�k���5���c�������V�R����]���x�z��"D�,>�p�Q��oX�HE�t�d���{�s%��MH�n�$����\�|<� Zˠ�)~B,hY��5� ��Cq�Y�E��Pw���%�������Z���.l�V� ���՜�|zG�ǆ����R�XG�O�&1���a��Ҡ�d,��o)Ǡ�sL,8gΞxP��q��8�yKмM%��.3����� y2�F8�NH�z�N�#hs�a�D+�/�[�s/ݘ�^;kq�Du��tn�Rّ^���8��J�5�"���Z�c�9E���e� [�M�=!���c�lQ �T��ϭ-/�v޳V�RÜX�53D܎d�pM-B��Ȁb�.Ax� ^�}�9&W�q5�_4Q" ��60���|��T�u+�Іd
�Y�;�>ٍ�*�`����O��ӳE®���z�0�w;���jb�kLy1Oqρ��hi�������	��,qY���L^2߶R�f��C3�H���"qE��zJl�^W�WJ:��]ݟ`%�7��&��j4����x�.^�8$��e�S�n���ʿ�g���3��7�t�DM�e���6���,],έ�/"�_�Ow�������_���EP<�f�ï�{`8_�"�3,/-���=t}�-����V�G���i��L[�( �8�"n�\����+$8GknOBۑ�R;�##�|Vt�
��-�f�n*$q<�@IpR�/�=>�����m�Dl�[Bsd�eJP_�)�M���Q75 D�w�]���k=�JHܷJ�dR�=�[<������{���|�iL]@l�R��+�VqXCI6GpH����1�]�Jv$nQּ�g�X�<����N@a3o�t�O�̈ɝ���r0b����9���|8Z4��~y��`�U��P8��J٘R�5얦D/�5��z��O ��H<��P��"�� \)�{�el���و���Ѫ����,�o�y�����{�r+�f�>KOc/�(�l��w�"Z�.�M�n̛^��Ee�뮝����I�a��猙��4�Z'���	K��n4o���y3��� gJ�ݢ�ӳ����c���L�a�o��j_}b��Ҳ!��H����r��ъ-|�b�t9SE�%�sKK��4]Bf�s_�qk�@�S�(����(�	 ���I��"��ׇ3�L�t'��wa1�:{/���ZwH΁��y��\O�ey��Ds��CH�#����u�VV����: ����5����>�v��y�|aC�~j�ÆSH'�am�6K I^��xE��S.T6��r�qj��0�W�d�W� ��@1��i�S�y�2Y�l�k �Q��&˧�fL�G��Ė�u?b�-�1b��2�dre0��^Z��Q|��� ��UZ�9�ܩ�ê;���"O���O嵑;鑎A�@̛7��1NM��C���:G�~�N�?W����Jf����M�B���p�.�m� X�X���5�a�� ��R(ps�k�G��+UFQE�>�.����ZOW�G¸�|Z�40y��_�������K.�co�pD�l>��:�i�>�:���M�R���g�VW�x{��A"?��F�<����J�EU�#��[Ԋ���ubx,#o�o�ـ.�g��4]i��݂�"�0W��}����L�tCkX�S��35FX8��}�p�ٱ��� >�K�!#(�O<���b�i��	һ:R�+��v!}%�;O�Y?�-*�ɻ�\!&�re�o����R���X�"{�en�!%�^��u�yL�ɟI"�t��L������r>� ��\��SWrN��Y$�_�0ź@)���{f��2�Խ#�ڕu��'�v�$,��\TD���4|�=�I���]G��/{��n�a�}9�ſA�f[r��	)a��e�c���͠�WcM����az��p���:���F��VFh)s�x�?��=!�F��-�Wr� T�+�Oh�݁LW��g��c�A���"�����)�I��t�Jc��\��� ��Ck�)�T;@���6Z�nYTH�t�]�>�:��ٜ���d�$��!4�°D ��״�t;��O�4��B+�B��o9`��h�mޑ�FڕP)1_8��"rP���Hf�(/�f����B�.	�E�F�x	GRje���e3̈R���]0G_�I���8r�x��\eI���
������,X�
]��7��Bc��	Q^�x"�N�g�����t
(6��8���j�m���ڣ4��w.���|�[�_��.sZ�
���'�i{cا�(�&}��+q@X�}d]��8�p��%���D�	������J��@\P[��PR�"����BCc,��J����a�%l�&`���}����R�Lv���3���˓��Q���*��!00�L��`i�����'-�ߡ�"	r,��i�\��pqf��S=f|R�#+VQ+��w?����
[�)��p*��2��6�.��5�4:��������H#�&ڋ��O�Z'S�sY�I8���M= �6z+�H,�z�q�8b$�[�����3�5Z��1���C?�18nQ�	�8�؎]`EQiG"�HT�5�������w���LAߵ��w�$����;'~w���F�Ȅ�7;�|�����8&/lUI��&0���x�Ky�(�F�K��;��3]F�R��̕]:
�ҁ�T�R�����8���V�8��M=�
Ã�>�-);z�$k��]�[�hl�����g�2��	�Nn��������>0�z������ai��c Kf��M�w/��&[Zn��`��k!k�'UC�%_�h%nV��,M�ͅ����y�+���)�#@�陚�����yJ�}iIP�5�Q��u<26��K���j Y�������\�0-r����[��ڗ�g��em[�.�9 ���x�r�D�;b#���`���f4�Z��	�J9�Br	-m�j�7������Ee
�L�\�w����ю�Usx��)����m926�78{��SA�{c�e�mT��Ҕ�a�`�,Ú��"�<�4�*=5��=���9�B�ri�G���,�{>'����?!-_eT�ǧ�?�c�RSd��x�p���Ԛ���������i-(R��ؽ55;M���h?Q�� U�4b!���"�Ƈ��~5i(��A�n��EC)��B��j� ���[�Y3)g堼���2��
ۉ��NJ�es@263zA(6�ěo�H�>�x���O�U.�~�c�0~�/
ї��n��O���/8R�$T�ڔ���Eo�T
��|������1X$̚J����dE��=p󪫀1�1XϞ˝k�Ս��Hr"��2�����2�U�Z��H.�YoG�F+��-C0)��Eê����]!֜�!�$�>:lo��1�D�?$�k*�=���e��AL�Z���rQX�Ɣ��~%��z��@����j��Lj�2��Y��Xd�5��%΍���!H���C=d���T��tEw����~ɞ
�_T�E=���ɖ`iTt>[�+����;k@��(���!J����Z���c�T/����E�	���'���|���W`��$f�fv)~�*6 �G�����˵mˋ�`W
�ܬ�w]D�j�M�O�N5
=ɠ�G=&Yɍ���!㏩�>�S`����ɐ�d��cv}��1��]_�I�ܸCIx�2N�E%�"�X��q���4�g4�d��Ĩ7�*����ȽJ�r(��E͡o�P�{�K����ܟ���Hw�j3Ȧ�q�K�rJ��K<sQ����sѧTiV��D�:��_�MHsxY�Q�Oi��V��; ���c��C�t2-������?��"�?��me��R�\0jvvj�t9TC��Լ8��sP�"�T�����x�k����2�c9\�f��zj*���:�����A�:��N�����|vzʷ½:��>�{ȡ*�D2_BE�K�#?�Bg�fZ%k� ��ŭ, �{6磟��na�`�ȴ�.����	s϶���؂�56�����l�YQ�O������M�47t��{�0��`q����o�.\\㞳Y� Ѷ�#�H	�h��Cd
*��y��yI��UGu��}<�ܦ`���8�ttku����*�u��[4���q?R#]8�I�6�C�~;� ����0�+iRT/-ѷ��am������=��i~�}�t���>]t���%#{�?u�R�ft��������Z<�CIO����%т�Ǘ��k�q��yGxr���������}O���7h�z��I�+j�tS�n^1ґ� ��v�c}�T!Z'|��
j� ��l��<B*��.�h,+��� �ƦB3v��U��Ua���KzǶ�+;��I��{o�H(����1J�Y��6^�DtwO�4�2�0j�sU�s����ܘkZ^|�&Ҩ�]�?m�+�7�V��Zz_��.��@�]����Cq�7ӂ��v	vZѣ8���)��|MX�p��-��Vdq��޺nPt�4(��-{��a5!ҌÔ���$�-4����Ra��c�V���$�8�(E�����e�6�&S�5<+� ~�t�����;B�?����:.گ�>�
��MȘ�c�U��ް^������ۊԂ�YW�|�<���&~*]/}C�B��z��c��X�9ڰy_��� ���Su�Y��+!���J�����z�!&�d���>�%m>�QL���u��G|��<�M�m�.>x�h|Y9O<&Y,���+w$ņ��n-�~:HC
G
ip��|@��q��k鋼��85
�7&LC�+��+�'�#b��K�v��bu~@�7����Ch�Җ�գ���i�r������7�~�ɤц�����L�l�-��v���>hT�L��"�0�~�}ΪŨ��k��MЃ��f��}���&N/�1̄��p6i�F�M��������a�è�V>y?�\����rZ_2�Q����m�@9���	��"�jռ�Q[I�\o�SF'�_�X�`�M~GJ;��8�ɣ�	�`E\*���ө*m���ã��(?�BӮ���-��Z�q)dk!į�)������!�?>�G���CU-�s�sos�B�Я���ࡗ�7��<xɑR&ߔ8��%�W'�(�'-g>�mr:P�3�u1.Z�WU4h|�ڭ=�f/�9^�_9���kF�ĺ�4Pnza��@]e�ۡI�Ss<�?����\�F8����Za��,�L�)~�g���w�f��M�t}���^�R��#5{R��]���P���	^�(U��X���c�p�-�e�+�,S�\��EF�c�x���e��H
W޷�f���I]��y�}\0���EZ)������!�{��/������Z�4k�yܘ3�X6�6n��S�&D�1��{O�۟sS���F��b?/������.�{����.�	@����ǭ��6Hx�(+�m���OV��b�i���0\dN
��E#3�V�f /$qB�g���l�@w>V?�nA�vb�#*��;eѺ�Qb�i`|�+M3��^$�N�8�u�no���P�R����{M-q���.ߋʔc�����`b�/S��N�WU/$5���n�fN��S�K�6",S�Wz�8���B�/YƔ�R��BI7�'��Չ��{js[I���
d�Kr?��-f�')r��BA���s+|�%t1�6뚂�]q�[�ͥ�֮��Ը�����-���+�*hS�� ���Q���� �G�wo�v����`fSo���d&���i���3y(d3t���9�`����G��r�GM)G��|IK��p�-X߀����9b���2^E�P��4�[ew��G�/J'X�a^�p���]E��P|<��j�� H�����wX��H�bÛ|���m��&��
�6��Mlc��/�d�GcK��tU25l��,6� !9���@����:�0�z��R�&2:��(@XgXCDy���BO�]��X^��K�"ݺ�S���� �.�|6#�8	D9O�ȡ?ƚ3�z'�s����"ǨjX��=cT�0�,��1�{�i�H�SE��6Ddҹ��I�=�i�Yb�.Y�z��^�Ǥ��ڑJJ]E�,����K�y�/��?�2�4<�Q����������VN�8rj���JjEY:�.�;I*C�H�	�七Ш=��o�ٹ���+D�t��3du�F����7Ⱦ#�V�r���.��F-���t����sc��A�(�j!Uuf!.W�?��8��ߵVke$��v�v�췪Z�_��6���~�Fzә�{�?� �ʴ'۶X�kE]}�\�ڦ���9v�t���ˊxQ޽�������M �w���fe�m�ᅐ8�:����KqrH8�U6��G��`LB��KIj�?���w y���M� ��xc2*�
,27^�P���a�� CKf��ުp�ȸ��� P��ʽ`T�;D,Na��,F�(�u`;�
r���|���>z ����$��ż
/r�^g��Է��ߝ���_��M��D����4G}�8Q�v8�B��4��������\/�a�e���`�j����[�fE��3�L��@Q��v���5�7̲����ݚi�~bK%��|�d��~_`��x��5�P�5l��-��� ��Ƌ��)� h!7f�~Y�����&�?���xpo?�e�Q�z����/���*U�]
#>{	7w���opjD.��e٣1j �xx_u����_�|���\�ۼ���y��}nA�Opr�&!&�@�¤�Ӽ�Y���%D`V����+�?��tt����8��A��"���ӡ��zY��Rr?�@�ˣ�7r��ã�.���U����H�%��q�w�?����W��v�<(23)&�.�ȵ��/���NF_��}n݈��������o�63W3i�(��s-�3�@3,⇿��������@���f@�F��6�n��u䶣�7FIu�~?l*<p�i��NE��>.�UOgQ��2G�j�·���Ě��J.��x�H��}hi-ڌS	-�hX �\Wɂh�;����>f:�{�������d�ikƖ�˜,B��W6� ��7�e�¬���+X'�/�6���Xܨ!,�(Z���7QZuH�+�֩����%�s�X.�Z�̡A���z�Vn�k6�+Õz�k�4_�wA��RK[����[�/���:{q�6�?��A>�f��|.Ck�u� ��2x&���$ ���G�B~����t��vѳk����Ka�w�߉�y�]ߎ\�
�ZK����{��?1Y�K#>7�H��޼Zuױ�U��=g�z�l\�~C�ƫ�� �P����*c��&����z?F5�����۸��l�QcSƾ �a��	�����S��.��E��T�4x��P�Z�3 ����ݐ�Aj�3���JU����C׌�f�k^fT��~ivf\�������0�ɳ�˓$�݊�p�����p���$2�I��}�T�����)'f"��|	�mP��䭐ܹĽΟ�wc�e+���o#l���6�sv����9�9�j|9��ph _ݨ���-JS���b�v��+pW�	���~U�� ?�H"�d�pѡ'���OX�,#�@%	v��U���@�<�I�ZT�j_'����NY�0k��dK6;�;J���!Аrg�o/��J:�A�̱�O�R�{��������1d?t+����^�}J�4���Gge��z��7/�H&:= �:)ϭ퍼���zW��_�?A���jE�G�
��o?�|��&{dz}�fW��{�
�RW�������!��]��7\90z.a�&��X���Kw�E�"�IX�wG�n����¡< ��.m�w.��F������]�B�:z-���7�Z�.5�+C;����(wp$#N��z��x~҈X�c�f��
:Ui��0����GY���/p�L�N�,�R�4В��t$5�x�?�/�{u�����f�`��2�?yf��,�M#+|Pm�+����ы5D_\k���O�|�ckȱ�oٯ��\����z��3v�m�mi��hM#s�<ES���d��{�w�H�E�?��|��B��2 
a����v�����Tn�-�47��P�#n�R��v5�2�D�R����\��OƂ-�]?���s�`d.vxpl�v+����	�<sc
uevj
2">U5��$�`W����˓�ƤI�?X_���w�
������1�~:�!���u&x:���ls7,��~|�� .�LI��;�<���7r�R ����A��L_:���W�(�L!�a9����Y��֠Ny`d�2���jB6�3��x��fֽ�0kBJ_�<yDnצ>v��/��񛵨�j���m�+�W��SVȽ�@���R�gR�G
�L&٣��+����,�Sw��	�ݲ��-6R��򊱇����j�3	�E1,��N �+.�x��06)ʬ��@��	�Zx�t&	������@L���/2��`��߲qG�-H�`��"�Shw�,F9Q*p?G�K*�t�W��gX�aBǦ{�)E��u��_�w;�	ZXf(�|0��L��-t!���I�OL?.�g�U����\
e��Xkag'֓ɰ��e���{�u�x���<���R�,�l��rac�m�,{�B��X˷�6ȁ>Df9�V�KO��q�z�m)ޣ*R�<�n�H��x:G�7�섡��GƘ=B=Y�:�=�������5�pN�Y�S�Q�@D���,2�K�8V;�oBn��̸R҆������ZVX�V�`I��m��~��7;���I�V0����:�>r�{$
<���7@�:Z`�[���T�j���R׈���pq���I����O*�w��9��eR���k�����ؙ���(�{�/���-�9���<.t�5ݴ�2gp��8��c�q���[boR_z��ih{B�M�d�O��=k��e�29	+�)'����Bv�!��Y �l�ml?�|����q�k�0�M_7�;Jm�y�|.�"B.�*���*ʩ��u�t�C��|�gܒ��>��"�QP�"���rO1ḍO"��"es�Jv��> R�m�O*�d����a�[�\�bfV� ̨=��^G<,�?�J� ��#Z�=��͟����[��̷	p/�A�.a��F��낡e8*{�7�#�Ju�����I��{�����Z�\c���#��`8q�hjNC0��J����w��~�e
r*ǂ�MI�KLq��#3���Cċ��u�i����Im�(�0�pp�W������_%�|N��Tݚ]�%�����g	�(��7r�NIׇ�x�hl�t���-iJ����>
51W�Tz�M��J�ۮ��H�v���bD��{!��p>`�AɄi]�^���X�����ڝ�#�N��%nL�~<*A��2��Y�F���j[NU���䊰���[�����I����.���h���M�RW+[~f	X��U�v@k�S���8��ʟ�n���wC���ۊ�}qj;���ީy�F���ӂ�<�B��HA���,�VD�m�\r���H�j]���g��$Y������ Đ�g-B*K�Ϋ<N�,.���&���ض��6�c�}���� ��K[u-�!-���3��N{��s,ME�E�tK9l�@	B�1�P�([K\�Rbj�b(�zf�hPv->�����ؾ'�C�~��m䡯{2��;ͱL��
�k{��L݌\b�.4�A�j��"FN���V��b����4�"�}����;R��l�K�yZԫ��-��
��Ow=���ܲ��}��=�}a�f�2ZNx�f�F�l���ws�13E�vj1y��YW枙�(�g��>Ab�%9��H��
pM&�w$%f�=��@�)s����G�Й{��]�Y�*K���mt֜Gg-���E&��o\�c�9P�՝Lh?�ͅ9Av$_�����^c����I����	�-��Qq�*L8���0(��	����UP�~]	o�e*h���w���C�y2\j+�G���\&ZCͷ�I�a�xH���Q�~�>"tv��'u�?���"�4�W�����"�0P�*;�	JJ	�:�w�S�����Λ��/���_���p��L�5�l}��3Kh����u�jh�uq� �(���I_s����fm3����S$5���'�!Tr�����䈼�aD6$]�a���ȅ�p�!%atm�y{��&.3q� ЀyHN��xvO��ݲ�-+�*K��t�B�r����)��y��>�9^� BXNi/�i�"s��آƖLҏg��uXs"v;��ڕ���<�H��0%E�����=�&����Vnk�.}��m�!e�-�ˣ�?䒊A}�tI�oS{��=��B#գ�A���wߨ5��غP��BD!��"TK9|kĘk?ɥq1���ɔ�Z���qmh.��k(��w#�}��	X�核9%��YuE^�G��F��7)猪:W�6��@&Y+�z1����1�=uBQ̥x��#±�蓖��N�Mj��O�t��3h������?�����쏳�%���lZ�>�r�B�E�M�r����+͒w�-��)��@�Js`yO歓�k�e�f���Oq�l�d����z�ҏ�'��(4���Ow�v��l���
{R'�*����2brqf�m�~�sSzQ����c�[ӑW��ɣ���pneX14��\�M�x��	��,��	�u���};e������7<O<ѻ5����"`�p�ċņ�]0%�S����n����5b��x�1���Ç�B"�0+�
�ӄGI�*#Wi�'�d�^@�>���/P.0��BЁ@�k=�����We��I��_����߼y+�N���X����|}�`�q�j�ǽ��]>'��(mc^�}-� ��/VNXK ���� �tШ>�z;�®Ҽ��p�w�$�����y�[�f�.��!Y 6�P�r���\�6�s�Qpr������Z�X�K���j��Z�T噉�c�x%��qJ�i��������h�ZD��P�`�Y7�]�Y��#n���i�����J���� d�x����r$���؅�b�G��.���e��B����O��w`�x�n��c�N"H��$)[/Ő3�ς	כ}��W�X1�tNT>#���0������V-[7���j`�D�����g��PoB��h�����M��z��<w�X))�$��͏=�)��WL�/�	�0 ���&�h1���b�/�t7��;�"=�ᢈLD��H��>szzc+�i���.�z�	WP�9^R�.q1�*��	[-�% �����:y�Я��6��-���c��x����Ĺ�v�m���E���XtfIb�m�]ƴ��T�i����[f�_h�;Ƣ:_�� Jy3��F"~��p�=�{�(K?�Aǀ����~-��o��O*���B��Ω�I���7
���p�n`��"�zZ�)�H�G�{�k����)وA��I�)m�Xx4��#es��ň��j�mP�c����/m�I�Ӝ�iB�8%K�D˒^O
�A�@�7Ia�5������ӱ;�	#�3	�NN������~W,�N��7\~�.�
�m����4b�X&������ ��@T�aŌ�wv4ay\Q����
sw�����9\�f�����"I�2#{�<�3ڤl?��۽��ڹ�4�qz��[ʓ������u	�GE;
௽s޿! �V�͜_�0Y�	q���bP�^���^����+�3��|��>Q�9Iv��ҬTtX��i��!���7Z�7u6�05�{-H�g�Y���%�� uPq:X�1��*��L��Ћƻ�"���C�`�0�����۳�ޠ)q̣X�15�-����_�I�'z��ȅ2M�	��N�I�������*D�r��!��rD�(~A"��=Js���oX���!ػ�_��g�������.�!9
w������ʱ򺪫BP�Z�Ί��������8�ȜR�a) Z�_�����&f}�}l�*�)!6
�1�}: ��G��#��] �$Aˊ)��O�c8��$?���M\h��葮0��a�g��P�˪�TQ��P`�$df�ؔ�����J�ڠ���Y
�`*��'��^S�2��U�%��FɿT^�9�g���n�V�sa�O�r{�Z�Q�+$�\۱I[�9��dE6ٵI4
���.�Ol�)��9�W�B!��$ϔ��:�:�kn7���m�[�O��f?4�t
5��	:3ӌ�ʏB) OA���'RP�?�mb���=�	�4|��B��p����7w�ٟ|��0�Dl����kg�o�LOݜq!����";���,� ���RA.�d�F�J-�Q��^���z8�Z��,�fو�����4�4�C�V�=������q#.{���5�MiCj��-^�WP�	7f�]��`�
R�o(�c��ܣ�Ў˩�uIx�_�YM���ȏ`�p���2� ��e������1êo�^���$��<�7?*�H�z@��l�W�K��Y��h W�'�6��%���h���j}����!��/`h-���4t�j���+�ֶ\�D�bM���G����R�=V-Wc�\�c9��z�����l�7��j���:���y�?.8�Be5��-��|�S�%3�L���̾��� S����1."-�e�@S���K�H���u2�틘,Yh�����{`�����~L `-r�)Mcn.�z<Px� ��x�"�]X�%�0��!��0$�,n�o4R�ڭ�v'`ґ�:�o�R�~��]�ךM�̟��T1]H���5���[����h�\���c�b�����S�W#��K�� 57�;?� �A!KJC��$��WB���C��^Y��kq�}Om�L����apj�!��5C��c�-�`e�g��Fw��_��kwW�j
܋��|��?(&�o���f��R�e��o�ͧ�[J����H����wY�������ᤨ�HΕK�;&�.�`�5�9�.�*C3�
R��M4\�?��YGl��kr����6|��
3�BZ#%n��m�*�2h��=����_x�	ڷ[k�g˴k��S�]c��	�v�������vl#RݖHg+2�ȸ�]Rbۙ>����j�G@�����ݧ���!�3W�f����v���E�fA���x��>B1tM���G~P�5E��n3#2��k�8��#�e�9�k�/�l�%�0r���H���vZUԼܟtS5��j�Lh�!�� �������� '���"���i�#a5\Q�ퟡ�P�U~`��Q��b�0;�@�Y�Vm_�0U[}��	g��Y'�yMh���?>77T�d�x{���et��'P��{����-��٣�6�@j]��|�mC�"h�a2�A�;���t�+h�A�t'C0 g]B�j�h9��m���	�c+���6���ɬ%q"�>~�&��F��Hѩ�iT�ۈ$�65�����7�-����z
H.�jVT/��5ؖ���&�o3K+�.W���isa���ǥ��|�is�����s�p����P�^.}�p���I���}�� >L��B��?7ɟ��O'U��Mv��X�C��8=$��~��Xƿh����S���yѶ�1'D(APB���^[zL�KS<�qg:�+��|Zߴ��ۖ2r��&��7�Y/yr�2���_�p���d��C�^�W �H�$��w���R�ۋ��r��j���?@��$��,i������[�3��ݣB���>�ɛđ����j�a������]��B��KW�#��5���1 ��ij�)f������[]�B��y�1�|�GW��Z5gq �	\�|���\bր�U۪&���kNh.֬���W���]1u�cQ
�o$���� �K��1YOJ�{��G�?��Ǡ}��a��=+;�́�ߗ2�Gut�3������n�<��L�Y�vm����aΛ�5�PG��J4����3�Z��h���W���͹6�}�s�4���3����d�*�t�yL>�F5XȊ}��"��S5_���;�cZ��x�Ӯ0 F%�fp��<�����'���
S���������D9�Q@i�Ǒ[�	�sI�޸��]�����z��d�On���t%�]�G��xjU�"�`s��L�ʢ��.}��	��<�����Τ%&��lyP�m�
h雰za��e���U���V|�H�,�
H�X�W��Q�&�؎����b��\e���+��lM��pPr8L���i��� /�O{~/V;&w"��ޟr�}r��T�M�xg�Z>Ɍ�Y�ИPu�7]�����{�Zy�u���	5/Z��/G8/@W���o8a'�e����f�C�M�ܫ�:��'��|�s��H��:P��P+a^V)D�n��������=nߺ2��ܑ@��V��b����8�c���8�N[N��ԝ���b���K����r�R��*s.��څ������΢O�ީ��as'���(����p[�&r��@�ˡ�"jM����6Z
�ɷ�
�~�
��k@��j�\K�Փ��ub�.}�VNV"��nd�����m���ٰ�|��%���7l~�[�8��2\�\К�;vA�Q:�� �fd׵�v�r;j������h7pCI Z
�y�=��p��L9�,5`�f�"���/�iM��~�bȥZ���#�⽹�Bz���C�-�e/�'S n~N��	��b�"ΩI�	��S��V�A�ݱ1��-��� 4��cn��JS�����IӾ�ҌM�1<1ԭ�#{�h�f�j]6���u��cS�ز
�q��sɎZ��1|���d���!c�Ѝ߬�l�ڦA�+���=���q���m��:1/�������Ɠwm��du���ͱ��W���TYq�f�~�M�e�VFQ�>V�xP�Ո_;���j����:K<w��غ�j��S`"?"C��a'P�l��,�L�դ�АX,��	�&������D�Ȫ������csS�/�z��kY'�ә�a���{���w�~'�΂���z���bp�֩P�mce_���)��O�9i�*�}��I�:)�1��:����3N���9�����fݞiz���kĝ&�r��}=���>lA-p�$z)s������p�r�ș���yja��C9$���z��籉Bp����Q��7.���(˗���7��p~�[���+R�z�0��V�~��6<�8%�����賠�׌ЉͫY��O�eU��#*�n����s5S�{aN͏Sh���^(/2�.�[��ؐ��j�C��Y���4��xfL�NA�����isu���z�rb�_ҟ��6G���C�:9�\�i�%�*���X�0ߜ�{e"�X�ҭ��Gj%v�&�� b����r[nQ(�� Z�N�b!�5=���i�*e+�eS�Ƙ�Sw���{/����g.sU>%}��Cb��o��K��O��Y	�c�~bN�|2�.$��J���W	�| �gl�:Afb�{!oјG'��?J��
kZ� ,6#�B�#�R�O���QY���cE�m�yJ��Ts���m��/��ͺ���dԷ����#Zo'WA�,.+Ɵ�H�Gz/V�����@C��Pd�ߩ������ɸ4B̺*�O��R���GE�7�j�/\�C���U�8ι����m����6X�w�
��bO�����]�c�J�j�SB��C"��	P���2y4����K�di��
͚;��ԓ���}��{�X|H	���".ڝʗ�RX�l���9�
��ф�Gv��bl��+�s@_��`X�N��� [NB��8^F"��v=9*;���?k���t!�����=�Z���ؿ�F�Ï�#Z)��w.&��YlEZ�h4G+�J3��[BR�%��=������+�;D9O��b�3���W��^v`�r(&ʾTN��B�A���>r��0ge���@��.��Z���"ߩR�%~��|�Q�����%����%�����i|%�G�����J�%�8�����ǭ��C�\^�$r���#]U/�\�n.�La�Ѳ9��+v�`r�ż���<X#�K�#�SZ�ncP- ��Cq�@�g��?�Қӓn�lW�o{?v�B>���Ez�#��|�8��2Ϙ�Ƣ-�l3�4V�r{��4v�>�U,�k��������������[�	���T#m����������)qv�t�P1j�`�*���ǰ�L��aM�:N�ݛ���� V����-��Uƃ��}M�2T���;�X�9��^BP�|�j�L
��E��b�N�h8������u�R�^����n��$����77��f�������$��TC�tt��zs%�2���Nd��rM��@�(f��l�9����_.��b���\�=5�@9��?�r4Q��9:i<f�Sd6�`�,�o�#'�+�����f(�T�2'�=%�OU���ƺv�M !��vZ�H��M�b���:8������6���`E;����E���c��ra A�|sc�w]QH5"�\�����-2��V�h>&�:H���G�lA����*��Q��A^��CK�Fm�t�Ef3P(��o�a��B@a4*�䯋���$�#�]W�<���;�Y��QJM{8�}T,F�����
���(o9�u� PY��O��G�D;;�w��Ӊ�a��_z?\/΋����葾������i1(_�c{Օ\�"�U��ӯ���k�Wc8��CY���dR!�zݪ�ݧ�£��[&2Kd=`aÇ����������Ч�n򤣑����0`j�`Ē�Z��r(����H��]���|�֫��ov
p�,Z���Iy,R�Ԃ>/�c?�R�'�N��Xr@-�1Ǧ|ȯ�ұ7;+���f�o�X�w��E�Q��6�#t�P�7D�V�-ֻ/���խ�	>���{�ߋ��*OV�^�#z-1r69�9) �`�d.�6V�'!�us}�s	#��ay�:d}v�z�n�����l�_�㲭� =.?
��&�qA��T��T�8j�W�M˖�+{���C-���?^�X���vf���P�TS�8�bD��骘�}��p|$v��W���(f�lb!c(�'8y���W򧺲19|�Cb��?
�U؇2��)Ƽ�8QŁ�I�L�"c���;0�VW'����;�Zݲ�
ş��?��m8�����b�oOg~�R��S���x+�s�W}�`M#l�����=7F��۪l�YVB�����`*���d�C\��5�mM����G�6��_x�N�"�w�s�Q�Ht&T5���K��-�@�4�1͗rꭶ��SWfS���A �;<B\Է��}�R}V����Û(%�J*���Ij��b,��˕�k57-��Σ�v���$I�ʏ�t��4��7��)��M4����T�Eb�/}}��d����O�f?�NEɺ��EZ�ێ.�N]�#�M��_�L
�w���)���2�R>�p�?��Az�^����ꏳ�a��ò�]O�*�~�^rf�7J��T�d��)�No��+�K��vtbXf6�_�҇��Nk}v���x���{|mJ`�K����r��=[ڸ�7���&�`}L��� �}��ac6T-r){w�О����7h ���zMyԅ$(���OŚe	Z/��P�S�!D���W���U�:ax��痳V��[�f��Q��nyv;� �xz���w������l��4�x5���!<l�R4ï�!���x�/���E�P���x��"zu��I����6��j�WH�E�GK�_���L�)>���������;�V�J���6 z#���j�O/�)�6y�n��ҽ=hW��'uU�ʐȌ�H1�+�<�/u�F��:��;qB
���4-`��B�^5}���,��P���lN�nЮC�[)'Y����U�t5��8�7�ݳ^��<�U��+\l ?L
ƺ��[�r��4�zv
$C qd�Ɏ����Ǩ~�S���l�"��o�`�q�x,8�:�:�u�H�|���
&g�5BY��]��@��i�%m��Hk|GxY��o�9J�-��.e^a������S6��` C��/r�Ea��Ƭ��8P`g��,��o#��y��g���'��0OyB��S�L]�� ;�6ʊ�P)�ʌѽs��?\�V=�Oϫ����L�-iY
Ty�;K�G��Q���U�l�-~(�Ғ�m����N�-3-�"#sz4A�u�&���gC"�B$wS��h��7p~�s�Ⱦ��WS��p�r9+x(Z����qt�m�x �|?ښ����~E ��[+P�%Xc��L���Aǟ��	U�*����:��騨�������x�7Vٽm@� �H3���i�Z�*mL��;��m_����n|N~�7������7�t�_ ��Pi W�����S?�N�'��,��l�T�$��x�h
x����l������x��A��QK�xuH��֍�T������*{:.�����OD���ޛb��n��u��9AK�_!�
��]����x�r�x�3����&�˵�р#���:�^!�� ��Pj�p��e]?�Lu��֌}��|�m��>GY�X�\k�Z(JP��Mꈁq����S7̈iڠg��Aw��
/lý�6��	޺���B}�*��5�(�f�6�78V
.'vW���&�6p��%S'}1��VĂ{�ʭQV���`�!�H�׀8�ce��]߹�K��8���YĂ,b&F
s���D���{���@W'�uBs������=K
v�MJ����1J��H�&��6m�Jr�-�+E�֍�h�Ke�V*�cc�*�ೈ8t��zު���
�G0�J���u3��zS]��HJ����
ѭ����&gq�8-��ܠ�9#�r�³��}��zX?�3��Z�������Xzy�#���
�������g9ޢ/Vm��k�^3��\*���^�J����{GZ�ES}�=$���C~��VI6�v��\$'�Pj_��OC)o���!�f�&JAb���߱�jA��ըp�) 2=������l�Y	"X���kȌ#$�>T~��Zq�-B�Z>|!���|ܿ��4�&P?]Lnz���1N�*��|ow�X�m��ā����J����T���y�uZzB�W��]�7����H���y9���mc�L,�ﴖP��{�6��)�]R�$r�L��.��q+��w�A$�ne߻G� Ԏ����MgP�:-��sZl�ճ����,��5��#���|�*����,^T0M4^/����p�#?0�D��u�5�pk5z��?���U��
ó;���2�7�t�*70�+'G�AJ'�D�=Hd��A?W��٨���ri�4d}��,���2b):���h��x=62�a�Т��
�}��)���Ԣy�z�,E@���w�l�ބ鄚�J�H� �j�}y��y;��\����\uR��-��������X�H�!��.�
s�s�$�G�|i���܅�a�<>�?�҈�n�,��5dE�r���sU޵����"�e1&�6$4{�Z�wv�����3�:�sӈ�P�Y�f��ǘ�>��@2�n{D��B�G�:�0��r3F��ڸ�d���a�*;������ ��mpT�/æƆ��P��`�3���'�
l���/e���P�����zj/��v�xz�q�2���7�9��ờ��������7�e��8'~��}�5=0��W�~�{-Ks����"^�[�Eҁ�oG�G��kiO�]R�������1��T}>@9�#����	���e뾯��Wx�ib=BgD�WW�$�2L�0��A?�5��� H�HH��>���fɝ���}�fkrP��Qv96���I��C��j��s�Q.��`]�Kr(�:'y����%�N6��)��� �=�v߫�Э�
��۳���\�c����n���A0h�[���D�<�F������u�q������׍G��wo��0�ˬ��}M��:�L���Lj@��i�2V����Hlu��)����ޙq���Mx�,C+��L�=�d�5��_�/H�z\e ���l�,����c�mp9J"�| ��f�L?��#���������K��� jmt��`K}ha��q��wY�Q�Xê'*��F�eD&��6%�BY��nݻ��@�m.�=����/���;NԹ���)�G,9EY�p$��������L)Q�8��B�g^Ā�b�>V���Z�z���UZ`�A��-�MV. ������Ml����������r��8jO���y�.`��H.bC�ut����oa�D��^=�Zl�+L���K�?��s�Ф�b���+�}��
W���mw��\�n���'�s�гyy`�g)5oM���!��[��q3�s���MR�&'�]l��Io���O_Dd�G���~�nl��u]�+�T��5+-^.�׃aj�Ub_�=���/V�x�O��U8*/M�Z ����ӵ�}J2��ƍ���ŠzM�`�ػl�Cq[�s3��$�N9�����[�B���o(H$`�O9*�O)F%�y�����ر������v�ƿ��uh>��Rl�S�'�;h�DM���f��;"O�iG~���gpÃʣ��b���S|����1U�������2XRQ�� bZ�V������k��Ɗ/�2jy-@�rG��m����,;�IY� 4�0y��o�8�?��f!u��P}�%��f�TW$���~��y.�Vgԅ���}��s�BՔ����ɳ�.��K�3ߨ��f�^c�8�����<������Vid�o�(�={��0��3��I?M��6}:*�!��� ;��}���Y��$������Y�=�x�ɧ#ި9X�[�RQ�|� �#���m�cNu�`�rN/����B(�jp}������&n�v��3�۰�A��V7sB�m���#�6h{�B ,��5q|���ZN���tN���:��T�ϥ@��R�`�$���ge�%���0^?�@1X�8����m>{�s*(���y���^E����M<=�I��2�tnQ�)���^�-"&x��?�0�QT�cKi̹�7���Ӭ�@P�xaT��=%|
��Z��/`���6��G=�������Z����u������,/{�ESe1]�~�T��xP����_�Y��F+|�˖�7���cl�?��`L�<�E`r�ɀ�nw/��	�; ���kF����%!)&F�!(�LI3ٻ���A��r����'f�̦�6ALWGZ��K�	Y{�&Ke���Q��i:�b�4)>J�y�(�2���������_���k��)ҙ|D������?�k��k�jn��،���U2�5�X���,�=�;a�Z��3��
�ϝ�զlvG��XT��v
杳bؖ8��92�����~��pE��ԯ�uWY��jf�m��V��AY-W*䉫�9�c��-͛U�&�ӛ���客vJK�r+�ϧ��f#�DC����W�-�z]J��ı9˖M3����n���/IE�n��s;�``^���j�ߩ�#ģ��;�bl��<�7�pD�0��h��	�P�Ya��׈�� 5�����ԋ����i�t�<��Ѣ�Z��]�=|·Z�^��ҏ͒P����w��5�w	$�&�UN�2��Z�X��+���*`�=�F�mڝ����R�=��;�����'�)&�2�Ū_7F�B�I۞}#n����L��Cmz;/�� G��p3Q�Ge���ک��6�u��9��$I� &��r9��۞~¢`յJI�-J1â��6�zړ~!�x�GtW�a�#+�C�=ayAi��v7aç�j&b�⾈	њ8zv����S�=������ �8�4��p�➬�W�x&�W����k�x�7?1g1�۞Y��z�(��5T.�� �D���%t�jK�ݧ,�7�>[���v�/,
	3�D��(��h���v�莉����j�!8��1�81�¿ <��^��hwH�?6E+F��d�'D����$��rC������X��O���6�9�ȲÁwe%7����9d1�Ѕ@)�e�8R����{�o�l�Iw����^�D��Ω����z��X�#��v�:���
���Q��ߪ�<b��@:p�����3�(��CI3��T�砕ۙ�"K�F��)�(��:��b)	��)O��C���g���B#7&�]���:{��N�Ks�aZH��"-����	��*w�"(�H���z���T�_y�9�$��"[fv��Z���Ϸ��'F��C[HU��>_��iJJ���@q�
�Y[S�q�bcݠol�̝�V�;����f��H)�sU毇�I;�T��4;�٥���L�v鶀I�yN�C����q�����M���a� �9'��qp�ʘ�ۼ:��H����Ud��W�m�?�?Tϛ���zno��9�6�C�~woїzi_�MV%]g�`����鄌P}KB�A�W�O���Th����紡�e�%1�+ə;C�!���_����d�]?��B{�.��Z3�(Q����B���6 �:E'�}W������D4Q>Z�<�Rs�1�$f`��
#?��|�p�x�����x\�u��h /�!�8�h 
{��ok��k%����eI�M���3<鴞KDr����&�z�@�3K��l.�A���0�	��,�����Ռu�<>�p@�U+a`1wJ�ߐ,�z�~���<{}�
v�SfH��F ���W�m'���'�4ϒc�������j�KC<4�auN��"���^pё�kV� u�(H�LSh�~���Zќ`͛�~3�܆����2I]�.#n��Ε!�0���r�_VSCV�b>�]g��hfkq������7!Y�7��B	4���D��x�`EE��R�{�ip>|_O�/�����*Q!�?zCzr���+@6qL�7{H�׳�V%�L��V��65�i82|l/�
q��w�[�88��/��N%1�����%6D=A����<�{qt|Z�ep	�5���:�%�@{1EV&�)�I�9#��q���,]Z#k5�|J�J�ac��=�	?�%k|��A� 2�������ϖ.63�B[O�N�7}K%>;�P�����	��WO�x@�&��?�h�ή���!��;[oQ�sr	SN2}%X���������u_��>�;S iӰ����؎l�7V_d9�u��=v_���
Eo�偱�%�k~�؍��NB6D�o��V�}D.ɸ�!��i|�N��|g��'|�.b�R{i��-��~�9/����x;�Ո�+I����2���:���G�Nf��.���Y_j���s�ʍ�/W�[~B������K��׬�������6%�F�T�vo�|W�ȅ#ל�
��K�kxiV�]� �d��V{����6�0�t��
ѥ���3���`5���ݠt ]x��ƥ��?+���q���[i���|�{� �Le��ÿ���\ug�ŋ(�ב_��7Ԫt9��xA�����>T���Q����>.6�g[]@[�j����Çb�5�s�֮��_d�b|�l�v1ڼC��0/S��u-JN�^�E`������,7yq
}��L�g����5܅b��&I�]{_|.P���!+��5�+�8�0����ИB��;�j���x�>�O"R%�h������˫�Un�n�@�b;Z �2s��Y�eAO�o��\�3��.q����P��UK����pdf4�|�1���k@�ҳ|H������V�P�K����� �_ �V%����"�Y���q��~���#��=YB��X�3��A�מ�
�?�2ĆY�o�~$�/�a%9��Y��/B�N�;���}Y���q��t �с�R`�\�ƹ�|���Xx���|����5:��+E��ͼi��/q%qg�f����J��絶`m�@�/!��z�÷�pLGi��v�,�H���:�^{ �E(+�|��/8�k�|(R��)���Hg������8��!c��)���_W�(�(A�[q7���U���+��N��T%�Q<`��_����ے����u 4���=�B�v��5�h4�rAF7�GS�D��W@��)x�ǵ<n�<tz�T OLw.{"Ӥ�C�p�p#��f.Z��(�K��3���\2�<^b�CƯ4"����y  )��X� �/}�`�=�f��tӹ�q߅���\��Bh�F�i�|�5�Yk{E��tmS�;�J�|�������+*��1�L*��u�Aip����� 33��c̼��/��0�#������x��~[PE ���랃(�%]�vV�/�"��#�*�Ի���m��;��\�PW9��I�2�RӒ�&�}�oȾ�����"G���a[i��π�d�d݌c��J�r>�
��B�?��4L�h��5�I���ɲP؛@��S�#��~�Ny�(��lFA�wۆ踳�N*����Ҋ�v�P?�M"2�ٴ������d}E�Ɓi�w��E[%�w)�3�:��i�
�v���(=ų�<A��3;���,>'�j;��C�����q�`�87~���]6w���s�A����b���Nٴ�c�$Sݶ�c$�Uݡ*(8����0�_ִ6��_���K̋��P���6�T腒�p�*9������'�A�2͂�E�c2ԉ���5e�j���@���<�B?�j��o�V/�c�^�h�l%
8�er�Ow�LN�1���\�bݞ"��%�|d~�v�Ԁj埓�)IꞾ�X��TD�D���^c;�q�7S��ba�a��L���
�;�5,�md�v<Q��ȳm�}�f����~��"M0\���e-t�+�u�����?>�1���i��7��ϣ��8�p�qu��!������}��:��Z�78��pL�eo�ר�ܾ��yfj���:�^����D��Q7z�Эm��ڳv�҄9	#�Č��A���G�@n��;����G�;P�Uo�e���Tō-�������$��h��\)̲�`Q��b�{��y7�IȿT0���?����?H�v��ڷar@����g�۲�~�4����G0�����Nx��&�����]s�n�BsCh�-@��t��r������x*Df)9۞�Ɠ��q�����3;��p��K?��g���dda�f��պ~�T"	��P��XR��÷�Z��5Pr5x�Rz�����M =����W<��7;&󢷪\��$���k����v���и���{/�;��-�:m.��K�� �m
�ߵ��J��Ȫ�b㰘�H��7Yq�%��������
��9�s���#���߄�Y�e;�X��Xj�,�F�ye@���f5�t���jB�v�
z��G�#���C���7,�E>ŋwlD����E[-� l�h��ןT����XzG�~7���i�_��-Չ� �z�Cz<�Ӹ��@8��ޤsݵ��)j���a?���@�g�E���w �h̶�{�vؚe�~�~���
�#�N�(0`�텚ޝIS������aR%I�%]X��S6ڶ��c�*�f��~ޒ�t?~�xTe�8�9V�`r}��`���� �빙ê��A6�c� rfU��|����x/f��Wj�pJ�԰t�M̞�g���9_�W|�Z�%�S���������c���
�˿Mp�Z~�;}u5����F�T"o~@��y�#|?�Q�{�yH�0%{���ek�C���uԉ�����I��Kf�one���1K_�i�!w�I��?i[s&��sZ9Sx��R��:�q'r��W��Y�E���D) �{���\��z
.6m=8��3h�C1-�T{�9���f�6��F�,�Jp�����O�����|�v8R�|���@8�'�B�Lj�o�E}2�w` �B���Sm�=�-�&c&F��9F�$(����h�}�"W�0�v�F̲p����6����=+���@�>�T�!�S;�g�/D=E�l'�� "�a^���5�X�w?.̸A���9Y����%��_Ü�=�|�G�}�Q�Y�|���}t�j���A�X�/iѲHg�T���V,ڢ�5o.�<j�����y�\�a�Pu8;�� J�߾
�э°��?�7��m,"3u�n5��{���lI���]��=;RQ�+���������}-���O�7��z�<�n�X_�)��K������%���)�^ݧ�p�I�ctŶ�,�s�tI0�^�c�h�Y2��ȉ`��IVc��/�~Vt�
Q��ⴅ���/�,��e����>ɪ-�	��:��Y^ު�oJ}�\��g����
{�����gz��/��� W�3�Ѹ�K���N��x�xy"`����a-���;��E����[����-:*��t��MH`��4���K���@���>�B^��q�M�IBBK!���x��|o�\"UKFOѡ��&��V����N$f�萫23��E��P�0>L�Cnpk+V�a�����>�����7՗}@���reO��Z������0{\J4�^k_2��4�(�<�x?�-�[�)��p�>P�q�� U(�ë�m��8��,ZV��+D����FC��	���Fg�/ۅV�BZ����������30��=�c�(6�W��6�������k�Ă�D����}�����.9��[��$iU���`HW�[Rx�:�%���6U�ǡ�]F�"WG$��y���?X7�{��z �&`u�xX:՛|�8�����{�,�VaqLь:��~G<9��"2b ���9�,�n8YN�ك9�ָ�G�dXZ�7r�K
����6aF��O&�k�Y��^_���r8�+��C �� ��Y���`	Ґ>�z���$鄵�Bt��9��)��a`�`���d-�`��f�+>���I� �20�e�X������ ��ʡ�Ү���EP��O|����+Z!��I�`��o����$R�
�-�'wTYC�G�2��;������QB9z�H��ޔem��u���|H�t�h\�a�$�#�6ʫ��5vN|'��MǕ�Î����weh@�d��ctM����N ����ʌ�7s�Y��T6�5�����U��m�)�	�d�WB��0��!E{�VF�a*�HT���1�.p�aO������yV'�Gv�z��p�3��E���t��e��6	�����]"|�t����V�z��q��H�V��8U+��2�Y�I����u��T�}�%/�y֎�Vs�����M�m�}�����0���o���-��e��jM�8(��ĭ4ER����Na�HU�S��c�A�#^��$�F|�K�$?fN�ϓȹD�x�4��ָ}p���wˍ�'L�P�Un�!z9F�-���w�VW���Ǥ�{�k���-y��ȃ}�[6�,@+4�Ԏ�x�ɽ�1Ԭ��@j�T?z�ڴ( [@�Q����NY�3��W�̡�Ğz�G�N��ѕ	H��v����xA����a���N"��Sِ�Z�VmC�PO����4��Y�h M��/��������e��+�ئd��Di6_p�����AD[� ��, |�_�&�x/M�eSG�@0��?}븏�����>M���?�k��	F	6r��J�@���Xׯ.�����HA8y�Ju���2�S�'-��ʎ�������<��U�9i�v���O
^�� �cd��������uvLR����񛹲�m��@�U��4��<�Wo� �����n[K��Ɱv�nW#0�z"-$�w�����JƔp�¨]��������� 4o�nн�Z� �R!����8I/kW CBR6��D�5G>�V���~�|L�ē�,<ɩ.��
w�5�����-]Nd��U����Y�bK�"����>� �B�Ɇ@��|;jal��[�A���;`�,zBE���W�z����@v�U�n���}`�Z@KKCOm{	�n���ä�~�H>S�F�7A�`�멧�}�0Tx�}W^+����#�)j0�#���~�qӏrZQ��*�����X�'{JdbZl��X�`��YC���� \��;*	}t�좔72�c��ņ�W�Z*U��1`�|�D�r9���� ��KoWH+*��t3:)	��r�J�bD��M���)�<�Ѝ���AM����0a�Dėy���r[>X��?1`"���MtV�χ����KP,�g�����J͑������22n�#�Z��´��>.����n����g*������/�N���O�\$X�	�S,�a�Yp��x�|Rj�p=�G��_�`��ȍJ-��;T����堩�$�|do�7U�6�8oͩ_fby0l�wn|� Z�@.��ta�2�jy��o@���>��U�_�� qr+Q�<?|�)�e��:��d��T�Brl���
���@��y��k.�-�������
��n��}�,ԯ�8�S�@	%H����d�0~Yz�B�hTH���[7|J��^)��s�!�ŉn�kG���\֤ދ�w��p2��W^�lI@1����&%{?��!'1���6-��iı�ݑ�����*�F=EՑ�-�;�P�A�(Z�~��Z-���;������bF�����'(�j�RG�I��pl���h,��=F}�ѵ�2$��<���� (���S�ͯ���V!����(�V���X�!�~f�e�i�޼�\�h`UO����γ9�@�FdC�v��� �q�p	�'�Z�ӊ;���\���,�X�'��e��P�l?e���������{���h-2�����h@��uo��o%(��fH;��V4�jWy=�)M�|�U���XޜvX�(ЬM`�G�(�!B-�!�O!��J����{�A�������_ǲ+"��=��r%|jO�P�1��ߎ��?b���ҕ�o眳�Q��C���`GG�FW��:Bś�W���8���]�F��R���-v�� �[���h"�@Ń��aJ�l��^�3�x6�����5ӂ+��� 5Vۗ��u�
M:��k5��*���
%�'��