��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�"��F9s�`&���a�oq���F�g�O�]�<ݲ����eCL��D���{�5��8̝DFI��Zp\m|Q��
�}�6C���UnF:<�jΈ�2�����<����sf�k��,jڙ�����2��X��Ss�HL��	�������+g?���N�Ż�����|�v7�{M��VNB
��Rs�゙�Ld\��X�'��R :�J���^�����kMkx�Q���3!P}�e���Z�Y?.�U{�RP	�)��lI{tI(S
7ZF|���[��xU���U;�"i:fǇ`Z�={%�n2�%4���H0n���q�S�]���	�b,�3�k��	ْ��i�ҙ����DkX���"�V�=�+���Qe��)�
	�@�w6�,ܟ��cTK�{���5� .z�a��|7=-Ҿ`�\P"�PL�2ܥ�j7
����_�5�M���e�J�FbK����-���jHBW��h4��rm�c�SCS����D���@�ǵ�≌��Q�sp�n1BC6�;�Pl6lgs��$up�{ ���Hi�T�n�R74�$�R��R|8S9���;����m	H�&Ң�EF�	M�0��VPi.��&�"�W����3�k�o�Z��K�c���Az�"� �>E7�.Fk|#��v8����-�-0�(<Yk��X��23~T�k�!�lG�;���R LTr��r���Y��E�i�!����~��-��2regr����%���z������QO� ��0�>Px���7���	7+�^2Y���K�y[���]5����e�#�a��4<����	O������`��������N��b9��P��j@�%��t�;�B���-���S��C�MR�~P&Ƭ(߯"#4�y�_'E���Gt)SuhҲ�{c�9b�`�&?��^U�_C��O4�/��v�`�k{�s�c��g#	�~w�8c�=/�������ن�ү��3m�(��.�������UY'�Yz6�����;N�5�6Q`������?��U�Mt�wag���n�`]-r?��M�m��Y;���p�3��l���:�/�B�m���Z�E�Y������خ�V����*J����n��nv#�Y�0��m����;k���S:"hh���h͘-�K���ff��W��@�e��p�Zciâv6V�l�<E�Z��RXL�_�A�d����(4_V��%ȷӃ���%�SS���=�H�5�w��wR0
��[8�hG��M�v��ZX]F�D�
5����9���0�0 �Njc�Rx7��W(YM ��f����Q;�Yﴠ��?K��a�K�}��3�/��܆�f}�-eI��SnQ)��J�5+0K3�����xl���,#�	ik����|�9$�G EU���'�����}�����@�K6�
�͆�~��b*4���߱SD-n5�/NĞR�v7N)��N��D�>���n���q[����J����:d&L�p_���ԋ|���6H�C����\x�Ȳ_w��`�����.>��H)Ɲ.�p���<d�u�K�j����?�ēí�G�/�P� �q����GK�L����Z�$��ҤG3+>�#�=c�q|�vFt7/7���^�lK`SBF"o_2�9��[Y8�QD��'9՞ ���`��hx��f��H+c�̋:\P̵jI�=f /�x{���&�M��o@8*�Γ�=���x�>� Cp����<�4�/Lb~�"�ZaL��/i4�.�44�Uvw�mV�� 4�$��lC^c;r1ˇ��U���>�g={ބ��Bމ����DcF%�'�B. bbh��4�dS�����{)�{=��<�n��^��a�UC�_)|���O��æ�����# i����K�#޺r�?��*v�kq�oU:�,8*C@�N�<��8��,�BkW/dsa����9��@`+��&�D��RW��;=_�x9j��Czl{x�Fz8��m|����q�Š02I�VV��'�Ė��b&�LLާٞ��S�'Q�B�Z���Kq4=� "Ɍa��S���cIʝ�{�V��H4��ǰ-�ST����X�Zw˸#����-�3��@
�	S�JXT���O�ɨ>D�|?�����w�5�.1�Zd��Ί=Zx́l�J[j�^�7PV��r����}�W�ҽP@�2��X5��Y�4C *�:bEh��}���^� ����6D��QX���a���~8|R��1�Y5��Ke\t���ω!!�X�=�K;z�m�12?:�%X֠I�ʐ|����I�R��d9e�XS���W�L�!�­Y�X0G���W.A�����R遀��2�mܸ��.	�ߏ�@H�6 �����b��t��*6�.�9S8�T� �[w!�z$�*�$��4y �%�8N��(�=i#$��q`n�K5~���ټ�r�eFB���'�1%��R�nL�ݍ�4�ȹE�?Z\.����;��s��"�,�mK��3/���`���d�]]�f�G���?S�-s<��UJE�	�8�+%	
T<���t6�?���Fs9�(��Bl�*ܠ�9�R���/����@K#_W��W<�0��*G%��v%B�.���̷E(�{1��ɽ��A�ku0,<bk�>�Y��ME�ܹ7��M�*Fu<��0���!O���������_�CQr�7�:���F!��&�=��Y7���Y,f@?%���P1�V�ް���E�0e��JBw�}e8�L�y����>f_����D���!3 M��:��*!�^h �c���-N��g�#��'WK�i]���%���A�i�#�:����;�����������l/p��T��mzT��5L��":cN�bڶ�v5y���Ey�ÙϻD6s�	���5���Y��-�$Q�/�#��ۡ�AtH�&0� �Y�?D����C�A�x��V�׷�07�[2��H�e�d�c�U̩�9�@{^/(��\�A�+C9�7�#��ɰp��Al�������ٺ�&w��f_�6OM�J���^?IZ9��L΄��S��#e-�P9�jo����֍=s��U�,E�K���u���dg�<��ԫP#���jld�q�|�o���g|!�i�6<:�
�Țaa-Y��H���ˮ��;e�b6�þ��ahSs��t.��~h :#�9f�{h��;:9��Vg\�|�J�� Dn3멗��8?�?�9���Rc9�P&�0�~�)��~������,膖�;�qk���E��+5�b�2D9H�p|J�(Dʩ{��$��g�T��a*�@�Z5=R&��}as�An��s{��`�5�힔��D���)G�9R�Oy>8�o�]�Q��*�;���&�F-�����Ay2yd��E{,�o�0�X���u^��U�j4&by��+�S��Cؘ����}��^m
H�v3,���!��"b�M�c���B�[���&��)+6	�6��Y����r�0Cb�\%��z|!_)��?o�s�)���]C(��dG28�& �6�0�4](*�2�>��ƞ(F��,�5Ӥ��4/>�shɢ5ѥ����y��*��v2D�Db�U҂Aɢ��̒H⋇�K,�j��lk��%b<>XVWI^-��f�\����b�Ze��97w�Oax�w鯯�0��A 3e���,LlIT�i���4#�JR�d3#�g~�A��-s��	�dyi�=���
������6�V����Ü�^~�p�T�uD;���噇��c#��C���"I-%�6�ff!�zO8�dh�����U�L���V$�N�,IKf���\.ы������7E���=:��� ������Ca-�8�X�~�yZ����M�u�
f�NO�|R陈!��ѕ�_�F�
x����:&�4ՔI�d�O�l��4���B������3����Z���B�"�|lX�vӈ�v��A�a��Rr-��.�|��B�<�2��K�D2�p�l�e ��t{�� �7��ʛ5t
�CJ<��B��Lf��l��푛x,|�̥�5B#8z�e�<�Ι�{2�@�`F�u݉ ]A��t��6��է�~�^x�ϋ��ٲ���t�a�� �Ɛ��6�La��ϴ��)���5��HW�P-��b�N�7�u�k&"�B��U"8c4ª}Sb�W���9ҖCQ]�\�~1:��L���pJ,��>�˻i�s�ߩR_ҙ4�lM6L| ��u5�B�f�Cە/�z68�����?E"{؝+%��C���?e!L$ ��J �=JW�i,�fg�����@�Ƒ	��R�1t������i{�%5�T�&������#SY�������mz�N�����)��KӚ8��V<Q
�3�U�<�v���[���"#���x+-�N��7�6z�G����?���{�9��Zӷ"��y��j��th��~.̏PY����g�A3�8�]�./n�
����(��Л}��;�.R�j��˄��	��dκ�%�i��](��Cb�>��9}!3��������1-�1�|��qkQ��P�4K<��g������������I��J��	%�-S�'�U�{�n�<+�$�5���۱�~�'��QZz:���v��՘P�8g����)���։���h)C-��)��*�����dD��Wj�xG�
� ���k6��ʌ��D�/hK���ɏDb�OrY��)�Q�|xX�2����7b-��\�B�s���W����V�ohKp�X��?-�^�y���|$+VxUҷ��ķJ��"�Q���O�G�d9��-F5� �-mOn(�fؙ����Ւ����0�=��d��l$���!����|Z4>q=+_�,˗�vؿ�z�[�Ő3�SR�4���"��97_3UU|����b�R��/B�&��-���C��[N�+l�F1:Y� %#B~y��`֫(J6j��Gֵ6���oI�p�s�Q��J�Aa
h;����2}�67=$3ضx��.��c~���BW�c#�Dr��')Jƚ<Se�}���fzrw���tC��>ni�Ѭe̤��Z�@!1.�B��4k�� +ݬY�@���vV��i��4UUYZA�(|���ג��o�&|�Y8�����6O�J ?ٱO��hQ�`��k6�=��G�� �n���Gݒ����1�����^*�/�hlW�k똁�I���p}�y%}��w�s,)`Ļ�F���4? �$�KHD�7b���c7�.�Wc7W�*�g`�'��ٯ�*{���kz��C����0�����Nӧ��S>/{bV|*��1���	���|�?����$%��-ջ=����- �p�^���b[f!B@��tlyۢ�9�� 
"9aw�����Ce�31��P��\M3xIs��A��x�T�n�p�1�����Q0�W��0I�L6����j(6C�����T��f!��)ŢeJ?�9g��ۑ���ӧ��"X�Ӥh�T��L��.���\�,H�x�m(	п#r��A������t���A����]!D��˓\�2xl ��VW(n��T'�9��r�Q�2|��lI��*�cc
�^@��T��{�&-�v�O�6�����O0'j�Ǧg���?�	Vz��\tA�<����j�O}��y�=o��n�S|�2Ѹ�w,tG�œ�-�ԣ��aU"z.����Յ4n8�� &��S<������P,k��K�:?䚞_�p�Z2{5����7&,GC�J����B�HP�X2�����Y/��XC�I^=����^��2r�?E��~
F�C(�V?�'cVdWŢS��W<X0�:��̖z�3�~�yxY�������*�$�G�o���6r�re5jl��75@���}S�"�z`������n@E7�wL��1%�g�
�r [���˧�ZV\�� <�p���?��K&�(��T�b����l�x�����H�<㨍�;㺹�x���*�Χ�1��SVξă7���b����6Uf�,�A
ym!;r�m�k��ҴR�?J����j�~�$N��,#���^"xV�$!*x��F�@�J�k�0�
4����}V��l9Q���x˥��)�w!�n*=bo��r��5h���W$t����X#��fJ#=5iaq�â�e1ΏX�S�aG�r�$��3!Q�(���+4e������w�K�%q�k^Y�c/�����Z��W	-����!�t��$�1���gl\�?��bi��J�x-M��JD��k[l�ׅ@�|�y�*6:��Bnk�xX;X�����8^�q���s��hw� G�ޞ@~͔j�8V�%���sOi���Y�	���<�)����z��3!Ռ%�/�x�wq������k ����T��0�?�O�4ar�kab�.��Ek#�H��<$��;eNϵ�!�����{�X�����~]}%��/s���Yc0��yg$)]�E6S4�>���ô	��
�C7�1��`T.��lo��Ȍ��,�B��۱�Hi���"�Ƌl�^�H	k�&���(���ݐ^JhW�;�2SY�����^e�~��s�lt>��(3]�Ѝ+T��.�/k=_й<�G��V����ܐ^&{(����hJ����eBBk��<����4���^��5�ԊM�k� .yOL�sv�M�l�J���3��5]��Z� v÷�]�i|M\g3�b^1�������`P�"��8CŢ:�RU����aQAc��?Jr�Yru��D�a$ � ��"��V�Y�w6Ir/N��R%�KiT����,��ū��%7�ӡ0�g�Nd��0V[�ݥ�"��V�]Iz���ڵf�����0)�p^��U&L$��7�t������uSsG�/θ�C���"�̙ʄ���*���	���_�{�U���B�v�Y�g��] #l8o���)��Ab�%q1�&��k�Ks��Ƅ�SN�����M����k�_B�Q  j�*M��#N�A⍍�T�NX�z&����"",����{Q�}���"�L��fúV��}�_.D��p�f��>�V.	�(UF�[��Uy#���q���ۇ��:j���Py�R\CyN�r��V�|C�{A�᭖t&��0M�4� ��$��-���c��%�=*�0���ѵOz9�>o;��+sѽ^�w��Ey�{�<Q�0d�����p�.������|���f�EX��J����z�-��͈�4�F_z�Tș�*�q��V��(<9y�h���"nJ�P�H��0��ו��(�8_���'U :�)��S,>���SuݘQP��/����j�<-ɽ�	��`h�S���@�e�'PB�:�Hf8�-���y����;%k� �,�0!��u�f�<����{35J���Z���J�YC��ѣKs�"�u$ˣ^O!�F���	�g#7g��y^��G��c�6����G�<��4hEV�W[�Ic�v�M��nݛ�y~��>��p�{�3�_�az�����e�ת���Q�SY>E�"ƈs��U���O�|S���٦�m�Y�7�|�h�uU>]��TN�#�
���kb�LF{AAٟI��z�O�����yw��J�:pd��R�e��*m�B|��c�i�j�]h{Y�����(�P{�Ë-2��_3���ƭ�Q���X���Gfe���}�-YA���-�=��U�23���t�T2 �\۹-8.�l��W�/�-��-����/H�Ⱈ��;L�4wI�͗f�0�9����7tS�OY_��n�~P�	5 h����!䜐�)2�h��"�Q=#�������CP�>���N���o��A�B(S\�\�
�	�����kO/oӒV`ts�Jf����ݞ�91Ł�ho�<�(���fV�d��Gޓϰ$vq~Ǝ��y7�Y�W'����7Km෍N�g�P���#*b*�<ʬ�B%��v��nt��X<4~�L��¼e=\R��e��}*a���!:�(�U-n��t>]��Vc{6�S����e������͌���)�U�u_�+F���Nc�U��v�%����7XC`;�"���ᦣ�̺rtv��u�v@��K���W$ɱ,�Q^P��p�3�Cmw�E׼�|�?��#���^Ӹ�Z�e���84�nD����9�"����PS���UU0�H��ǚ��	��[�/堺�6������n��}P�~��UD�K�}�t��/}D����Y8�.�q�|�-��7�u|�+Jl��}	�UйQT�R� )!wGN�3|�)\"��z�4��E�+Z|�tтCa���bX���FJW->�V��' ���镀�l(ȟ�Z_���2��;�M?�s�]�t�������λ���I��3�[jjcV{c���o(�}��T�s��:(;�9�fQ����ŚE��@�؆Cib�X�k�n�딮Tl�"|����~�r�=�����cX��}/�;�}Ҳ�!0������<(A�?����>z���w=;��YM����� �mv} 1�(�KAW��w�w^+��*��5���ðG��K��~�������{Sh�^ř��ЇZ>C�	9�;4j��{��N1s��	āJ�;���$5�碤0�(}M$�!�S�����v8��F	��5�#3�M�~��FO��U�ns��GI�Mlk��)��G�a���A}�I���n���&`�KvY���P����`���!aM��!���>��H����ꥦ;��e�uG�98b,���/�|���.����x:��P�
@� �j���C�7���ߏʧt�9(@�vr��o��gT;(�Ay  �f��Xl�u+��?�,��t'�p!}��\5�� ��bԑh$�]�X(�ՙ �G�|��#t���״���%=b89���c�o���W#h���+&9�C�6�=Q�7�I	���V��>+(y��i��cKI�����k�FS_�Dm[J�_��.���e�o�ɞHZ��6#F%�� z����EI>Y������%�_�Y|f/���j�m"Ԑټ�x9������c�����޼p;e��_�2&��<��-�?�C.�H�������A]BףI	tņ�RC�ש��5���5�uk�.��Q��ئë�#]��O��8[2�X��l,��+Βo����'�����������L�o3*k���b�4�F��/��$Md-n��>���G�]ъ������lu��v��tN\w�8�;%��	0�9|ɛL�#���ր�Og�(b��t����>�&�T���"h����_�AA�{�0q��Ȕ��Ł("�ք���/�Z�@�Z*�������JX��a�?���fr��.8�� �g�_B����w�q1�W3��"Lf�[��,��9D�
L��A�柀h�N��eQ9
 +y���p�U#@���҉�l1�h�ܔ�p"�n�|�%2�kAynB�I'8��`>�b�IW�񚚕s�8F�z�	l� ���\�j&|��uf�@�u�# = Jگ��x�"�N�$�}9��X��i#n�%���Z�M���_��tޟ��YChg�	̦|�N܂�����x��I�a�E~�f��?���x(o>n���8N��� ��r�i4�q��F%M3�&�VMm�)��Oj����{�T����Q[p��Ն�6�`�.�t����G�LJ����bpA^�j0��1��+����c߅�C�O�d ә��1}2+�Q�ef�%o�v`=��t�o�(�N0f*v�h��hI�\��@�z�`Pa�!�`��]��7.��SP���&�{�?�	d���TѴ�n�op�P�zw��;1��#x_4h��U�3o�R�iu+��F.�zwaj�!>� �W	�E�r߲
�2��Wi3�ڞ4lH}!�	����o���ݓ�3̱�ފ]�c��9z�q���@/^�w�"�P���U1 !��� BA��Fkj<��}��p/�L�"�ş�-�aSN*���%&��d7r,@���	��;� �=�PR��ru��g�/���õ#��3"e"���4�@�/�,������\B��M#��9?��w�`O�����M�cEOn�K~_��������<��R�7J���T�zIis��ç� ���lp��1�I��n�c>4�d�roH%y鲔���1�_���$���}5Ay��`3��di�y��0�J�&n�
�W�#f|rC��_IשD�'&W`�:��m�:�suo��ݩ�3��Y*�4���`X�9l�ȍ 7�� ����W��I��ֈ��ȴ��n5خSn���4���(�Sv����+��"wD�g�:bm�8�Vn��X�4��LU=0H)��X���z%J,k{��_��]�w���u������䶻��Kő��v��W�5�'̧))�F^�I�Gk��DE�2�y6-������V>�w�['�{=�'�|ŧ����'@:�8�[ֆr��<�Mw�!.6�{[8.�￫Vw��j����/��Tk7�b��G�;�L�.	Q��4�p#~V:�l_�r�Jw]t�dD�[���v'�O�����e~�-�]��[f̿`ey��6C�#,P���X:��CKoݯ(�ł[�u�J
�]<��@���"�0H��7�����B=�h1F�(��t�? �*�xYÊA�d��w�#𼻘��'6i��N�1��bW����f�n�r�Mԛ��qх���R�_��^U.k��F�]�@�pfe瞎�ZW�����e	�;Q������˝����ރ劒n�3�Ak�&;���p��BT�D���1�B�>�b�Q];��'����V��$�D<��^��x�h�̔E�f�	�T��o-K+	�_�lED��sTe�V�����te�zFgPL���%�
%eS=���ea?[�)���Ƒ���� �\����XQ�4�@թP�lR���X��1d����Z���d�h���ȧz��ٙ	�Ń�{^���?x��\��?�,�k7Ň{ Iq��h.��WԪi2��z+�&G�i��ce5zW��y��~�
�"�����E�N<-��tg-�q��k�O�T��0|W=6]�cB��գF����j���^^3fz�2��\�����Y���'r�
�����?>t��8z��=g����%m(D��h��U�ws ϸj��R@E��GkE���
˙�wΔ�PJ�< ������%%�5��~J����5�z��q�+�bu�j���d�U,Udqpʹ�L�#�H/.�xĭ��ߍ�q�܎SR�7�e��ϿA���y�Ӆ��e��]��hy��}����^�+Cl��r����vl�T��V�L�d��+���V
�&{h }��=Y���-@����5���r�v<��9x�s5���b,{#:Xz���Τ�����o�)��O� �tI�+���EK��ը
L�	�7
�B��
�0g&,��nr�ϕ5�(XG.�e�ES�V�~T��&��B� v���Vp�y&��y$��0���B�FG����K��"	z��V��F��b*�벵ۓ"/wj"�q.��t!F�h�۩��y��_��@&�IVh)�!w����)�`�?%G��$�W�����P��m�I�2K;?M�+��� �#+�5�-OP����-��cV{��ER��3N!��WkU�>�J?�%j�B�-�����`�H'I��(�{rJ�� �u�,��ڬ"? ��w���y�x���C�,�/����|Ɏ���G[�G��K'Hnh�x=�k�o���(�����Iww����#R[����X���n)�����5֍ř�@%?�]�"������w��p8�K�ԻF��т�B�<�����!В�����!���O}c1h���/`b���u�DZ�$�q�Ќ����S{���Zh�R�aPAoVQvN�(�_�gAo٫��Z�Fb	�T�[>���|-�{�2n$H/:���V�k�'�vd,�b�������&����(B>&^DA�vD�Ӡ՘ߝ�����(��8�vʬ�!� ����9��RJ5�z��s�P�JF}w�`W��0"�О�z(�ː�&Y�<w�w��ψLLj6 G�1Lo�1�fU±�	Pՙ!���>ϒ��v�j���̅�5"��OS&�����+�,�7K�,_4�B���0��ڵ1ʮ'����"J�{��
Jó(YI�t��u���9@B7|Q�2�rK��c��TC�\�Z�[���~"�g�#H���q-�'�1{�*麷w|��,��z�ccM��R��C��rr/�K�X(|�J��S��d��lc��Z!�fg)�²�%��ٝ�mj5�YRNZ	T�'��H��H��f'vD<N+l��{1�L)�J�d�Jd��#���6����vg�dw��l��t�7@���s���W�;� ���a\շ&S��`�T��w%�i�UPx�' Lr���1��r��n����a�8F΢У�ˤ�,F�i�d���&��}W-ם�����֦�X�~�� JZ�"�@]gIH5�)p�j���]��3Wg*L���Ʉ� �<ŉ�̈t����Q(�a5\�vV~s���C9�e�Yh�4����}����z,��z���o\��ߔt8�bw��q�֢���2>���� !dl� ��T�^�j�(k�j����<���J���w�Y�����Ǣ�c� Y�ҳLB�1q��������-�W�P�V��Y���D.�h��=�e�zZ&g*���=�vh��z��
P�S��1�L��j!DXG@����s�i�5�)k���`�1�:�K�C��}�nS�ԡ��͊�\«j����&A{������A`�!`�����g�g���d/$#fKo�����Y`6̝X�d�})�Z�	/o�nS#�o��]��x) ��GT��^�ɬ�����Y6֥8���ǥ��<�ߎ�ta���GO�`��������_,�_{�cM�؁���� ��ˣ/?2S�p��;Lc�Dǽ�+��\����j�Z�J��� �;w�