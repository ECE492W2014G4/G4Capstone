��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P��v�"<ߞ��&'��k%P碶�R�ӣ�sĞ������FY&��{[��a������ b�Y��8s1�>{+.��H���96�r%�2��+Mwchԇ:HndI,�"d��N�UL�%?^�EH��.3�!�mX�_ ��S5���T��M��a-L�-����R�!�M�-�)|�Yɒc@=f�應@&๓�I+�&�$�����К�W�r���:[�e����=�*}�N?��[�n�����.�k�ԡx��O��^9^��0J�I�`�q0�	�,��:�UJ��q�_j�^�,�I%=�%;�w�s�l����%rWM��֮R��f;Le��?�.�h����TNb|�xyp��TV+xys�K�XE�[�$�Epo���Жю�/�,6�&���0�!z�7a��]�b�����.�:�q�߹UQ���1N�CYh_c%������D���]������2_����6���x��M,ebB�(���b�ႏ-]��m���e�[%`UNi��5Z�?���"`bl����r��`�d�s��=Z΅��D��B�e��lLV�̱��
�-��A����6�YM�S�H�/��}a����s�z�p+y\�;α���!�bnYW�r�d�k׽-�?�3�����;ܷ��x{���� �y����F�*0�G����s︦H���R��*�	�6-,#���[��vl
ps� cro�˝�z_�8n�<E�@͂P����*C�pa���0��?�Z,��1�.n^"GE�x8_+�y�q�,����O)ASij\�V�>�6n��������l��R�b@I�F�ēH�%���:�o�#�Pr��i�V-0\��^|�>����c�Jbe1zeÉ��F0�'lZ9�h�g��0-:���c�Ѧ'�A�?����!���6�8,[ �9�Z`��pn�Mf�PPa�G
�<6<���Q����^��Ȧܕ��������v�8��謰��+��N��ț%��ƃ��o��K��y�!�e(�0�e��{�Z)�$�X�W��%p+I:�iq��x���!���?��?���`��,=��҃�8_�P�]��
�C|�W7���y���w�X'��:Z��k=}"�-���G�$������Dk��@�{�Ib�F�Uo�*;7T�~�JQ�ʓ�G^%9����?a�P�O����0�E��6l���bUUr"�y���¼�Y�ٛ��<P�h���7�ټ~��Om�x�
Ȃ����-��ǟ��%��6�����D��Tce�dF[ ���eU�~Y�|�Գbw�j"7XĊ%,&�0��c}�}�a)�0��4�aT=>�a�����I�����\��qz`Ж��"�!F$�N�N�Ϯk�(.j��j���l�����4��|9H�p#ZA�F�^�_C{ ��Z�M�}�Nc�'��\DH^��z��"���R��R�нO�����i�ߔ��|����-��pI�z�^�h>� ���A�E@&J�<����s���v�Z7B��P�� xPӅB�۟��K.����OCG�Xcu�1��-
�D��F1��"�'����o�`�L�I�;�ۜM��)�O�t0r]T2\ĻחN�@�l(�'7�,E�4K�@o�u�)��̇{�D�&g��A_A�H[tM�-�&��K�9
Ī%���څ "~^� V�Q��	��ҝ~)��E>�<5Lr�$(AP�A�w���6��t)~�g&��E]E
\� �-3S�%���&����t\������J|�����	\cVx�V� ��7i����=��amuJ1U�n/��	���9x�>��/l7��L�a�_2�/>�VPn!z��K����o�+idV!��G���k�[$~�U���� �WW�(>B�4�g	�$yU���.�cL���,���w�ր���<S���l���,:x_�`�5�f`e`	ۂфP�\a�j�b�{��R=Au 0i�Ҟ���;��W��%ڙ�w�t�����qq|�(� �'򈈜�(����+����	ņ�+�e��B2��uU���@�t3�y7��9?�
Ykn���=!͠����d8�t~7��2l�oԿY���6��O��Rv_@�묋�� �[��M]�g�/6�9iDm�=F 9	�;��3K���3���o�^�:t(�u��e9i��=���<nU�4���s�IDA�M�)����D����!��T�yJO�'m�w�b�����+������hνE/9xo[|ѝ�B�}�^���k�2>����j^v�jlg�8*����T��b'ˣ����&��Pbl�0�A%���fxw�|Q���K�/#���Ҡl�V?��/dC	�����Zﬄ��vy�a�q�������?'5�8c�*�O`��	�qs��z�Ɯ��3�("�/�^��\Rt�։7�Xֽ��8>�ŷgB�ճʘ�я8�=�bd��=�g1�����:U����.nt�؆�|L8�h-���,�1�Zs����&C�=$$n�q2�H��h����Oj�[I��M[�.�dА*i O�7*��[�S��B|K�]��}��>�N:���81���x�����W�R�Xg���qr��,O�2]{�辯�G=@q��p�0�����?ƀ*�x�bk{��?�ʺ�/��By��9G#�%����>��1�@��"K;�3K�Q=�B��(�5�~t4�����*������Jk����Ϛ�lZN��,<��v`&_M~��������v�'g�����P����PT�6��,��������=*�M�}��G��ـ�]�J��r����ӱ�[I$��!�$��9�M8��~\+1~�ݾ��X����D�Lx�"�_ˉ,��>��}K���j�����p�i��/h������s�/��,�eC��XY�hrc��^�NےcJ#$��d��dt���Cח׉��4��F���QF��D!L�!U
k�%�Hӱj�)�2��N�S�_������0�OU0�1���6zl���Eh���4�~'OAȀ�KORu��D��ڄ�*ԭ/�n`{{�A9 ;i)�k��Z�+�"=���#E�2߄�"Ք�M[-Σ���zW�AC^�TF` �rh3�5d�q@9��(�3f`���7���<���r�G����8v��4��O���V�X�P��3�����"@��S�VM�����f~A�J��z.!�6��������'Ũx�I�q=:��e���rͳ�R1��!W�PE|�f$ұ1 dP�	����_����Q�I�U5���7���X�N���Ƅ�����p+4��1u>�L�k�%��i�!6b�������x$�ACh�Y��ج�oS�E��қ/,o�p��)Xb����M��Ǭ��� ��ўɥ��TJ�a��Mo����\?z����{����w�I���	8R(� �����������^�8f� �`b�c�u]^�M��{��}u��:rҩ���}²�q�q�s��k0-[˔oL��F��^C���i��HX*N�� ���v+n�.�L����Q%������&�k�3]P��Lts�V�F����Vs�M% �&�P4����ƙ��C��k�\�=ف�S�	lT�����4�)��x��`����T��$�=���,$W*^��P�n�f��n�;&|�}(��(e��C:H�M��޸����>3g��~�ݞ�F)`��O�&��*hx��.�K�E[���)��_޴j
{�=�Sa�:�_ ���Y	�	F��sχ9�=	�w�噜����_�����mLx���ˌkQ���f�KB�ӥ>?d��>;5?�3�c/x�"���T��0hs5rx}��[��^�;y�F�NDЬ�
@Ĩ+���c�)X�Ȗ������m6LLٲ�ț���p��¸�#c������U��U�IE��n����4��xko ���*��������!��t;흒?�Pf'Z �9~ն�м`�/E��oD>�
ӳ�nF��/W:�=��]��$���0���m'T���y�P�ƴ-3���O�t	�b|���IA��x ����$)�I HD���%z�x4�t��=6���T�O�ʔ ��+�u&�-F����XҘ"��sY�L��?�:�B�s��b�����54r�Y�J8s�M^�:�:�"�{*�zT�,4f�e�z�ȍ\����9B}~;�u.r�I�2	=���T �F���#��'�փ�7���-�h�W�<+��o\�T�%�Ɋj[���$��8�gڪ��9������fBl!>��\��B���ֈ$gd�nz	p_��v�鯁��D��� 9���G��3fR�E�#�PT���fZ<���2kюVO��,�V^LJG�Q�LB��/q������;7[��C<&?�3ztM�9�l�L ����z;����|`���p�"s��������a�����q���(Xd�S�� a��|?���H����m\���e�:�Ρ���zKhZ�:X"B�ԣUC�������V�_��l&���ʑX*v�
��h'���7��m�'����8�塆r��o*i�=�f��A]�V�w���.�����q��%EL��o�^]Pk�n�!�0I�3�<J^t,���DU��3��s;���^�,FzU'S�ų��:�(�O��J� ȑ�U���ֱ��q��.��uF}ăX��H&v�7��z��xЯ�i)�����b�I'ƇQo�L�:"�(	M�<&����~�$�o�"�
�_���N��m���� u܃Z���D7�����nB�h`NMt��ݾ��AxnƊ���M1ܖR���[<J���5%��Aq$�L0z�ԅD�Kl	�v1:���A�/��I1�S�)��f+Nz^�/���S��FY�Ɗ�jDg%���Bq�E�o����H|Y�8�?VTM+���^}|�~��C�8��6$�ŧ�F�[p�o�T�7�ƭ���LǟnB�x�������_�ו����R��(�]�#7\f3�&F��NܮVh�ART�f�h����N�#�5pb��]@�Y D^V�oe�m��Ek�/K4H�+ p��D� l��z1]4N-��(�#B�d���*�A�fJlš��dc �r������٬� �&G\�y���	�����ݟ}�)A�=�$� �Ԇfc�YX�j���F|��x�3�����AwM7&��$���E����o�u�v ��Dm�wp]Ӕ,�Q�ON�I>�f�/͉󦽔�iC��ǖ���`�I �
��������~D��Iq�
F�5��P�r��k�]^�t�TXV��A�xth,֛�,B��'j�X�imz)�w�g<��ˍ�i�[�(yD'h`[?�uCH����@��9P;�����>	*s�,h��σ�.�&t��g�iE�#�[^�r8�mJ7�jüy�,/�Mh&j���o.�`3Z����nq%Jgn)�ܧ`ZU=�Ҟ��n�P�v&q.~��
|W.I�Z|��^["�D�xpLfP}�u��,3�=<9����,	v�ƈ�o��h�У���;�h�����_�}��K��+X!��3�$G��� 1��LV.N&����a��&R>��z�r���#��(��.���L�	/������k/'�\�PF��L�T�kʾ�\���j�\�:l���aFr;�.�s�8�X)0mu݃8R�Sn�D���r��=s@S�F��7���G88���Z�zz��e;�C�r��WJ,����K�xA�_}�ö/ɗ�^�5��+�7UƇ���&	���WC9�&�<.7UǓP�b\��W'����E+���~(��ՙ��5� n���;��]�V8����6�����B�R�����^�<v&���q�Sn�{�*ؙQ�z��.SM�Q��[����3W_��GoZ?&��G*��Fl�����P�j�T�M;��jۧ!ƪ��D��>j�
,ĸ-Ehfù��t�M�E�V^�^8��Ȭ�C�������[�.$|��]2��r�I~��_�|{��m��LӼp�^ hW��E�g��q�r;�{;�	�;��3\�Ă7	"^�qt����r�F%�׈~���W�.��D��G_��)ٞ:�pH��҉��x �ү��~%��L����廴�8"�%���1%�d�ͅ��vW��zނQP��G���"��5h���H�~����y�U���Qif|�u��BI�)��5ey��TU���6!����ȋ[��>2Yv��\uV��e�^��A�6�3Z������Y
 Xd���h���|0�(e�E�H�J�KL>�o\^~�?�E��&�l5�s��c��3Y�;W������q����Jlo=Tc\A�v?$*��A�qr�[����r0��$�J6ٳ�'nN�wwz~Dp�N��:El�sL�=�\��$7�Ԯ޳�iT~�S�
�.������__���s�GLY�j���rO=:`�8kvj9ΆoM���l���Z/lCX����䣜A��K�`�^?��f��^�E�ؒ���K��W�X�'M��M̚>�9;��%~�4G�@�Z���
���@,/ȱ=���)��`�Q��7�܊p�wP.A�|C
s�Ƞ"��Q3h@M�`I�Μor���H�}�WL��Wʖ�p
%Ӫ'�����Bi�VzÍ̦/{���ٟ��3��A�)^,h)b�t\>��r�ep��k��-uM�;��YN�F�U
��
��'��Ws��ġ��e-H���ԗ⥦��/[�2��`?P�`���s	��2Ƴ���.$7/�K��K�v9]�1��B�y�cݬ�w�JgN�x0��R�E?r�[�*����	ʱ:=5�4�Ӆ_6������ǈ(���9���q.��[Iޤ��>YK\!��:)�:�U� �;G7t�}��=��L�lX~����:��䇡�w��w�ݘH(��O_��r*�PGvMD��5m-�ʇ�9+@��RU
4�o!�|��+�q��VA�͌��4�diݡ3��'P��^�J��.��H/��� _(�5ܙ��}��H�RU)������Rj�g�P�>�����a4�x�Ik�B�n�a�"6�ȧ���5�`�i2��"�w�չ�5rZ����W²� ���0��6����堞�"p���Ӹ6��N9����}�V��#�����*׬�v\���y��PR�9��Se_$��Jz1��c�x�7�"�DeM�����u�Q+bߛEB�5k�aPL��,ɾ�faρ��Z��� � �4.�y<D����b���l��8z�I.;���P�����βJ�\I�+r�PW!Q����T�F��
�ʲ�}<2~������&�א��C}��4��@p ��h��\S�p�t#@��ޡ}�;�\/���8�ã��G<0g���k���[����T� ���!�����K)+�	��R�oqKS����s���Ic�=E�͗^W����E����xҤswcF ���dotx��Y?����c:�PR>�׾𐶚����,�2���0{�n���)ɠ�(�;��gD�8��9����';7+:~��+�p3�]��o��UH�q��J%y����(�-��bh䌫i��x��I�H_��	$��+���Z�XG�Δkk�#�������P5x�Yk������G�L���L�U�S�TGV]���5G��'q��V�Zd95�����>[���:%�1��X�_�B�M`�\+1wZ�Ҏx��%K1�k��G?�����)�bd�:���	

��X �q�/MZ��x�%<\���c׷��jH�B:o%h�N/y�HA�eB��(n�u�4Q4�b]���B��4�̲��	{�y'АUgl
��av�����8n��P��Թ��0�.c�4��!�#�ׯ�\R���}�?VUS��~��A��']>��ǿ������<�K��G0���BK����N�R�F��3�S^%"L��:<����ʙ�;�&��z��t�ȗ������O
]M��[&�N/�G��J��	��͸�>��P�Mv�"w�X����(ov��O�~Rt쟀�W�ʦ5�?�o�����f�`.�n^��������j�7���YE��ŕZ|Ģ*4��8�`��[��: �*�q��Km�i5�3��@J �-���1$�Q��i���H  ~}ڒ�|����]�a��:����A\ �"�3RN���]��k*۵t�S3�X��c[4����U^k�>�`]���Tǯ+�]�s<���*��c�)���P�Ɠ��{7��J�M�i�j�����,��8o,�p��r��U�����a	MP�t�Fڔ��
�H�������r��Y�Xn��/�>��ap"E�w�=�^0�?ȮoA�&��̞�Rt��1�&tFw��>+Uらy5<s����W�D�J�w��'+X3��H$&�g6���[_j3`%���B:x�ڥ���=F!�%��9ẗ�j�%Ӽyj�M�`j�I��)9�LҤ�R�Aw��ge`���sd�bL޸�@�Lp'Eڳ�\�/OX�������h_-;�&��uX�r��!�;�\edI�
�!A;V����I�X�	�J۠�/v�i�,����͒|��Z����N�ͫ�+"G��->�qZ���`�J���l����!љr���c��o&�>b�^W\vai�m��e4`N+�������x'@#�2�VQ�B�B3��Ue.<�����:��?[�em��=�4�Gdr��V)5w !*/:��\Q�'.�p)jQ�Z���w�����dxۇ4�G<����!䀍��Ax1�}3u(/�����(u�ͮ����*o����a�H{��	1II��y��Zik;:�n����v��|J�1�!A�4L�͐�hʠƲ����0���̨�2�]�ִ"�����כ�<�މ�!���%����f��|d�ZP�� 9EN_�~A�ׂ�o5>KA}��Bj��|0[_��U���xx��A����C��E�Tr������ox�4��F��1s��t�=r���f�r�fyAmL$�\ l�k�o��S��?�͑t�Q"P����Ւ	�ΡZI�(~L�T�0�� ]!q�H���d�=I'����t��Iw��.�lQA�e�cخE�	�h��eE0��v�!�@n�� 	!��v��)'����e^��7Q�Ԥ�sM��P4�i�`'�=�z&��o�c/��?�m���)��C-�Oӏ7�A}7��H!B�wD��>x�?\2�.��4��d��-,��d�G��0,���c�v+��އj�vʒe5�!�*�n��G�B�!��Da�K,��qT�o�1&M����PtÔU��dH��!��.���I�����ֵ�Joq�Y�m�Ô'I�m�ҕ��tAg�R��>��޺Ҩ?�%�eoQs�h�?�i��}Q�A�v�4z�v���9����h��&n����X�儵b4�a�K���r �+,�$Q5GlV3��k���'�c�;�\�P�G���pމ@3�a�3�R��݄א ��_�ݟ��.2"�{��%.឵@�xa�a�^HZ�&�@��$'f�4@3�*nV"�:����?-H�D��kf.�L/���p�!#K�;��*U]�E8�N�;s�WjO�;P�|X�DF��F���]����2�	ٵ�R*[��mL��J�~����aI�~�~�i%*q��������|fxM�b����-_�<�k��$Q�CΒ�yZ�#�*=�w��K�K�ԦB/�z�&nut��B/<�]!͔t}yTф��S��)P��̃���b�M�^Ǒ��0�&�/�����ݺ�ŎaFE%��n�@�Wϼ^�ث�����s!۬3��ƶ�&�`�q-�8K%���|W�[�Ap+oކ����]��}�f�Y�e�9�tc*����p ��@v��o&`&����w����\4�w�i�R��g���V�Y��1�Q�؛��-�d՝�7�v�'��l!kU���4�d!�mg�Z��H�
�	��f9]���*ӊ�K��>���6��Ja���e�!2�L����XNz�^Ѧ�Ŕ��m范�@�ㄒ��ʖw�\�ˮѻ��������<83� �r0CP�,��S��Kݟ
��-���R�TR_�N��;(��&ڜ���5���.��lG���j]ã(B��fG�!���MBk�O.T���Ci���?�œڒ��h\�ѐ5)�p��;�I�)|��g�����:Xi�nө2�=׏+z�_��#{�Cyj8��e1Հp��3ID~��$��4�xʔ��?�}X4j�&����G
�<j�����a�s�J��2Q��^\ڇ%|R!�X��� ���R��;%���W�b��f����	"�����?���(�u̜��cY��(�N%x�'(a���B��Ƅ>6P����H�00�(o���z��Uf�?=�=�nTi6��M[�c�~T��Mk���L"����"�d˥��h��u����O�1{�Q�ئ�)&��Ë��AIo�ļ8�����?�;�T��}qD��RS�/�a�`�E!5�lڰ�|��.a��$Fc]�zj�Y{���(�mQ'�>%XtX�X��hDI�|:�����G_7����5�7�J���C[�Ŀ�U�?$��d��'W3��^`�(
G|�#�B�!��>��=�n��M �Qǖ8=�i�]>�7��W�ߓNSz�Hjf
H%�!�'H2N�vf ۉ�q��:Ւ"�w�3���T�PX'��w�ǟL�J���z�v�W���[�kU�\���2�r���}��[�� z��*_=#K�<�ǋ��Z���#���!���u0��VHq��2ªy�����0?]]���Ӌ�1R��q���/d�ǯ���,����e���_��}C��P���''6��}B��	hq�n�4����jvlV1]�#�g3Gj�t\��Náw�{�i���v���7!�U6��n�G���ݐ(L^
�`-Tg��J�׿�oR�Ľz{$؀FD��R��0�`�>�XV����1tm�2���d������d���m���ު��F��m�3�s����� y?�VY��t&s���� w�Y���! �)�x��cV�1s�������'��ٶ.�טo�&�O�����8������Sh!}�S�n�/�_,�[����$!�
q�t�ݜS�����8ٓ�u����\,��Ħ��@ތ��Z`���-��d�	}�H�h+�����n)I��cM��� ��N66��{�4-��_����]��#����չ�Ƕ�^T�W�ק���$=�%����˅�}9D.Y�l.q� ��@e��|��8x�&��:��!y����I�6�����H����8��v
�`H� !�)(' ʐM%;7�(���.�@R��ׁ�'.il��j`^b;�hm�z"��$��pf�����l=K���#צ��e��'J��!?a�5��:�}��ϟ9���FOHWkK�߷Q�Z�+ٮ�������6y��O�3�=I�f="Œ5����z��Q
T��}Iܭӝ��=?��)i�S�"h�j�������-��G�����o��{B��1k�gݤ]��dr�,�n�_��:��b��������i�
ԡ� /�R���1�
#��Ògm��X�Ʋ�;��-�땫��X��;M@-�"��*�W�^���R�x��U���5�O]EJO�vvmb,��	-���<�'4[�ʫU b�mU0$^���v��o�l(NA�P�Q�+��L�c���'l����Jh\�����x'�*���8����Ĥ�Q�7�&eH���=��T���z�vZ|�Rh��
z��Ҕ�4,��(r�Eɰ�z�7�cu_��{h�V��t@����ٳ+�W�7e��11s~���Jj�(q*�HE���� /k��z��:X ��Ro&N@�����=��n^T�),��q��\�'�<Pe!
}�"�ِ���J��Zk�����g�4���@��VlN��
��=�0ߗf�C�hx��J�b��n���F2��&�<�Y��e�@@����gv�;N��I�A�`��6_C�ΤV�"Vw���G�
��g;�wE�����D~,�m�nx�̓�ʄ�B�ɯ�|Y�J��K�/�a���ź�׾��������JW�n/=��7�a��Z��9B�� )%ߨ9�l(����E�!X�u�z������	4���F���s��q䅥O�;��F)Qw�}7�$�&��	�r8�Cf�*ok|�ܘ
�7�~�����=�dzqlq�E��Z,���N]t=7'�Uꝃ�[W�NG�1gP��L/�9`!����c@�?rܑ���.�BT������#����e��q0�|���d*����4�����1pO�du{���p��YY�_�� �a�h|�������ZyW���^���}��Q�gQ	+��|�PS*�*���ܩ|8����U�`�������c�@G����G]�"�����Ȧƌ�PԖ�h�<�Y����rÙ��P�J-��sY�W;ɂ��I2��,:��{��]�C:;����fBwL��ٱE	��� �u�wuB�
)Fk�K����iPM	����Y��JcW,4�En�m.$y��*iD��.�q!LpY���Q>��~nF����)����c��
0'��4�&i!�p�L��T�h�M�3��Y�M$����zkE��)\�*�x���'�u�M,2�*YU~
��^(�����k�w>��z��Ss`]�7r�e�(�� ק�j#�@��B�P�U�!A �P��kJ�m�
�h�2�����i )��8a�H-(�P�N]�?��ۘ���0�P�gT�;\�yp5̸T��E�U���n<1���� .�3�2بE�j�*�r��X����~�.zÏY�V�öm�E�Pm8L�K�#F�Ɋ�(���	b�[:a��+�G��²�h�Y�]�|`�7�P\�*Ґ�	1�u���>���1-���j)�+�/�|g�d��[�)*c4q��
����aEL����M�����bM�¥���J�Ԓ͡� `a7g{�P?3�6�Z�;.Էpis��J+;y�
G9,:o�?.�I&s+��E#9V�p{z|���#��r�T���y��dэ��6̼���֥�4�u�S��ӹ2`q[��+9�}����J{��AF������dg�UU��L+��.�9t�Yh���~��J�����s�Ef�_>��,�dƁ��jF�^�(�l�8g�֮3�'Oo����S��@��`!�I#�r�kJg-+�ē�Ȳh[��qA/.�_Ф�ԛ�AQ��K�s���0r03�L��ڗ���x녛�h�\ҁ��
��1�f�*{�aAT���Nu�:���E�̒z�[&��̄�i�ُ����3��J�u��J���G�{�CO�jwa��4��s۹�+��2=�9$K��G�c�G\�*
B����'�������J��Ք��k�~�Ù�@��22th����H3��c����"<�R� �/i��֣k�]��ޚq��,!�����M,/&��m����X�Y?V��9uE�d�-76	�o�qh���n��ٿ7�Bi�����g�"�V��3�k
�O��q�q��$}Z$Ås�\�L���Gs�
M+#�Ns�c9&�#H�m�M�3�1��d���BH5�� ���^�X�` �n�sڭ�p��K�:��*W����=����2E*j2�j<�^�����f�K`�$R��V�^��5F����F�제/�bނ:��)�V�}�)����#�ę8��/;Hf�Q���Ϙ�ib\ɛ��d{ h%�>Uz��p=���U��έ�z�G��zg~Zv���Z��GmF��=��6��8���O��˟��1��AyB�jȰ3����%g?��Di��*�>���Ẁ`}Vl=��fSx��(�`\b�CxMg�>��l�����b��� XSE��U]p^��Y6��m��l��B&��V��W��?����[�jD��ͬZzpu�L	5���A�A�b�j%tj�f�J��ޡy�4����.��P��*��Y���R�`+1
r��N�'�N}��_Ǧ�Ь�G<�u���T(}�#�{��$-��s$����`S��B�ZtmH�/����������`�+Bh_�4�"i�''���OkH����u:�I�6��Y}���|M�W�f4���Q��BZb��Xe��HN��u�q��NWD�*mt�o�W�q0�������ґ��z웱a / �����hOϰ�x�{^Z��<�	��i��B���;�Fۑ@����?Cw�A�u��g(��SD��B�D�4AH���[�u��:��/�&��8#�E�-��H�0x	(Ѻ�ur�s���^��~׌k��4#x��8�vX�Pk+z�֭HG����;r��jup����Y,�ӻ�wc�E����D���%�6�F���1�/��U��0�0S[���r��.6HL��35aa��d�h8+�j���ew�]��*IF@�Q����5���m����4��r@�r/� �n��4�ɡ�9*	6�٩����q��H��U����,�Α"��{;ք~�K��o
�[T���վ4��o��3�W���Wc���i�$�=�g��Okܴ.����}�X�]��0�7��da\ApP��-�:��s��J�!nfX�;FNW&�i���v,sⱋ�	/r{�)�U��0�`a8輅�J��0��.{�7���:�t�։_i���o���&�ds�,n�k� ~�P�iA�{����nđo�9�eu�.)'�ss�e��0��j��u�;a ��q)^_,y�9+$�q#ّu�u/ ?�����^̓mS�m�X�7|�~w���.�a7+�IW�X�f�%�%\�o7����Z�ڮ�Ż�����Z��3е�@� ���:�#���<N�4��I?h:�u�V��i�k����5l�<n�Y�e�g����A�v�V���0���R�i֍A��s0�����1뉚�RH*�{x��+_�(]7����U?�:^��o��O�cY���� ��58�5�t84���{�N^�7�GӨ��_���Y�!)�c�if�ݨ�����\Ur��F��Lw�D��j+⌽���VNj�y,+-#B����zP-00l~�ZC/�d�G�O�x�	%�ws��5�
�ÏqP�bp5U�>=��Ṹ�'�0�/��|�r�v
�U���{��m\^�̤9��[�~»�7��3����гd�������#y�u��.�M�OP's��7{	~��p���iL��W�B�~՞���D>X�d*��ts=]�m�k���g5X�BS�&�U�b��L<]`�6���Y�ù�3«{�ի�A/�҄�T����?�!��)VE��z�Zǲ��;�Z��ແc��:����X+����k��6�6�V%.71����	����X��f��%�ؼI�5��J�Z"n�!�{j�A��w�ƈ���5�j�mU,�0�o���΀1適+T!n�ˋk�ExL��H��Y���	���/���ɥ�J�Ʃ<��Q��O��8F�O�t��뙇���^�b����w��'�7p����K�	TO�z\�M�Px=�Dӳ�##~��-�:Cf���2��IT�)��,�����g��A@|[�C�몁`t�9�� +���}��v��bQ�~�s��۟˙t�F-��.�tB��`��3�j���}T�3�Qƍ?�v�+|f߄����J%=�wf�f���`;�4}�N6\�d<|�pk��^-k��S�S�Q����z�N��P�J>��,Z�>�$��McD��m�H�\_/���<�ʁJ.q�$��]� [G;˘� 5p��j�6֯��V�ݡ�]��W�<�A�d�~ёn��x�\�|�$�	sh ����Zl��
�ΒE�ԃ��~��\��A}#����aN�z�y�h+[Ԉ��MEL��M����Z0���e���@}�X�W���E�9r�j��;�n�FY��F��̦�ń4�M��edHߐ���7�ÍgW��vy���� |�*>�l����o/j�0
�����v�˵1��m�(�nB]^<�Q��s��Y��r���6D�w>Vv��=in��i�%�]��p�d�)v�Xjc��ojȈO��D=�2����-��D��,��-�.�(��sс��'�G�ҌLf����Q�`�Q�C��r~E���ô�Ir��g�xBۖ{6�t��o�$��5�O,�iVѬW���5�N�B@L�l%�����G>��Ĉ�����co&Oa/H1��M�'g�>���t�x�3��uzQ�-x}�(���n�j��C��|��P����S01{�$6 �����n���k��q�m�	�ع����n>�$.$kP{�2�=v�D3V����2U��{���Z'\52΋��B��ܣ}#y���[��@��|ŝߩ�+m�j� ����1���Q���eT��85��u��h�~]����'���3E��<�؆x�@T�f�x��QJC��(UN�N��B�6�(�q�s=���1�p�?�[y�Ⱦg׻�78��i�a��4�+�H��3��P&V�t���Ό"���e�>�ZJw��gھ��L�4N&+5��,�#v��%��}x���LbI]1�U��RXd���^g��Jī}�r��Σ߇��Z�`����(�!eT_��6���|iG����R�9ѭ��)�K^��U�W�2��ғ
U� q���d�6�_�P�Gc��t��ߏ��;g��P�@�Ʃ]���:��	� <f���Z
/� A@Q>G�6�zE�I&�=J}4�:��4C;?�1c(m�B�z4!M��"��{(~�#�$]��#d��!"��<�h��t��T ����LB���[�_�ȼBz�ߏ�f�t,M�ڴ�#�&���·D�i���v�{�`P������67��d=tv@���J���!\�l	�9���]�vc�m���v��A:������]	��,�˶�Ȇ=�R�B�ĝ��I��F�)�啷�����u�i����y�f��<��Æ��L�#Ӓ�#��q0(E�7��)���x����h�5dz���0|c��NA��on��>���3��8l�LHkǊ�#��oN�ԍ���ߜ}��P�W�
���rKc±�=;�֎��r���
h��4O���bw�1}��pZ�|�'۝(���̑��?� �ŽȤ(R�lVh�V��� Rn�D�y���eg�Gy� �z��i�ϙ���nYӵ��/2
�U�� ��)骨cTɹ�l�)������Z�ж��E;wO���E'�m�����S��A�%�¨p8$�/6��pU#XT��Xq�_�>ac�gA0X/�')��_��/]l�4>
�M��ډ��Q�|��QX��N���v=�u�� ~TK�L��C�:�&�&��O�~y޾A�K�?������o|����%%pRD�C��t��w'��:H_LD2�=r�_�vR{X��P��8��} ��n��/�3
-pi`������P�
_�jy��'h=?;n�ݩ�D"��8�Cb?س���B>�+b�Ҩc���j0���#
?�R����4�Iw:l��}3�8��F��z+����é$�)y�U�p���P���y�Rg����|���ڶ�Y܄V���#Y��T���m�Stz5邭3̌�'&����g�A���!��~
����`�VM'����.�L(��(�3�����5#��
�<���5�=y��ߩM���;�u4���n����J�+pg"wɣt<�����C����	�Z�6ܴ�3�S_���������޽$����X�(�Z��Q�݄0�%�q�s�Jv吞bTc��E \g�8��'�}k�)�����]"#(�`qbM/4��&5���U:*1���4U���ש��1Z��&*�������Vڏ����~G��4���`�>���C�y�M������XZ౸�a��'�����0���v���Բϔ"���Ԅ(�?��\J��j��O=�x��Ué�R��;��"� �>���D��,�T�'���T^[]����N�.�ˆC����{�hN�\
|�/?�Ī5���n�UVQځ�!�~�JNJ��J��~Q��N,��x����؁.�j`�a�.,Id�t�ls��1�*g�3��A��Uǒ�=g��A� �����w�^H8�?����� �����~m��S�a���j�`��c��$�����QJ�uK^����c�n�%�B�zM����E�!k/��DؖҽR�0 �� �pY|���/������?��ڭ�cp>��������.�7���q�!�A0/fE纇�Z-�6D�B���J�zr���bt2�o��&�I����C�=�V)�ۍ����ԩuYܵ�"�n;�EM�U,	`8A�I!#o��8�l��2E|J�ݸv���~ĚG%.�<֏!Z9X:*�m��#�",���߅�İ���J�g����A�J� �mc�$ɮ�0g*�T1I�=�".Nr?B(Q���kP�'��L��%��q���4!��Bo�T:�%c��|�`:V$�B},rS�}�<��Ѩ�4ֿ�&��*m��R�b�Gr>G��ƕ�ij�kE,0�D��V�L6��<%_���ϧ;� ͢��X E,�O"A�h�r?�3�`��M�i��?��
WZsu.�Y�JuESa��iHjƕ7��`�������,?)�{����Y�b���h�<��_�V<֣sݐ�G�C�d5aTd�oȶ0��}�+zJ�.��x�X/6BZ�?4������KP��8Cw}����9�Oa��笃���a�n讍e���b�0���Cі>;A�-�~ϒ䃣�	��I�"�9~ȳ��9��58���z*��R3A�5����[�!,��`�蕸`:�S�#c�E�KD��||c�0�"�U2���FԷub�,mϵ�5�s�t	�-(b���A��4w�i�z�f]��pZ���!�/���B�����V'а���k|�����#88c	Z9�e����J�o��z�%%�a؆]>�6g�6OsJ��
��кu���7�:��M��]���� ���c���}��L7p���8�7�����&U׺���IP�1va�f;"�e]IU�6#�Ŏ��ـ�&#�X�`X	Q�𛰩8i�τh��-=�D�W!��C�R��)^ai���Կ�i8(ʏW)�j�\}���xG�{�m�C�'-���C̝6o��Xũ^ȶw�D댂��Q�'kIT�Cͼ����Aqa�i�MmRbh*^�G�:�6BxG�T���M�o�{zl�Rǖ@��Bi��&��;s��n9:j�q��.2�yC.�ėL)�u	�����v77��l_[6��f����{1g��!*= �F�|6�v,{�ᒶ#�A�_�]<��A�c����r��IkG&|�J�_�;�X�Sa�:"9_[�9�NW�|��?�Wr���|�ڵ�<m�}1mv7.:o;�a[�Α��1F�:F[�f=�͙��Z0_&����VU=�Vo����:��H����9�Q�V�9S;�(�;�7v�e�C�$�/�����0����~��K���0]�Ą�� �=#z�~����-��������A�a�(�uT`;Ë�����=�rW!w�����N�����}d��U�V>�'���v�Ft������s4Un��.�Ţ�k���BLVtH�T!�<��E�#g�~7�KO�k�%j��q��Pk̫m�y5I�id���� ������fd��H����UjXw��X[�9ߨ}������1�M[�/)���<!��SE]�	3C˵p��Q.�'M�-*xN��E�R�3�褐T Z�'��N��m
���5�0b�Z�WT/�V��1
�W�`(�z_�D=҈ݛ̓r!L�>W�-����`X��,��v��ǂ�4�	#%0��az��,��@I-��u�&��%(E�ݯ��k�J���.5��RLї sn!\R�����%.�b�s���V�Ǿ�y�J�{�����x�(�68g�p��°��#����g���ݔ�֓�&om������!�SoP���$Q&�%-�{PS���x4m�e���]-���Q�^Є��q��j����0�+�k��C����0���rd,-rܰ�!���)4�`RS	��0n�Y����+����/�_�%�z��	��Tʊ��@��7�d�WB�!�$�?�J�/x�o��.g�z&\�W����!&+xe ǎZ>e�L!8ͷ{�E��ٍ���[l���-9�H|̋��z�V �>�L�᤿��` ���k}E
ї�Xj��JBOX&��8?_�;U�=s��%�'8�0�$*��h[jw�O�;C7��p�h@�e��p_k�����>j�e��m	�恟(.��cOF��X�ܗ�ŨTJɿ����A�[ޗ����LE2N�J�����4�qzd�_���uj����;��4ņW�~��oa��%�������\��p��H����h]��FK��x=¸)����;��.6i��T^�d �����~�8O��z���~}9��Uxq�u[-?����M���;�H�V4��E5+�Gh�E�KP�5"�{3^w]94"E:�E��ۧ�U�K�2z��c��3�Ҫ��t��(���jf��"��P��<tu}@rXj������-��v�6�����V�xɔUթ;$}s�:��(y��)-���i���H��kJК�4Mt��?�v��0ŤԢ�P/YޣC�#0�bjv�;��Ll��'gnm�����j���&͞�ı�~i���P���-8�ՍU����Ķ��?iJ��>���[���w'��=~b����h��x"��TCvJn��]�U�����F����״p�!H�����a�׬�H#��G�B'=��nmPL�����mAF)�$а�
ߌ�:Լ��b�d���KY��*�� ��e��MX�MJ4�uoj�i�������Ֆ'�~���c(�.�θ�
,��dϓ��K���;�K����u��F�^?2��}<$���%u�
��7)�d�7z�O���#N�Podc-��I�=�ǧ��_�r�X�6��Y��_.+3�6��2��G}���U�f�	N�vOʑ��6�&n��;�|Iɜd��~{�rW����[�p��MZ`jݸ��:_�hEB���G��#�Zǁ�I5?�l���5@��G�|yg\�aPQ�d�Du��3���ͽ���}��ܺ���޻3e�ُ��~�^��T����.mY%^�	{��c��r����Ts&�H�,�Α�+�ޅ�����'u� rJ�-��Ͱ�B) �����weK�89�isq�j��%�6^T�Oq:!�6�ޚU�|�}��B��.(=��T���_T͟f�{��?H��7�@�*����F1T�݃� �]k�^?��mx�V��A�M��F�ǥ����P���)(� ��1ͱ3��9┣��_����O�Q-�"T�=��i����77���F[�q������د�	����e�S���\GÐ�8*�c�,�uീ�N�'�[
k�����=7�%	��{GqU�$:c��p�=���4�^+v#�QFm?/��t�/u����:$��ݷ}��;mu�e��1�����ݶ9�m���
�{��TAK��_�:�p��[6�X�W�8S�H����F��^���G�-�	����3�����@e�4���̜�Byۅ��Gn���i����+�6�
��;Î�=�}4��� �Ct]W'�Y�ɚNg��G>��J[=��W�W��e�5�+a����g��]\���S��j-֢�1��)�#�ޯh�n�ŏz�ԟ��X��M���{�Sȉ��|[�(��D������J�9�%e�uՇ��I�Xq���GC��5]��i����/*|5�EU��*D��X1���y�{@}�
du��@��ZP�e�������!^E�0���'rWz	!��ݲ�PE��i,���R+�7�Z�L���k�����2��:1OA�C���9�N���~��u��+j?:ە+�c�i�V���[��=R�	���sk��A{)i�U�����gv`i3XH����		,�����uV��%�G����t�S���<l*�Qҥ��v-7b�����h�\�Z!~dw�
/ׂ��?�B	�h���0��
l�C�=\��%�G�C�.�x��]��`x&��z�y'��Z�����qxj��ZВ	r��IX�����E����κ�/vT~�R�	��X���ЅaA��5�s�|�XGX[���|�/J45(��~T���d*d�0̌�V?�vj�ƭ�Bģy�;�bATg�����U'J)wf@I&C��Ŕ�p)��#f#+������l�*=�b���(g=�M�'� �y��)������w ��ь�Y#��g^��J�?Z�#}/��L�Y�c)�9���X�W`�����"R���ڙ�ոR�"�8_�+W�]�?.r�A&��-9L?��q���=dK1w�XŨ�M�a���Y���|5����#O �P��R�f�I��6�LB��q�-��:���/������E���=מL����# ��xh���{`��M��&�%EH0�?rd�l��OJf�Ey���9� O7>�$���g�YNZ�����F�G��(��U�-��<}�6��?X�;��Ί[��gŠ�� nm�8N�L�Fo�(&�"-&t\��lٗ����٥� �*ܢ�u#Ɂ)�4\R�YXVGľ�*���D����F{I,�o��0ǈf��_g���-(��s\g0&�f�D�n1��j�����=�Q�c�"�X�pI��T=�S� `O���<�]��A�[����&R	磌�m$�)5g(C��7=����ߛ��'��S������sc�@�2�m�A��d�IB�~��j���#iD�'B����J�׶����4azk����	^E�0);��JQ+�(���U�<1�
/��[����"=q�x�ۓ���!�x���v
���	-��gc�%�`�.�3Ź�9��(�a��k�T`����*&�2v�`��6f��"��ʿ�{��Y�+�dMsO��	E�ۂ��d0`�8dK/4��M�-p��0$J��%���GV9=Ih�MF�����.6J��;v�L��i��,�J�����Dʇꋙ�ש2q��B@2t���a�h��fDdЄ�w��Mב^bY=���_.|圼G����!l���| w[s�D9�?E�y?�<ԛ�/� ��q'�`Sǃiv*��2O����wt
0 p�8(=���4�k�|�.BSW�?K�N��&��F�;�؈ܥ���U�&]��Nl�f�{�G��k���7�ʚ�z��,��ԝ�V�/�sG��%��W��$:ܰߵ����m"�]w)�f���' "��_��N�d� �\ה,=����5�7dyȣ���� �a��0�@�*n�ʌ���(���a�ئ��m�ݺ�,l���#���=+a��>�1?qJ-�������CE��[�O�&�W?�*	�uT��px�}X����st���j��H}_��1?],}��Z2�X+m��$�;�z#��1�n��Y�'���t:uO��|������h�H�+h{;dB���@�aE��ؼM�p,&�J��?�5��{����캉���P�� E�kJ���ay0�$�A�vYbO=elӊ(N�Q-MhfQ���Z߅�e���m��
���:K�8��-���	D;�p���J�!��L �P��.��1��e�ey2EV���͛m�jƿ��}���a��4�jH���/�/�T��._�J9�\�;�Vh�2kˏ�m\����=ƟM���nƢm�ǯ ��v
���ಢm�)5f��E"v��C����5�)��i�'�HpB��ꜤȄC����0�ԑb����y��]M��i����� ��ߔ]]9Fy���<~�3X�#-Ϲ�W[��;c�#��썎���U�����b����S]YC[3-�Mwu!d
��W���H_���B6����FE��C��>����;��LoƠkGGf.m0gUğRߕ	{?:���XK��Pf-�	��A� zy4d��?c<� ��O����V8yL���PD�`�&Bh� �1�H1�{�*A�5��^��'��o�p�o+��ճU��
�B�eD�Ĩ�y���a�g�sKLXKNN���u������EȌ��uD�]��L�,C:�k^?���@/$��S����{���J�V�<#���i��K�[�ExI�E�`�s�}P��E������*Qgbn
��^����,C�/u^��� ��f �]�~J?�=�T��M����4��-k���
Q
"��C5剡rL3nH�y��E��1P�Z$l�ev����!�v��wEz�k���\ ��n����O��-%of@h�K/� ��G�i'Z�=��Nm�}:���}�(��׫��Aާ-�O`@|���9se�\�(�� �s�cpp5�w�ڹ�xh��NP?	%��.���`e=Y�ҿ�|�$��� �A��?���6Z���
��vU��s�`�a��������k��Iy�~�6Ʊ�� �E)B`�s�űy�Ċ@^���7E�2����6���x�p�(�6x�K4-&e:1�nf�YXr�EþPX��R�;s��]LȎ���2����u���}��hS�;�q��;c;П�q�~���A��� �]N�@��8�Q�p5�ڴ��(h;;�݀���m��Q!�_^̯�58OX�e͐��gh�ZbQ^�Yk�jԩ�&2��B�߈1J~ /�� ���% �L3p�z�E�I�K{r�N��d�k(�X�כ�[=���'k�Xo@_�C�$9�R/N����h���t)�W ��jD׎<��T�`�.'�A�룛`�Y�̕�^��DB�Y2��-������?#J�	������Oy�����}���K�U�zI�C��Sܹmq�W��D4�L7 Q�X���0�a�Sc��>��I�b�?���������C*J��yh��d��ue~��IP��Jp�.IX�T��3��J��������$�˲g��Q�J5���1�1�e4�sP1*a>�n��J���	o���I�9u�˹�(�s]�ի�m�v?Hn�_�<X�q��i���T �,x�C��ag�_`ծdc���ɧ�m�������p�ދj14�Q��;jW�/E�~+��"��qT�㉣̿�����M��[�$y��7+�(�i"��%0c�����j\y�X��,
�:���u�W�*�kq\;�V�*4$u��v���^������7�%�l�gђP6g[G>����-]P�V��cgz����!��;F�oT�����6w���
N*��n�	�͑�Dg��ܣ�_�1T���]�����A}q�K5¦U��r��SrY{칱���@@��*�Ѿ�N��N�aN�}�Aj�a � h��G�ө��p�v���O�W�+$�|�]K�,�4r�@�vYT���	׋��܄ʜ܈X%H�J��:l5:�8[�Ύf.BahVKdR��r�vO�ǜ�/u�T!Vo��6��|o�9���(+f���VY>髀���Y��@"��?<��y�R~��[�C�*O��Ft��\�~����Sp ���k����,�D�P+Ł1z���$3�h�B�uI�D�m���f��hJ�nm��O�f�5���gE�$U-��7�t!��x0k	&�����|�/���c
Ϡ�����#�.��UF�^��T]Lg�E�l����а7��Ɔ�a���v�Ӡ�_���L��w�4�I�[�f'ĚͰ�s��ݕ��kH��H��+v&�Y�=�,���b:?`�AlR2��4D-�7y��$ӁNII}����F���1����ά�����;9}�G����������MD2>k��ku1�������K=a:^;����1O�bN�Ab���B�Ǉ�<ť��dT'������4P,��I��A�75����y��gst91����p�12�/� ��0��;������͟Ǐ�a#��eN�
���q��i������8�V�f~p~�C�6�� ����h8�Ya��ng�w^���G�貒D��l`|�����{�$���eW7q:�F�W#_7�in���<�[^�R2P�I�@�����bM_U4��o	h������@��bB��&���/^�;!�(�5z��{7^��[0`0��!۩X��f$��j�^�q�CQ�Q�I
gA�wQ�"�����+D�����+�ؒ�y9�UAe��T㯇�o��)�z�n�u<+�y`��3��u����j�苇���_�'�܂&9z�&�x��t�?�l�` ���L}Ao�F{��<|ko�J^�#jb=v���ѝ�L��')��tM���j����w{`��e���c�
8Q
��2o��L����H���;E�N�?^��l�V\�*��dB;���p����o�ȉS6WX�q ��2����3���(r�ݙ�*�	{��K�ܻH��ۀ�{���S�0�r������`&��{�Bݳ!��C/�h,v�(.@��
"��ܝ�"H�����<2��n~�I6��ZV�c�}���+�h��)⬕�n�^�8.�hk��+�B���yD֘�3S��3��U�\X�`���V��<�ؑ�������m�$�$>J��V��Dbm�5z���J�!{���Oj,?ń!�N%�r.�]+�U�!y-�4Qy~ъ���G
?Ƣ�‵(�!#K��
rK�P����0 �=?�dZ}�/N������ҰD<5��g�O�Q5:��b�ߘ;1��e�����'�ƸT�M�JX䬨�]�4�
�3�:���'���Y����Jb��mr(k;�E�}�,~9��Gɛ��������/��M0y��lt(��I���{�`�м?O�2:�N��tt8t��~U��<]��t����Z��g+��}DUs���ف��`���T"d�q#x����L��O{��ʆ9��I��B�������\��>*�A��~�������������Ӄ��{"�n���&�g��<�HƷT!
{�qQS6�}%�;�v���ۛ�1�
г�z�͋��Kmnl�'IW�{  ���.���kw����#���CɄ�?2��Y��N��s�2�Y�r���6��p� N�ީ%?a�#}/�QO�еQ�KNv>l5ê�Y&�yj�:��O~�YM�&-h��ń!�9�����"�\:�i�eo~�|�U�	��'1����苴옒�tq��ұ� 1ʎ�Kʽ�@%Lc#����"N�_���1�]�n��&!�1�)ށ@̟A:�<�i�����5���p����(���u�?���=�7\���y7�zyNu�fh�ʅH�4_Vfzh>M?�^�ľ�2��'�|�&<O�� �4g.�,z�����ij���>��Ӿ ��u�g����Ro�t:���G�xG�>h��X�B�oL�V�B�Q7
�㧝tn����Bf��Aɤ�_�H"8W:���d*4�B�
�ՠ���j6�D�K�i��t��+��b%��Ǽ|�eؒ�4 m1Y ����?R�^;�'@�����?�����ep� jH3�ċ_b�,+�vf&�oX́/������3AN�)��3�8�~�VF�����/~]yv�;��o���k��V�	la\<�J�4+��[���h-��;�L�ɑ�Q��
���� ���{4?4���b]	�^,<>������7I������~ϒ��U�XN��r�p�	.�e
@G4�«�eR�U�=��e�R+�6��pvt�gJ�P��N��d�?�d`/j;�hf�w�7:ZkGc�j]c��&ܯ)���~�O��1֌�A}�N�����Ȫa �<`km���KA{�
����˼���<�a8�"�;��	2���6Ve �Yaw2p����8ԘX}L����?7���r�{�=X:$�88C���d�ry�
���={j�J�\���H���\�#0�v,� � ����R��?��ziJ:���4�'�9��i4�j�1��[w^�/�z�,s�`�����Ѥ3�Ws�~�|�� �1����e�&(�\���$L�
>���7�yx���_�.x�&s���Cm�h���5?��
��_X�|��s��<lT���/'�KtƋ�C���
�Z0��WԚ��&�	�Э�c�\�[xP"Q#"`z�{/��H�
*�©�i�z��a�`�w���6��bߣhN�z�>���k14bY�n�ΈV���=��+՜���QNh'��4��#Rz�X�YrW��#��Vb�g�PҕA�<��4m�1S�|�ɒ-����[���Hx��p����,�O341�*E�l�4�v��9�0^>�1����Wa�fV�;,Y���eDf��������T�;
��\8���|�W+ݛ�CR���^&~K�Ay/��$�]N>��+���0�S�C�5�7Γ���"y�7�CR���[�VM�_B���ӥ$)�Ⰽ�3��F��}n�d���Udt_��k���뭴	_xu���o�M�bt���`���Ag�nA�Jn���\ѻ�D1O��l3����?�>��bzY�Z�>���+�����u!4Gp����H�[�\��P�)�ܱ��t^�#�?���:8ӽ&�������`
����s�2v�F.C����  �F!9s����*P���|�d�3�ؠ�#)UV��6�t�#-���Ie��9���/�?4��Ԓ�[�[�oxrG�}$;�+��ޔ�a}�3�6˳�!)Z��L^�:����Dм7F��%6���M"�X��F��7/ _�Z]�b����m�0��+���8�ǉE��Ն	2ս	x�X��n��48��W=h�p���"ü��L)i'{i��&K.�I��;��r�K��3�X�"~�?�Ef����z�I���&�!�4�jR����Т�鵾7�5�̬Ͳ�+�Y�T��{Ǫ�]��L1f�؄��x�oZ��C��K!��ٍ�1�� k�&��jr�)���;s!��=�>��06c�܊�!�L���I4q��e��<��OK3�˴j퉹W�UJ��h�!�O��U�/�T�����6xr����K��ixF�����/����Q>�NC˴r�E�^`���u\�޴T�5�d`Ea@d�G
s�;Vj`�d��1���%=�E�J�A��t�ʰ�~�:|�L^�m�������}�g��8�l�:Ur�ąV�8L���z(8^]�Ӗ��#_�fYe�"��.����;(Ă��յ�\:�%;���<����Q��2�ˎ���ޭ��V{[ŹY��:�����/��L1���h���7�����N��3ɔ�Hr��coү���n���!��� ھ��R�܌z_
�'�`CW脣>���Ͻcj쏴Ҩ������x,�o� �ǐ���Ԗ�(;V�B�p$���w�z��(p̿�����%�կ��ؗƖ1���_�������Pi���3����=����ƛ}Oz��\�;	Oq`��ɲ��ŀ���G�v��'h$��h�r�ą��E���:����0#se^��L�{���k�O{��9./��?��~
�\��v����I��Y�cX�ɱ 7�:P��U�G��9��4����Bs���ǂp���Z���٫<-'*0�>�����t��Є<N�����§j_y�֖K���w����W�a_�]$���~Bl��y�\�<�_l�rn��g��_��oL4���-� �C�3�s����7�?5Q梆JJ�^^Ok0��E0�a,$	��$���a��T/��~�6{5�S�>H�<w},�)w���.�x��t:g-�z�%ʜtБE�N~8�lWm�0T���D ��q��z�iy/>����pq��WE�S�_$�si�wAW�q�y�[�6��0k �6��v�Bo�~t�2�1��K�gW��Rk�	�l�P�p7�����aWr�U��
v� ���=�k҇@��Xٸ������ʍqT FXk�'h��2�n$����T1�gC��X���(�l���*|���Z���!^�?��U��7"��4�/*Yԫ� Z��RP+�T�o����w�gf���u3���Rq�( ��������r�(�������&�����5��H�!Q�<GkyLki�����̭��R<٠�=5�r�J�5���_lp�wR���}��_��:��:��g�����i��퀓��7m	��T�cf�ۭih&�>�iW���_�)��mC�-���{4��թ3�o�����8A�^��+쩷J��o�� Vs>��O<��/������N��_V]��?Fk���B#�hq�(���g�t��I!�̙!�s&�߸�g��l��*D��� x������Q���ꊤ鿎y�d|��
���{0H(�>��>�_xv�?f�A�4�����f����eSj���*�_���#���qI�[,��ˁ���K<�<߼�vG&���w:R�*9���9��$��k��a|&r�*�q�[�dJ�9�eA�c�£��J�O���b��%�l?�>[��t:BBV5���~E�66��V�]��"�S٭C�)&�i��tċWH�M�u[_Y��{F�c=���3f�
�끎@[���Q��:�ߪ��g��MUʔx�F[p*��7��1Q��Dp����:���.ecT�M���4�>T�!{��V4]����4����z#�� 4�J*9Cv>h��"��>�v ��a(B�z@?�Eg�O��g	{,N^_�Eiʧ�M���uU�ۗ�bZ,Q�+i]��ɾ~��h�
�cM ��؜&���
�q��42�Wݿ�"Z�"������Zk����������X�\/��
���`�|oG�zӌ|},+�1��Kׅ�AV�n8�;�hƒ�`�F��$H�����1F@�n�N@�j�0�!9�l)kQ�e����8D�*\�˴�("�
�J{ �:p�7wp�w�������[�'����A����J���}@�]��^c��������\�I!Ƕ���O���ʰ��#Uo�R��Zͼ������!D���8�Y\}썓;��!M'4�6����P��0�:��nn�
f�x�����p�����taJ�>X^���6?ʛ�x2����Mm�p�vk�"�V���r�"�ȏ?�y��
�X�|���	��}u ;�.�! X����cr�J��Ge
;O�@�ᡖ���~�k���Mֆā���>�g�1�-Eξ�ڜVAQ~ fEݟX�:*�v�����%�I�p(��#�:��aVyf��K��R�B���7����{d��K�8��~�tխ#b�m��D#�n�^~B�R�N�C�
�-�O���.v�_����Mc�8>��'a�L�@oD�3.
�u����1��{TzTBt�a���ӹkRjz*�8��`�l�W�o�����r���!g/�>�0���GY��k�X���Tբ��\�Wx*ZL
��؇�_
�y��������n� ��ZKr9z5צ�Ͽ��8;�C�S��.��U������?�A�sK���dDﮦ������X�.J���)�=�F>ro�iǔ�gx;Y�r��U�գ��BB���-3�tkrD|#�yĩ��hanY���cM8ro�{P��6o�^Z�2���Y�1!E�����T�w����Pu�v�����$�xs��_R{��4�[���c��,�*Y�}�V��8�|cz�w�T��;��6�����rӪ�u�d?�o�CJ!:�u���Sh�\ګ��=�5(&'	| u=��l�G�#.4����}mG��pJ[���E սA*/1@�ea�di=Ɨ����$��{�q�F���y����&�V#�g���7h���Ê���mj���cԐ�p��
4�J�g��v���+K?(h��p�e���e���+L���).:G���}�)/���!a�!������K^*��o��< X5�`9�em��K�mq����ػ�/��h7�}?*���N��^A���u��<�P���d7���0��,���9�G
�1��*ǜ^@{]�̴����8B��0�Y �t�<�4e��s�T.Ƿ1�j��_Ҏ]�5e�)7����"Q���F���8�X�m���'�8Yx՞x���]�Yiŉ�y���Ú�0�@�N�D���c
be�ю�e,h`��G�{,�7a�p.����� �iw���1�S�����[Z���Lu��78��U x�Mkߕ����� U�1R��75R]i��dU�Zhs�g�p��Cɷ�=�Z��¤��ʐ������?hP��`-,��j�����Lak��Ig�r��:_!�n���=�@�|��Z�O������QZ�Ek�tc�ϕ����З��k�'�X�[\d��9!�$���gY��5�=�K�HnA��S,ئܒwB�X���?8����d���:㏧RE�Z����`�#3L�۠f��|s��7IW��l3k��fu[y V��� ݛNR��A�),4��a�߹�P�H�нL)�H��'F�w$Z��=N"�18_����R�]��҈�%��r~x����5�4���L��q��νu�ƒ�*����E#�1�e�ʉ�z>��O���x���<_=	��2%�s&���p]
Z]�8p�|��Fn�jG>�N�yn$�LaL��G�eE��扰��o�ط]�S֚�e�$�CM�Q�.���H��ِ8j�C���RtH���'nԪ(d������O>�a?vq�W50��^��r�z�q��n����"� r�s�IN?�mK��ߎcO��p���?��
9t��K�,v���5� �,B�y��EWR��{Hb�=��!��z}��ϩ�b�9�c�r/���%��g��Ǡ�O
�w j��0����«���&k�cZ)����0��rr�f��fH�$�9��yh�`������ku�%<�%m./����0Y���3�+�;�g����k�+��"ÄA͝\�X� ��؟��=�����w���b����HЦ���ķ�Q�	��b~7CE��l�=@4♪����#b��p�Խ�ϣh��3�˜Bn��O�U���]�jg�o�doD?�>w��C;]F�����#���N��Ҡ4?�{ ������y#���7�������A���#�U��ơ�GS�,sJ>j~�z���4&����r_���(T����1�pw�\?:��`��Z�9�&��! ��v��Z��?�sB��	5��y�w��8�]� ���|,�����}�y]�WB��� ț�ӹ�1R9	&uP�$�W��;@�
)�ѯC_H{��/�a*W�u�C]w�Ix��G�o�S�����ڨN����G���j�A�!Q+��+bZD�_D�g��s^��}FVU�ݿ o���h�Iic�>�%k���cou;�|�~����)J`-���)��e6Х�W�޺Sr4^/���WHS.��6�[j�R���}ҼqlRrm�egO!,BU��f6�ǵ�/Үҷ�������'�]�!)�� :���c4΄�-��p�����H��ʯ��n�	�#��>��A��iE�\`���4j�fn6�`>�,�%
r��G�0���DYq
�߮��"�:�ܐⴼ��o5O����%%V���ڽA�	Z3�)��7A5j��v#_}C��ҵ~�\�����
�Pk�t��?�����=u�1&R�k�<Qܭ��'0�wh��[�)fS�a���2T�p��"���񨿞=�:�O��\�F���Ϲ��)��Ⱦ��L�tg�^�*q������\(1�� ��¤�	��x������?�;�Dp�,ݭIsa���F���,(�7�̱��<�ې�l4-�(OuYEp�?]������.��������N��̡�m��d������ɚ���3+�p��yWΒ����A�$�u�Ruf��J�	�J�K��˟�\��78�jf�u�Թ�h���Ѫ���j)~{Թ��K�V���w���1?��kU��A��;�ǖ#��A&K�
Sΐi�RU=�@�'^ �ǚ+����6��������'/"|��s���YwI*V��\��5��a(I���p��mp�1g�2f�FI��F�[K7%e��9���g�0n"=I��ŋ�k��+�����<�����y��i��ňy��F����P�+Ɗ�7��x!.Z �6��鮄r�9��Io�d�O��'\O\xl�Z8�A�F���y�B4 �UP���TÁ-��%�����������x\s5��U^���	/g�#��f�'�R�fi̽��a��gG�%�y��������@˫l�h��*V�\�E����s��R�5[dK�D���Iɔ9��k��?��g�:���tiL�F(g�`��5�PY�,8��zR~��ƞ�?�c}�����?�<lR���IKs��9���B(6d�.k�(j6�%�3��^4�׿N�w�����է�J\k��m�|Q�?�<����@���a����0��^��#����O��3Fo��w� ��{�m ��9��ꢣ�U_�k�MW���0�s�5�˙���7˒ɱgڛ��7�����B�}Kt@����"qa�̖�j�JI�6�����9%��҉�I.dΫ}��II�6R���<�nO��]�l��ۉ�%9�b>5x����K�梔�q��KƧ҂��\�e���Od�]iw���_�߹gc�Ւ��/�`\E���� ��n�9��^4�"�_���Ք���s�펤�bi��:���#w8�fo� -�`h�����=�r� )�;�A�ph���'������ J8�C�D��ώ�t�L*5�0IG�G�3I�D�w�&����KX���hL��\�����Gܩ
_$��ʒm�.���aoؽF"&�D>'�������&xOw#�"q1����n���U;���L���k�c6k:F7.5I���J��@��c��veX�/{�zob��ށ]�z�R��_�/Pb@�H�V�31���+454Gp}t�߾�:���՟8c�J���;'y:؆��ƞδI.�Hpdᐈ�����''𚺳���Ð�[5㷓� �\Ԉ��.:ɚ�X#�h�nd���<���nD����� �VcO+F��]ɑ�T���w>U��z�i�CM�z��M�v�X@j%\*�N��@~�4 �d�Po�������S wpʘo�3+�y����PN��@�l�O��r�-����W������^d	r������e�vp4��t���OC*rF��TqJ�U�aMԮp��+��*� N�*����Uܠ@�v����
�(�3."�����<�H>�&$I~�.�=����P��Bż9K!�e��κ�K*�\_�0�3(�{T�P;%�?�M3c2T��8#n���aE��/��Y���<Ϋ�L�B&���[�6e���6����l�Q+�2�+��Fk�[+�kxӸL��� '��u�v#�n!w���� ���i�oM�±͟��rC�S��g�S������I-�y�Z��j5�`p�HS��:m���&�[&A�	ZF���o�{~R��ʒ\N����p��H�)��9���Ol����eQ�� �3CuΛ���o�r��9����d�����Q�|�R��N_�tbKǔc�%�AI�	�����i[�
}$���W�:�����@�iS�ԙ>l�G�kX�n�j�TӆW�x�C��CҼ(r.$��l ����o4|�
��(���'�'&�]� a��~��na��3PD�>��xf�'c�=fP�];�F���Rs�M����#}�Y�wGm�۟�*xR8��F5��1Q�1f'v�-�Ek��1@�J-�D�|{8��q4�J� �F��{�}�Þ
m�L�w������X��;dw)_��&62��:�@����HT��׹�q���)���K�%C}�
��a�3 �E�ڜe*�ے�/�����S�8v`�x���9��[�aq�N���I�c���[�\�[:��y���.(���c?��vH#\k:�B�uG�	���X�I|-�Io�����_�!g>�Au�gIT��ëd����5c��h���S��A���"mdL ��uI|�2�m<_�O�5����K����.8�[Ml���U_�d�������9�O�T�hf��F�[3�n���1��䐣Y��p�\���ޗ�z�:�ݓ��R(}��ɵ@����(��J�s�j�j(I�홧���I1Nc���m.�T����LT_E�a�1\��ۇ́���s;S�MW�bx�PDU����g�+O �ǩ��-ފѿH��K����pi�Ke���H\E�Bm�}��g���Q�N�H�z�r͟�Z������Q��Lφr���K�'�H�N�g�ΗoU/���	Ǣ��f�l2��q묮�aJ�הQ��=I�W$�
w]1�䞧EA�𮓁��qI�"~&���'y�i�[��7�z�H��#�Lj�.� 5kWi� ��M�J^���V�5��3zR` h�lK��� �yŲ}�'�n�%�u<�LU��$xt�܋�T��@��Aq�L?�ȡ���^{Z��p��:|�C ��Q�ř���h�)׺4���<a�g�y<�Y�򙉵�Ș�HCYcu�ۅ�0C}�ƃ��Z�����C���́}}3�¦V���_���s���H�`�p|[�A.�湪�@g{�5���*�#+4���������#�
��A���7��x�"zѼA$a��xe��e۸��Hw�����n耈�}6�����@�6Gh��Kdۯ����ɬH�m�����_�hL��ڇ�S%Vx���N��[?Ԛ���hx���sB�/���	�����+n�DKЙ[|��a� ��"o�Hي���y�����3!������qo�<�(㔶���(���σ�R;]�u��q�a���[*6Wy�B/�M$P��|f x��Ұ)kI7��3���b3���+ju�K��_��lEĊ�	�zE��>��dF����i���W͞����<;�6pVPH�}Ǘ3�Yx�N�k���b��"k�,Mw��B�D+���`��kY�u7۽��h�� �,_�6�m��R��RC�3��	���\�8Лne�#Z
yl*�A��J�'���'����nV�f������$v�>��$�ʰ>y��h�ݭ&D[w&7���6]���*�) �SR��9�=OL�ҭ���gX
��T7�Q|P�P|_C�J�R|LRJMp�{�����k�4Z���"'�A]��-#�,�K��T��=��GUA��)r��z�^ŵ?���}��6��j]Y��g�Ë��fФ�B�l��-��X�gG�����T��VI̯}�b���,�Ŧ"�!:x�?(���T}	�t�	ج�`�B/��͌�'!̚��I�&�#Y
�7 �����Vg^�@�̘���U����(sf;��g���IV�3ЬM��A�d<��EgnʭFĬz6�~�k�V^���o���J|�?�f&UK�6�h�'����9�l$����A�T9@�m��~�Y~�ѥ*�à�?�ej��F�$�a�����ز�9&�Sy�c �>�
>��e������&B��O��CW@$�$"8�4t<p�o��l��I>��{�~_K����F�]u_*w��WP:m�-^�����s<��|X�}el�x�a�H��a�Nw�n,a��"�@n�P��6ӡ��m#^ʊ�s�rl���P����>���#]?�Π�%�4ӌ���y-�q��Z�Q�FK���]D�����zLwT����g�Z�[}��#�l΃'�j�/����������/B�G��IU��R��*٨z9����Ώ�k<�YE2|�O��%޻zH�\�?�	�����+Bpo�D���0"��R�F�H���e�-�����#��9�4�[ڟ��z��'�4�8����WfWd�����2��M(k�dv�n����r@z+����9�NZN#����g*�sm38���Z�rlZ�Py�$W[{�'�w&���Qf���T�{]�7��X�#�����l,��W�:0=��@�����~���O����}��z.�)T���\�T��k�Fp�T|�3y�����܉xʄI5ڊվ�(5��h|q���9�+�*,��I3w_a��T�x�~ñ�q�/[�e���d��3P�I��g����1R�y��WJ"r�"�Km�ل����'��\ӝ	J���
��?�1xc3���`%.#5/�Ѱ�9�ժ���{������K$L��h��	Z�ȳ�Sw�P�Yd��-�C�q蓱\\r�&݇�p��Me��0�{|��Ui�P�����L�8�9r{RY��k�cs0,����2���d�����������m5o�ét
�w�{_��J��Íi��]���%�Y=�<9������\^D�H�/���	�ۦ2qM�9 u�(ۉO�`��J)p͆lEm�XZ�0�}xzj���F�4 �{�d�����z�����tM2>�0��N�CA<��/��~����Y��ҝZ����౹���-rƍՀ͖ׯ��o�R���C�Üֈρ8���k�ᗁA��B�{�N;�����׀��!^���7N���=$kU=��I0�_4�>�X�����Oe��ָ,j��]��-���.���S���=3�����]��9�H+��V�/O�7�@�� �AҬaCC>����5�Df&��`\y����cHט�d�kv�R%z�":��~���
�4���k��$�?�gm�5"T���^�����~u0Ѭy��c-l)���N[�U߿���w�&�m�vP�_�q�aA�eV��ؓ�޹d(W���Ҏ���~�QY��,Ŋ�Er�1�9��\�5��`a:�5mZ��A�T)m����T�,���<wh'���}2��Ч�ǐI��Hk����\�W�[�sׄ5IsfÝ"ް�[��k�Jm�b��E)O�͝��oI���������=
ι�9W;`�=x4��i��F��=�I=}�M��}ɣv8��Z*��.��n���6���㽱�{/	��Ǘ����;y���k�0\V��r�V.!�`/ѓ���۔;aI��ޫ"Nsf86�{F>�����oBÁZJ�q����|��q����!œ�v�)�n�h�y^��5�m���; ,�&b[toe��U���/�N�1�渚̒RpXD�#�	z�B�䔹�54^��Ԥ�wʽb\`Ϭ�e��U�alaǤ�dcc_��͆/C	m)�Mʑ�'�ʒ˹�X@� ���l:��?�l!�����o[[�Z30��{��*��e��x[di��yE>�.����}����R��LnVg�^�|`�n��K&�:�O:2/�����,mH*��M�d����Aҝ�eR2�qrG;v��B2l
��Iv�EͽZuX^C&�򴮶���r���]���W^=�'|Dx�P}�u��Z�k9Fm�����pM��7�+�$���#�H�6	�p\ƺ���Ke�����9Eo�[����h��ʵ��	��&�o�6_�RL�A���Xe�V�*�#�m�{��}���a�w���RcHx��M���m��˨�B۹oq�O}���U�`�����E�}W��?Km���hh�3�߆�,�G>�go�9,!�7i�8�}��wU�+ٴ+�Ĕњg[���?h"����"�9���������:ݎ�`[0璾����9�AZ^�/��T5��������)F�]ƒ������R�!�k����N����������-��K�q,�F"5�;�¦T�����m�5mX�L��9���.!Iw�	�/��bz����g&�n	�b��m�'��j����ϐ8�s���RzqB����z2��]��z_�ݎ��//*�B�=)�2�}�К �m$4MQr�
��W+�Q��>]jB�z;�G1{7;MR�v�(����n5���&m���b��[)����,ٙ��*�6�U�	��0fN1./p�a��<��Oi�mq��Y7�}���yc�6�Tha�1�}Lp�bȝ9%���3"�]�G�N��֦�D�
�exB�*����C�98\�+�9���1������@1o^��p���R|�G��4�Zض���B��� ��I���k�b�EB�)���]�X�&�6�"����yώd��	����˝��٧���Q��ݺ%w�AvD�-�W�P��S+�z���#L'�̂��ɻ*�Dr�������Bˉ��8Sig{�f�T�vlB�O`}�u���JQZ>txz�U${)!1��Y�er�V�_Qs����E����x���T.!�}�4�(:q������P"�3}l͊0E§W��H�N�t%��hl0���yW�j)f�H�8m,�$M��D�a��8�pX������ľϝ��B��1�ov��<ƓG�E9w��`'�kO�,�;v�r%�r�@>A~�^�	�17yDgkڣ��O�H���KQ�����yh�Me���e~a��<n�V��|��Y֖њY��8	�Ã1���h ��؇�G����pK����վ�":�slVM��'���l;Vo�ҋKa���h�Qz�F�-T�S��[ln�?z��lX��!���k�cI}���6��:uȧ4�Hĥ���֝�"��I���=Y㰾}ģ.L�#���.�;f�4Y�����1c�RLm������s��V�J�����x�:�v8���mT�a�S(-�۹��Ĕ�(��ܴ�����/��8%Z� �����t�'@�R��+h�o-4��:����9��f�-���AJB��|؆Q)8�
�t.i�Le�-�0�;�F�g�Zm����h������hs�<虷ڋ�&�aE������pt<��[��L�b6��޳H�K�0����)0d�kV��	�O�҂k����G٫������l#8���Xe�E���'�_��fJ���ڪy7QEwң���=��Z��o���f������tֵ�`/@���lF���}�c�l�"�z�W�.�d�v�,�=�@�0�u��{���������&��5�&L�/ĪD�����V�(��B!�dΠ��s��c{� ͎ 10ĥ�3.�Q)��jQ���s����xy�4}�.�M7Z+bL�w�eE �婷ܸ�|N��G�z��>::��c�v�KwQdެ�Q����Yj��\ߌm,Txr;�4��������B�2�n�E�\m� ���|HU���C@ѳ����P\��v��P���O�,��7�}Bm��-QLwT�hf(�Jv��IP�8����������X�֗��!���~�1�Ulϯ���*��78a���Ë|�Lb� �vjŢ�|�uEچ{0.���Ԅ�i�8��S6?��ՉM�gaW�QC�U�1G�X�%v�4� NT�umܥ�U�3W6�k��O=ҢG�w�I�*$؎j��GTC��Y^ b�FS5}@�g7� E�\�;�f�3k�h!Z�I�I-(30�>&�ŷ���هl�N�-?��w��(,�i�
��3A�F>����O� �=�@�*�E#�Q�{+ӣo�~sؓCܢ�t������𵙞��-�-p�\��tQv�㖮����$ꝛ&]	��V,TU���c]�Q�G�;�ٕ@��(yv��XJ�?��tq� R<F#qL��}�##�[X!�9'�,O�n���	-�f�l�I���e[W� ���Ae=/}�O�-
�u^�Z4�K7p������S�༑i~	OG~�CζHD�C��$�u*���l}F&]���w��1��d������l]�l��7�Q��~<��S�z��k��T�ңp���xځ�z�Y�����\�*V&t�
E(#�����n�G���㹿�g�`���3���b�����s�
l�}���e� _=CU�aw��&߼l�G�)��M!u�P�H�mea�SJ��G�8�Xb��c{��'����a;{K罡̢���q�-	�d2���1�z��V%�sC�ע�S;%X^��X�	�&�, �Gjk(�.�1A5ÿ��.9�R��侧[1s���	|�\G �w�QMQ�$�f�j�B���&Hǈl���#s�]P���,2�)����������˪�6��El������g�W^z<z��7�`��1-�V�_���M%O�](Y.��
F`Hǳb
e�z�˜�����ρgkw��ۦƸu�6I	���`�un�����z*�I5%�2�J2�'�B�c��h�G��3�Z�{PD~@�)��ć/6<�$�q�6>���g���(�+%Jm��me�Ɗ�@�c�'�ص��� ̱����gP�k~o�1t��0}��m5w����J����JPֿ܄����4�iBN'Q=�@�b���w'k�}:]���đ3ǰ��0��w��l����v� �K��x{�r��^+ʹ,̀�N�ɒ�<�b�yD�I�L�9.Z��@�-�ձn9�v��pY���h*X1�L��_ϰOI����0!6P���'����X߆1g��V/��J�.4>���T3@�wM\#&�}��U)��7ŝ�Q�	���td�p��p�q}�ȁ�ر��[+����
�X�g�?oc�:���M��ēص.����p���݉��X�k~���uɦ9��� ER}�.�
����F��G��/��U���V�@�t�L�p>�h��x�o_͘e���t�\B<P^��ײ��~*<0/!�r�j�[��t��jJh�e&���6@��ԏ2}����A�ٶQ��� ����͝gc!��;���?�p�����-jfU[���f��M(��X$l�X�f����Q�!t��s.pv?�* ��}`��ɋ����3>d{�m�<�H��{Py/A���l�g@y	Z�H��U0����q �<ǎ>���f� �b��4��Ac�����V�؆Ow�Qϳ�2��雒�ͷvX\$��q)lMHLm+kkul!�NQ1:V�7�l7@6G�a$�B�(AC���M?ZJfe����a��G{̇R|������E@DTХ�Owp01����T��l��ҋ1��RP!���{�?G�}Y�#�_<V5tw7{V'�=G�U����nw�:W	�zsb)�K�����6�@��]���@�<�Y��"	� ��|C�._<�L���o�����4!<,��=�Ο��ֺ��QYg��!_�ɟ����K����p�D����$�M�/�B�R���LehA,Bڸ��LMf>��f~��x���@D{�TE�ko_�)��9(CSEg�^l�,�5�6���c�	Ϧ��f�|S�wx�b����=o���ƹo
-+���H��X{�~^o��"�Aq�v�
O�s�"���n�h�!c�'0�Bz����w(�����R��
��4H#�a�S��^�����( ��3�o'��P�<I5���ض�Xb��A��W����Ϻx$'\ƌ^���.d��H_�;z�7�z��5vE�r�-xֳw4���I_Ok������ԍp��z�G�VR(������0��E8�6�|"F]�*{��0%C�|H��'���ju��Z���}l����Y�;
*���L�I�l��d��G�ӯ7H�J@P��|1r�Yh�E/ß����(���Ir��[�O=~�s�H�e�TP��?�^�>Q��`w���D3o	�WЉm���d������.���c`�\a��h��	�	T�jGl|�ŕ��#�(-��
ZG��{��)��,� C����[���{�'s�?���U����$I��^������� ��C���^�������ծ��<�=����bi�M.Z�Yj�´%�K:�2��Bd����y7�$�2���7��[����{�۸�F�ʬ!�����p�ef�Ё0r��&�t�օ���0��}?i�4�'�@6�)�f{�Ɏ�Poay!�.OR�,z�n�v��g��,�$��ö� T-�;f*��zp�,"
}
&�<F�|�Ԥ�GTo�R@��2i&N�����S�LD��k���F��?�`q��)�4Vu���Y�2lJ>���3��/)(��%��F�'�ӹ&�[��aA�W��L���"�ve!���#��U�	mA2�#W��O 0qa��d�<��=�=�d�rp��j�(�.���)f��ߚ������r��uq,�b�Z�7Ka<k�f�/��#�S'~�a�������P�pv���;�$�Jq�M���!�j! B\I���%x�kg��j� ­?Q.�u<e��z���@�Ch
�:-���j>t�9z��j.;�:�cbwt�.a+0��vg�5���r� fL2�s±�W�ۀֆݘ;C��:pr���1^��t�G'@ލ�g�Z`����z��EN�7���HV�WfO�E��I��p]�VVߕ7�T���!ց��o�zf�{n��������~��5���tO�Ф��C%�ڑ�Zg�h�O��f�U�A����a�ތ�Y	m�=�c��袒�6� ������t��k�6��@"Z�u�=s#8��a�	���%�yDd�b���Df��&�%_C���6�RK�W�lJȱ��vo�k_�gt9�m0bm���M>�F��/vuM���t��A^��yU`��}=]@��⵬�{�.��c�G�ŗ�3�'6�A�}t�#��$NH��R�rp�k�mdV��i�����)�Y����@\����Y�0�3/���[��݁������.���>�0_�(Q���mC%*���aq���pC�Kv ��2H�!�^��X���`E"Z�a���[ru.3�?Y+�/鬇A0�H2�~�L85�z���0�����*��&W�_)�eY�&�U��G��wq����+3x��c����O�21��"F�19�z�*,�D��(�����S��k="��Y�FD�w�9 r�zJ�Wc�f���9���y^��Ca�x�r��L:�#Q|[PI��ale"�n�8sX�X���P�����a����"|R�7i5�0��2�.�x9\;e-ʋ�>y������Fr�Z)ެ��ʾ̄����5�LKy��O+�<�5H�L��S�ʣ�d��u>��ς���N�����W���)��`jl[G/���e�������
�e?lμ�OM��NFţ�]��"
%1NN'�k"�LP%��M;ƖBb����xx�#hiO�'h���iC��d��>p�2+bVT�V�D�m��5J��F�l�2	/K�([�F�G�	�k��~��5�w,\�\�̍��%w�&)8��h��n y�F�MD��M��ߪ%�7������v����JT
J�����~A�aå/��2�8��l�u��W/FH}bn
L��"�P�K�"0�Y���^�/��(�F�:��u�/gp�h^���:�e$�:��ޓ$��K�֭�gY����/'�O�"�7[�u���� uj��)�Q�m�v� 5��/\uB.��+�澫����T��p�Y0��-e9X�����Nhh�0*bP�q~��W#s�So��uG�����?���"�ۦb��l��c�W5�v f���� ��El��$�>*<!��mYw���ƀA8(��3X�q/tp��]~���.	e�V+4�xX�yMa�7?WC�u`� t,s(Iqng��H��cd�ɇ��
䃷��7�t�[�ᦒp#���/S.a։m+�5V�`K�u���αR�[�h	3&x�ްuS+���'s[�#W��|�3������QA���a�@�����ڴ~Ԭ�N3��B1n�IB(tK��ڻׅ�b��2��o��O����V�F�D��DH�ݵ��0Ӷ��/b�����I���(�6DզY�E�{�~����R���#La�&��Á��q4l����<��P�~� q�����q�]R�ށ���sޮ ZK�p'0�Oz֤Om��1V��cT哷a��g��-͸Y�(�V���u|⎎�:fF.0tMC��{�����V��Q�"�~tU�4/��K��sk�C���;A)�8�C�������h%�4�S�s���A�x'�~(ӆe'�
x�-�T� ���=�3�+��?�pWY8�Mk^u� �Aj��"V�ɹ���E�#�ŕ�����N@��Ӟ��?W�bٽ�v�B�ywy�G����-̮/&J����Z ��Q=r(�Bp[�jÕ��:���;f�x�P �$P��&�XN0>�㲄���!v�x��%���'xy9�phY<��q8Ğ������wXb�q]���3�L^�`.��6����Wp���Mwֺ�PN94�N	�
��P����2	�K���@c��[�V��/��]�)(ǥ���"�"QT�!;���jҗt�įsn�Q����s��[�s�"�lfS�d���7�7 �dZ�Н�"����d����I�Y�>���Q������,Y6\���!VX-��w��$�����7� hc�,Y9t�����r�9�M˜�:.�(H�4T����eD��?	�T��Kq+n#�����C-J�B�;%ϦvM���,���L��W�� �d����$�EƉ�s��p�Z�"��5�TG��#��jSl�)�����;)O\4��z�6���} ��i�ů�9�O��\�.� +Y�!���t(�ߚ̇^E�������������O�BD!H��U>���rJˇ�1��c��������p��߈)e���w62h7�X~,2���D*��D $ 5��[�Hq�|�0O�!�H�̃v�&�-g��^�&�U�Ė�>�����j�u��[�Dֹ���"9����-U(_m�qρw̭��D�e(Æ'I�u�"�
T��9I��8�e���uRߕ'+���*�}�ͨ1cd�c�:�w��{�g� l��р���\���OU��q�%��"�3�t?��A�q��q#צy��p�
��|}�:��Ɏ0CT;ރ�9�BS���h���x$��Ͼh�Җs{�\9�T���w��Yk�i�9���������������V����`��!F]$�j�p�f��sL� _p�gB��Ϫ�&��z����@�U��'��|�铭��� �	O�JR����s9��S��Ń�/��)�P��jҝ.�Bp�Zb�^v熠�)г�{�U��ZO�C�ׂ4�����Ը�- �/�����$(����5|<���Z�.�	<�8^o��vzb�����5ut)"�P���o��gyL`�����TsP|��Dʬ��9H��+�C���	q��j����1!?"#����O/�l�;���KpW\�WKw�\�o��y,z!A��]�O���O��BH M�LJ>���K̗��Y!��x�lQ��C����~���>7*i����Ruo�jd{P��G�a�u����(�^�����|Dգr��M�W,� yb�n��e�r��`�\{��,52 -j�a��`X��?��p�dUa6<���D/F|�e#�~$)䗙/��/�Ehvc#ƿ�[
4 �Z��3�a���U�0�MRz<b�6�;�J"t$F6�K�ݛ�tne�p�~���ؙӞ1ۛ݋��K�$0c��?͓����"�,]\`/�1�tz��Qݧ�`!�i�uP�?O�P듛*T�;u��?݈c�Vri�a��b�e�� ���N�N����Z
dfj����l���mj�c^C����;c\x��e_�&Z����&N^��C�jfi��"��^uE��\Z+}8�9���!-����c..�B�P@�hY�N/�̹(�=�!o`�MP1^O9��/�#5k�����>�3u=<| u�`���V��)t:rƛ%"��f�~��� �e�f�]x@�e6&�KN��X���Q}��Z�j����'o���f�قpVZC�rs��.��|_5�9.�����Ώ�����4r�h�!z0�y�%/�
ol�A�n-����(p%��x�mq_{♤�@:W� PB}ͯ��������ѻp|���Ǒ�a��$�M�����µZ~����v~�_|,�?bBZ�4�6o[J�� ě�����B�r@?%��A/*�!1��D-*�!h���_��լ��+����֧����9����{Wy�-�:}a����W���
=�Jj}|*�:�P����v��Sȭ�h�+D���uE��ǚ�Qcg�B�M�7*[ak�ҏ�*<!B� Cfr�4��NeE3�	�����cy�=a�f�DB�Gnn�ϴd='~#�@�G��7B�ޥ��0<$W��CmUg��0��K�F�}Yg��I|�w+�+��k�{Q�l��r��u�5�`	?5;��ŧ��6��l[�'�Ż�k+�^�>1�����S9�:k+g@xYm�\!ג�o��<+j���E��vLB����Q���
x�'���٩�sB0�@q�%���4�H�/�2�68f��U	��ua�آ	eNX�o@�>/T�趺⬡o�R#��z�i��t����]���Og:��	Aƿ�s�"~<���L߂� 4��{RA���Ԝ�4�蜪Z��n�_�� ���fy��Qض65	ő�Β�����E�x�cc�pT��tt-xW��m��	��	����ZT�>�{�"B��P�Eܴݵ3`��� �k����9/�1�� �c�ߔ5,�斛J4tyI�Pj��t"!ެ	�cG�T�Rk����6��\ҺۤXd$�G&g&�X����R�	U S�`a�ל�Pwe�P�ڗ�rȇ�tb���oV�6�TE��:V��������&P%�Ђf���2à�h�����A��~�zAgB���!��F��z�s0x�	ҟЩ��D�N�����觕�+��QF�Z�JS�����^iP�&�fI�|���|wj@���	�[�3-��ߥc6�7H��L	����P��L�M�ؐ��aΟ�/ЩjF��`��	JW��������X���0����n�-u�n�$���6dQܮ��B0�v�M���� G�lF���u�ĠAzM�Z��ԨW��M�ɝP�̃�J�(h��\�,�p����c;�۟R�`pw|��L��y��Q�.s��D���P�^����͘Kl�p�6����Y��eآ?pA0� �U��I���_Zk.���'����>��|]f(�{��d�di�_��p��wQ]�f2C��1�_J�F��_�o;�F29C���2�1�}-+�w����1�k�=D�0�:,�_Ǽy�AOԿ�
�x���m�A6w@��=�	g��L��?Lo�{�{���s|ڵ��=6�j2�v����F�7�z�=�jzn�Zn���lx_�,���6���fK�φ/�['X�ܥ15�J��jQ�9tBf���GC�ɵy^ �P�����g�`�B�i�/�v�?�@5F� ��c��s��0��d?�'_�C�!�|)#3r?��HH��u��N���⻖��,�L�Wy(];� ��.�)���	鳺�!/X[e�tc����O�R�h�����������Z��+���Y����5x�x�����2� K-*�nݘ 'Ksf�v�js1<{�>OH��ɸ�]��ist��a�� ���%;�U	;5�e����3�������ʄeJ87��[�<�a%\4	�c���'h�#���#�腢F�9e�D�.��>���'l�!�;�)!�<*hO�����
�����N��|2�@�˷������εg~ז �]i���N�Q�-���z�@�5�]>�\gB��O�U9�ê�i�� :M#!�u!B�b5�����Ok`��3?��K(f9�Q�`��h�F��6���x��԰�/��*�d^��#^�{r� A�n�8��x{��~�A0�|��
LV�����J<�^U<���L8��틂��Z!���� �x��� �<1�c<ή���$~~�WCl��%�0I`����C����(���$Cv�+����!��U�
�5��D�\3����e3 `jݪ{�>�2k�V\��29�obyri(l�{5O���.t������![�)z	ͪ&�v���$�� 
kI�8p��Hռ1E�f	Ej���
�E�'���Gj��Z�/�{[73��#���wf���PY�4V{t�1PJpѪ۸�
���a�%$�s����%[�F¾a�'!A�p̓�����ʐ��aැs�k��X�)Eċ�[�<�G������$\v��O)�a��|��h����E]~Q��š��q��\��(Y�k�}���E�����������T ��M*����&�����?����5ri
�1���{�-����ւ�����3�Σ��Yȋ���;��6ja��}SM�N�se8���-��N�_�BG\F+��6�2��'���U�hL��"�bK�a�#�	�%�~F��M�F2$��zV􍩆p���u��2D06]FQ=kQ��[+L�0��#�<���+�|�E�Фt���K��|A��a�	�丣��D�
�]���O�����G?�r��f��r_�0�>�x+Ka��d�9Z�4޻o?_#�-���au�:��O;��Ѫ�~h��$>�~P� ��,�9�&���}�[Xt�(P�U���M8�ļ6!5�(��$ed�h����ɷ�0.���3�+d��A��I}C�8�\z}iW����9kZ���wpL��&���u�3�Z�`��=9��2(�f�4tz���Bt�u�̃�
[�{�k,ڥ7J�u6�>�ySy�����x@5�*
S�c>B)�E�i�Y�趷>� |�e���) h簁��4a���n�&�D�Д���f�>�M�m�x�IA�mz�A��W�7��Ƙ�ZA�WY&�B��3��V��Co(.�^�n'�	<5q��K�:<i��C�R��na{�\�K�g(	���(#�U*2�Pu��D^���^��6�U��7V��ѓ1�S0lm��\�@8���~��) ���"vܭS�C6�[H��!a�M�	��s��%~�k���Qj�
�����W���}� ��䭈ciȜ�2-ę�,(r���.���Ԏ�F�n�7ٙ��RREB_�,kk�a(O��C֠��7sY�6�y1�F��oO��r�?kK��^���3�	��LMa�Ő���b�$oߘ��,�Q7�=G��n������#��������0�`^߁�{���p�=~�P4��w�L����u�OeR�Kৱफ����!�wHM�y1x�ͭ&q��wVݏ�Y��!�Zn{o/���`c7][��]��ջ�<˰?�id z��"�Ssfr2L��k�y����,T��b7q�ρ����oOb|r1̳�w'y�nKy��*o}<LM:��x2Үjf�5����c*�q ��cN���JDړ^���F3�I�Y�Xξ�%n����wS��s���+2Z%�6CA{�����g>���o��y��g��nHK�y�*�Ux�8B�O|�X�"�q6��O����i9U��9q���؃����9�u&�w�Ӝ����lIU%�X�g$���*#��Z�F�;	�I���gW���i����M]r��-E����q�i��C��j9 ���>)Ș}+7�:&-W�|��n)@&�v����]_;~u& ��	f��6�����U�@E���_��X�H*���c�>'�v7���o�A���WX��OR��gH�%�XM`��u��n�k�mU��S^.A�a]�؁V�]�VQ}f��V*�y_�m�0����j\o��U����՟��y���c�m>�D�����E���V-�t��S�ع�3MZQl���U��L�m�����@y�v:�Q7-��z9�`��$��In�`���mB0y�P/E�:���R7��&�������m������nw+m�6�P�`��w?�|�'$D�8�ʜY�:X#.篾�R��Z�ę�~mg촃	o �G:�	T�G�	�}�R��<����D/V����>�ǝ�V&��7��
���8��P^�gP={{�?I
ؗ�7l���~� ���>�.T#�9\���;"Z�����*l��$�wd>���j�{��I���K��h0��=�F)���R琖m�#��ŭ7FI9������ǖ�����_��es�G�z[�G:�wRtx�(|,65m��ew.�`Wn[	�Q�� ߑ�y<F]-��8]W��]��G� +�3�U�y=q�`���#�Ϥ4K!]�8P6�jA�vO�,�D����A�,��mK��f���I��T�%s��M+n�#���B�W& ��`��k�$y���A�Tg��9���E���Y�i�u4��+��[���J��i�jLs����g\��iJ�i�~�c���ģ�R�#F����� �	a��G��զ��V�uo��ؙ[@� 6�{�4m���?�W*}|f��7Y���u��&��Z���!��j��#�K鬠F��*��)F��D�s�S��_^9o\"q��c&,GP�_>��Ѧ-8���&[� ��
�V<I_�{
�+���XK���]8��4�g���.-i% �q�gNH�G�a�*ceіXs�d63���[�c�MC���>�g=�T��S"�Q���0,��袤J~���tw.ѷ�Rld��`�9ԉ*l�n���[Dȥ����d"�r[��(Ͻ�~��p�����BEA�k���}ߕ�:t����=?� ���Yd�>ў/R����{e����.W���H?�3�pV�N��o��wp�4U}���A�.=�M�x�Wh�)����l�1U��� �F�Z��
�t�L(�,�8+t�P]�l����|������H}���@�Y|�HOʓ���gP��qZ%n�[;'��&�?MA�w)_�����M�P�[ɦ��a�_s�^�	�g�~���Q�.r&q��ʗz�yo�Y��㑄X$74���� �'`�O�b������ŭS�x�暤��+4��p���n�|$T�T�;bs��	�SՆ�g�[������a�)��e+Q��e)�k�Z�1ȋY��1�v��t�KyX��!e�{���V��d����MSi�]FV��t/)����i��e"���m��y�n�6>��W-\�v�Gz3�p�uGx�vI2�g�$����-�z	T�6��7��@�����S>�[C�i��N7��8e��O
�l���d@5���W�C��t�Y���j�F1v���Һ_wU����,���ein��A��6�##b@�k���f��5���a�2�V��� PH�[(��'���ð�*_��T��Z�L�l���<{�� �:�D��p���Ef9~xL���'^�����+�ux�Q>m��^R��.�� ��P�u����>p��2��r:�
°Ύ�+nw�?3$�$�c�FP��+��#\�����Ub��Y��C�$C.���=W��WTZ�Ш%L����"E�ܹIƉ��U�e�q�k���=l��&G2��2��bQ9NL���qZHf�����-����}�p�NN"��/�.�y=��5��V(�����廷M�$�R70C��������N�d�D�:T�?���/9�C�tg������E/�=_b�.a�U����ޝ�v���M�n@V�WVȗJ!�uſ��/�ALe�i_�Y(��Wjwx¼,��j�$��+�����!����6A@k�B(����|�&����Ђ��C�^-"WwM���^0�T`�^p�^�}|[b����b���G:kН6�W����X.�c�P��؉��ᇸ��Ae!̬m6'�Zt����	�	Y�;��ʊś�Px���N��� M5ӎ3��VF�'dl��;b�{Y���Ub>�(*��*������r 6�/pl�Y"���O0gH������i��/`���Z��I�ü��c<��_E�|`�������T��-�l@6��YS���J��Ư�2��	�IC=V��}ahut:�_��d[���S_g3��{�~�d�h��SH�
*mP���qx�I+�q첾���s�(N5/YbO"A���1��~>�e<�t�mC:�{�}�@��6���2h�Ւ�nL~uA�P���s�v���2���LU0|��%������ۀ��q輱�E07� �lv��am�W
��z������+���.ɇ��]h�ȁ�i��p�>�%���_x�����z��z����M�����5@�(�������U֣<L�+	��D��]3/�W="�\���Y""�nT˵b�g�
o =-��Zb�֦4��,�j��\#�;-=��c��Ő������w;�^
��=7Vy�J��_�x`5���sZ����?A���_��(��Ǖ�{��Q��Ux�
<8"�75�G0�ʦ�N�ܚ�-v�G�ƕ6���=�}��8���bܶ�w��r:�����H�M��%I���L��d��f�(�"/1K�{5�}.��ϭk�Td#I5C�ح�I[����Ͷ����&*�7m�$9�7������!��)���Q(�w��6tqׯ�p)zq@w+�%��^3Q¤5F���G̨�[����O'du�@K�n:�RdnX�~7v��Q4D�3�mq�T�d[�K�6�x^�� wqo07��/�*���|q��j�k���Fi��C�x�מ#o4D�a�"-5���BMÈ���}��u_��糿UD*{,���Щ�F.d?r�q.|�%��/����ꄥ�;��"C��A؉�v����+-k��䨣��X���7$���f�UI��Jׇ���׍�U>���l%�"2�3��L���.��kd�n[F5��w*7��$p�}p$��ce��ǿ�a��R���r&t�6�]zww�f�+(��V��A��L�̌x�������4V��(��)_�t丰p��g"�]�o�^��5�8�o/��.�"�~�T��Ni��0r�9��5Se����t�L��`D��ǚ�.�:� ɷdr���\�N~�d��
eo��O�u�Q��hy(�X���TG=�}�L�}V�!~)*wŵ]�V��;�����A�/<5�"Q��s�����pç�rw[�O&��i�b���S�V���3^À���Lv�g[�7{XSYܪe��<MN�U;^�ʢ�<O���lܤ�CJNs�[��ܦ�  ���pkNR)��=dI��%|���@�W<���W~��ص����
P$�S��%����ڪI%{8r i�K3�΂�iS�U���w!���2�Rl��K����&p=~V�0�۴	�o ��|��(H�s^#O���2��2ah���q���wDLׇ�����S��r�.�N.Ѳk�lH ~��>�Gs�b]���yפj��_"�[<�mɗ�Wf���®!��Q�n�n�f2#A�����h���\hy�Ͱ�~�����!�*齛#� ���]y�~��D>��0�ۧƗ8^^����!gmC�
�X�>�Cj�h�6t��o�Z2���R=�!Y	C�K����[��z��0�2��7�OG�Fy�?����9�f||�wuA����϶�~CiU�C�у����̿wq�NuDQ@��f��lN4��[}t�̓?h�?�b%���!>���P���Gy#1F<r<���k��0is�����1�91�����I���/Ӡ����lŀsL���Gf�OD�le6@6>�o����72Y�7�Xe���g��4f-��z8r���̱��9֔۾���%�-�@�:<b�e�Cp�����8	߮a�l$|Z��W(�C{č��e��g�Đt��2��%`0�[�Z0K����t����v�1������^	/d3��O{��z���ta��D�� K"���^�0{�w��q��Z;#X����ڀ��Zk=g�8��ܝk^P��C:q?/�Zh��t �=���;Hhg@�WX�v�&sm?l�w<�ӡ��2$�0Y���EI^Ù�c}Ҙ�Ł��^/q��*�m
�M�")�����]� C��\�J�����&U[�s�M!��v�M��Y�n4�*��A�����b��"�z�DR#O�`֑<��&��iz�=i��勢�1��ɷ�&�\:��J�ڶ��}l�ЛF抉��3t%G6�#�:AOґ���q�mV�<C��1�Xе/#���iro��2�&49a?��0u��S�%(L#��C�	oaȉ�A�x�﹙��&�jLǉ�Vs��Kip%��O���Q�����(r]��B��u�^��?&���9!����=�,��*�� �c.�����S��27��D���Ϟm�6H�bf��z�	�����2	���0�E��ySg [�c"{d�2�9���!A����)�kaܦ�(5���}׿Sp����i�.o��(N�ɒ�Vٛ���۝+0L ����A����
�05���S�4��T�[�U=�����R9�4����w�
ԏ�������+��D��l��JP�����Ř�d:w�`R���-��e���L�V�o��ie� �w�����3�Յy�c�m5�Q��^�j�̛Io�������}I�����%kr�-�>v΃2	�H��k���A`kY��&��h�����!��S�9T&Hdvh�y��P[�+�l,�P�?�g���$`��f%$!/��F\Y�e�~��̸=�,rGd��Sҗ-_9�\P�W]�7�N�g�A�*���UVsR���9�;gJ6Pm;�S��Y�=�=7m�:4���cg���	�1E��3Vd|�٪�lW��sؤR�\$>�sy&�﷉xh��vSj�!�W��B����)"Jx������E�s�	&���'���e	-�w>��m����V�@����ݶ!W���~�N)�M�4x;!����w�6{�T��S��sWOH}�q�.�˷;:�i�~������(���#K=�cP/k��z�?y?��/oY�_wv)4�R��aY�!M
k ���s*Y�X=q1��A4%|U�h4��3J��������MQdc�b`nhPM����.J�[� <�֜�CD��\����Zڧ�ѬX� �$S�;�UBY�����#2Y�|cj.��o�T�u�\C-7i����)�;!�t�92�hϱ��Q. f�����Q�2\�G)oJ��Ek�g^2�*�fO�|y&O������߰��p��u�X�_\��Pu�0����x��BfYe��V�t<�%� /(5��)T������"��%Z�:�zT�Z�Jg��nh��{�96��%g [ ;���lF7荆�m)o�=X�_��r�3;��Ej|�z��Ƕ�p��E7M�I�=�|�O�0Z�A�cȂ4���6,����fĴ���4��.O����|��|�x0"=��^)�����%�r��,�p �=e%V�*�0�1�4+���ϼ�פ<�U���������A�c�:6UI+����i|����cm�4��?�_Ep�Z�ܪHuk:�Y����Y1E-9yT~��m; uG�ڍoe� b ����o�YG)�@����I�Ge?3��`����P�g@�/��z���@�#�hU��6�h�[�� 5B�0��vn�ʖ�4��e��J�vn|�%\�S����)&��>��~]_���}��4B���\��Xm�fuN����OL�5 �ubX���i fS\�����Ѿ��d� p�ߜ��K���E@�,����|�J�����\���E�#鍯�mQ푌=�;{�6C�T��*�!�C��?��rs��0~���ΪA��R��L
*��@��1y��l�x�D��)Sy)U ;p�%��Uj�r
�m�2� ^�5���K~��A;�H眎�]��|j��)@�ꈶ�W@}*xh$���sUCR$�����$�n/Q%��m�:Sp��JUt��<$��+���ظ=��~d����=DG��%�"��;��tQ=�	��)0����Z�l+Bc��l�>�[�"-Pd�NV�Ul�X�1���Xm0G��L��1^�q9��4[|�9��NC�<�l�0�J�ߌ��xƵf�3F:��Y4~a;?�6p!Y̘�h�y@��(��/_�`="H���Y�:��eI��pve����[Y���>���O<|�h:�W)����e{��Ph�y��N[�`:�Ebp�nKKt�e�J��v2L?��g����\�-#+L��	S\�&��sz�1h"B�I�w�n�	+,��FQ��	�^�sߦ+Z��T���8Έ�A�쓄��ܪʁ_G���MjH��5r�UB)�8��Ug<�VQ��A	L�>�k�l��F|i[�o�7qDg��������W���y����Vj�vi��u����_���(uu7ͷmj�4Q	������,�$�V��;ު4��s�T� ^GY�mR��O�����tL�Ao�~���Y�&���Ʃ��Hfzi,����7��i��>w:@M�%JvH�DP;�/AZC4e�M���3����X�RY��Z�"�t�%�i݃_��B�ԻOd|2��ڐ~��)��#��C���?����_�{*`0������f�n6r/�-?fb��&�:��{F$�V\�vܕ��2��������Oė�<'x:�3ձ�sr����~)��ʶ��^bB�,r��oFAu.J<;	�	����T(\�h�����{��3M<u�@�W�Q��J��<[Q�L���8+����-��w�9cM L��!��|��VB�.�����F�����bt���M��Gן6�r"�abpk��Z\@i��^"�7�����3N'�<3��o����q�K;9=_��t�{�v�Vs����� ��\�6��{��Ϡm���l�.�
��p����#{��%�a�<)����=��<9�K,��%%D��y���z}��}�����5>�N�D�gte�I������J�OXf���Ł����|����񷪽�ꗿ����:���z���� ;x	��`z�R'|���i�}�����lԜ.|�NX����dr4�h��Q��f�&�Ħ�dݵ!�`��n�u��e��;L0���x���>�/X��<��}O�Ns��'��YF���Ҡ���/������Ŧ��۾��7�Z!iy�L� Mi�L'N%,�V����+��ލ���3M�UKQ��9�hgG�o�Է��4O�aר]����G�a5Mr4b�>�rdba�gK�=��.�1ÏI�؏u�ئv�>.!&�]�����~�#�1]Ǒ���� �I����5{�֮����1�07}^P�v��W���_8�{�s����0ȏ ,�uJ�7R�N;U
��Vj�
��9����F�F$��g��B�1o͈��3 �QXU�[����W�I�%àpʥ����s�4���3�*+�vcC�e����������P�R2u,nF��s%�7Z�Ѝ��� �V]�\�|�.Ɖ�D�m��q�}?�H˖O#œ4�b�!�����L�a�±UKUF�7��g�"�f��r������@Q铲�!�3�����2.
���k�.�q�AG��]���'����ӣ>-�Bw338&8;W�{�=0��ܕ��c�#{�z ��n�S�����8��*.� R���A�σ?vuDu]/�I�K�4z�Kc�+#d~�m���g�ܲz�R�d�������'�z�o!�ƙkB���R�!�/�U=�5&d_�̵#�����n�D-������-K�!�
E�	����_ԧZw'����&��v�!ڰ��ϣ�;;3��ÆHt�7;���0A��N�١���Ć#���s�:�Y�=��0�^U�8{�}i�b�Q� y�|�n�2����ƃ2�8�����O��P%��P�Zug�S9����5s������`�,�۱	�	;�u����]m�����*{�Rd�˪�"~�6�2�F��ke���tD�ې@F�����{��]�'	�쎐X0��H� �j��'��m��M+�'߫aN�4j.�
2�Y4��\��z��'ÆՖ�>nUD9�U`x_�
н=<�m./��03���ظ%O0����16CNl+���If;iu�4���I
�Y$K~�t�a�(�������]���@Ёq6�L^s<���q��L���%Bq�:����J/���������sB�V�i��1����o�H��|�?md?�l�vW�����tz`�23�Ap�.9�����RR�o���������vAFO��д*���Eˣ1�l�c���K���h-�{�|�fD�Y�d��n��VC6�#{�]�5�/3��S3�3� ��Pϐq��lˍ�HԜ2�E����'����u=Gs����)4o�J�ɹJgW$��G$��7�1E��l$SQ�\ �ͪ��+b*�M5�x/_�M�Ӧ��N���/������	���IJ~M�c��Ntff�|d�Q��J69�f�J�قjb±h4�/��޸�����X�,����HPh�-��i���t A|NMT�Fڷ�(�N�G��о��R��2?\ԥ`b�n�(	��M�E9q!u2�����"�u6*��څ�U��Q��N���7Gj,���V�8���3߷�y<�,���_Yoa��!w����2���e���U}�	��?bU�W�O�N�JBW~x/���\�/^���lP�s\�i�O]a��W;e������^����P~�䛋_�(� E y�psģ#&z�LV+	V���%��'XP�<Ю����F%P%ԕk�Z�q�@+xa����t>����-��i�Z2���RP9�;e�2�5*AX'�,�ҍ�Z3����F�����Ag}γ���77-��|ODYR��e��L|��Ԑ���-� ̅m��[�Jiױ�5<���{��qٰ��qr�|���#�Ϭ�
!��	a��(n��K�\�$�4��v��C��4��*|ک�>d�bg��O��=OZ(ˋ8�����70�7#Zo�/��0�_���-	b��a���tS�4d����K�i1����!ҫ]Md�{��gc%z"@R�N3p������oT�M�}Ws��_w���qm'�7S�8{FtR?�Ī�j�[�?�-�4ȧe��c�����:=��Ӡ�:̊#�Ƭ��D�H��m:(���qvC_�h����/ [_Rہ7�5���/��ɴ�i@�_U��ئ�L����HZU�b��~�j����+��rS��,��]�%�+��Çg?uBj"24�g;�؅3֐�L��x�W[�#�8�X&��Ҭ���lX(��u �\��V�Q�f�Vn,��ΨT��׋+ �8���Mtˌ�sq���&���.GǠ_+`�%(#w+(x���*Ĭ�О��x%̤.� �-v|�t�˭s?yP��3�WC�v�g�4��@>�>�Ni @5s���F۟���af~�[��@�y������r�i.��C�4!rۙý!�c.Q��u� �Ֆ�RU)��:��9� �`�7o��Q��@s��F|���Ç}8u��s��-�[i�����w�w���! �����uR�����m��F-�A�SЬ)����!�e�T��7'ؐ�K2�(iHv�r0���yC�u��#�@��K}�b�� c�⮴%���ߛS
�h�X\U���@#�J��ɽ=s��Al;���=r�$��D���A�%W{��,�o7�Cՠӟ�u��]�F8�zU&�Ei����@��'�o����E���%ΈRp��,Y�݂L��d��s�#�P�W�Ubo��b�IQ$Ef���4lT��˻R��J[
N��Ĳ��v���qܐ��K�-"� 6�-� ��BR�tjj�"Ђz���d '��a�����p�5��%i8�=�fχP�T��mY�ARb�����nsؗ7eh����_t��/�M)zk���[ g�;1*7�
���C��e>�9�݂����yi�lsp�v͆#��O�q��$���b�!��t�g}qulBr�sPlu��Tr�ØZ@ 0t_�����J�ҩ��0���Y�$@�@ �"}���lW�<�����&ıWF�f��%��hS0�c /�Y�\�2f���X���ۣa��}�Wm
����oNx<�[n/܋%��*��ۅ�F�1�#lh6F@�c�'7(g��[ߩ�y#��-��P�����}:�������C!1�e��@\����i�}�]zs��[���8˯�� �I"#Y�W~��W�FA�%��D�P��J�pr��$�/�aڳQ�C4Oon�򷶯~B�֩,�H�%��ì�뺄(�?��6��e�| ,��@��Ph�f����#Y�*�A�����r=s��OIL�9����wh�*/P��+�߱���j����F��0�P3+�������.j��Cta<s���<��5�س� �\���'K������8�s��{g������ ���X��>z�cKH��U!�4����	�ؚŰ�Tࣕ$m C��gj���C��)�bi � �pF���v�s�N;�v��D��f'f�D����Q=���r���.`���ת���L1���!���ZK>��~1�����7g��H��%E��!'��X��k+_������<97k%i���MÈwD��@E�O�J@�a��<J�	6I�JǼǵ�$3%��� ��)�xE����`#�a
#�-a�^l~�l��a:d�~��������|��t��	[_��ڐ�C����<זM~�D�;0���28 6[z�N@��l:"ڞ�E���X�Vx�&���CP�L>p� ����n��oX�_�0����ck�HZj)N A,���]�O�0�"����*T��I��^����f��%��k������Y�����p�*��mظe��ڔ#���4�KA �'�����g���'1-�9!ݟ�@u�U�e���������ASә�#�H�H ��`��f�Q��<��>���$��k�&�≬ADbg'�X�E1���L!�7	7'tћ�6����c8oˮEHd��^)[���uõ���\�S��mˈ�*��L[���e��`ـ�j0�K&~"�4���:>kZ�.aԹ���-�S�TF�{oF+��>�����mnŭM��a��-��@�]�B��2ؐ�� Bֽ^��n����<:/sU4Q��hM���|ʤ��Do�j��4����&����lP ��Ǖ������G@��P��$J�+YT)�B*��Jk���i�8=Д���/@AM��2�3�υ.$�UC?�p8�Y�)�>�Z}��ı@�>��%C��u��Η(޽���T�����jJ0�8����k��Ԇ���b����\��<:�6�R�tP�E��]�ML,*F��:7{vd:!��C��v�����*f����j_��<=�AM��0�!g!&_�V��kBF�E��M7��U���M>Ԗn��Q�T`Mfj�z�s�4�:>-�.^��f�+I�PiD�~��j���;���C����n4�o/�_�*���M,C�,؀M6.���z�|��+G�?�G\)to����Ղ����~�EY Q�o���wC�m�?^u�m�nk-�^�VfC5���s�I�@��H]��4��T��VO���($� ��ݙ�E���i�Y��!8L�2y�Rqsj"^d��M�~�!%;�^hU#݉�4W�u�&?���~,�k��� ,���^Z{D������Յ��'(��3�1EX\d`$}��g:�AX50	�+3cv��f�S��כּt�wb��TvM3���J��4/@z����~�e	�Ӱ�m	��r�2�� ���o X�dV�
V>+�Ӯ�I���93$k���E�Y���cB��D^2쑯���G�ĚШO��� U���Ɲ�5�NtO�WF��Q�!�ԒvsXL��}B���a���,��u����ZR�oFc-�U�0�%���^,��_�����$�Lܠ������
.�g�'L6�4�ͩUk������r{��8�_:C[�)��}"�K#���s���Be�s_=��2��vtcwNo�"�A���K:� ����Ҫs�W�D?�°9���ۿ���3�/��!-�R~�L `lޏj�����k�����������Xbs��<�:�T��ΐM��Nka�b<�ᲀ�[�A��;4�<P)+�!z��J�� 2���b� �5/�m,�(k�B�G8?�n_&��W���:$Z7kÝ~s|��SZ�~p�O��� ����H͙��>��ϩ�=ٜKDD�����5�V���10��"�a+�W�*�t� Y+�����gzX���ϴ`+U��+�%I�I�b��
��c��-6��s�.0\���	�|�4\��.2��O�#��B\$�T$.v����4���|}����m<ȋ�A�����#����#�Ɗ�y�Ɣ��Q��]��ρ�cZ��d7t����Ǻ~J��̓���R�;�Z�q+����R�φ�iD	|��N�w�*Ӷ|8�2r�7L�Yh���n�v����T�\����_����ch��A_E�k_ٺ��`(-u�2�e�`�3�-��Q:o���tN�RQ��^-�\�jkd�MV�G�����5U���g�.Y��O�6@���N~(gM�R'缲�JT��a1�Nk�c̊Oi�G��73A��,|�N/�}i��A��ay��&`!(�r�����u�T]Kf�`WY|���jA����;v�]����/��/�2LzNUr~ZO0��E�RӨ!N�w_Uz����;�x.b5��t�up�GW<[�]Mb_5<��FS+����O�"
5x���h�؂��Ma�p��-,�V���}� flV��qtٍ:���������c`r��ri.,G�>1@z����8��%�<����?�GT�q�%�v�X��A��h�6�]�6��v�a�y���1cv���T|5+���s)I�o K�&�*��؎�x�oI
@��H@-!Kb���v{�_�a˫߽T2�}�猔�H��ah���m,��I0OeiI.9��=�f�I�p�)ӣnO�_W�$�h۽�O�$	�v�ú���r����3j0ڽ�Il"��KK�?�ҳ`ABa�������W�_�^��{��^���=n&�w�3Y��/PK?1q
�{�5~.�a�^�J�80��Wi��\1�tw�G��[
��Jc�a T�?q�!��$�TQ�n����fG�et$˝q
t^��bUрk9!d�3E�}�akq�c%���󋾫��]Ӛp[�L-I�&��FN��z�8���~4�_�{.T���zׯ�ȣ����+�ș�x��nv�@��X��/e���i�{�1�?Žbs�о�c@U4W��I��703�7tM �3Ĉ���K�{*D�7���;A�YP)%�?�fܶ��|1�NZ��N�ڦ��
�/��<��rZ�`��R�xf�?'��&1����Vi-v����Y��S���q�Kř��"Z\����@56*�6%�N8S<����e�n�%ӌ 3����fٯ�X���F���N±-�@�_������?�KbC73��J¾O�y>��h��ᥫ�V�W�Aы���ԩ�Ӎ{揷��'H��K����z#�%�3�RS�����F+Ĳ���4� �#�s�L<���SZ�t�F^��z��s'�X=Ĝ,��g�{)\)�bu��`��.�����B��]�h����Ju�7P=��l�����_1�Ԩ:~���L�l���%�ǹ8ңS��Д��A~x'GJ�=���GR3
�P�~]
_j/���G�SQx�L�XX��aD'�(�.w_�PƯ!S�_B��V�b����Q_V�E�s��IHu�ٿ�< ���W�m�ҿ�.-���Z�՘�~���z��z�T?��D(�@���G�'�����*+�2�?�?��1hU#���Ul�]���/��	�:"Nɲ��v��|mɝ/(�����9�kg��w���y"�N����`ԕ.1��E�r��}�"��WW��'��p}�E�Cg�E�W5Y�%�9^��~��5�U7Vfn'��`��	,>]�+���._����>�I8<�G	G������9�W{��ܶ]�e�%j�o����k{uu���q"5�P����͋��F@N�'CgE��,5+�ޢ/��X���NO�����za��z3�_���
3��CU�M@�	EI}�ʜ��&@�P�x�}����E��^�F֥���b����4J�,�jn�S$تjHo^�1!�Û����bvo�3~�lî�)�G7͏�$�~;��x�E�!����"Sot�e"�e]c�����`�B�lZ��x��`1��$������jtW�����p@�S�|���f$=4�G��Xx\7�i�\+�zM���0۔���0��:��f�uŉK� S�'�Z��§�(9���D��x���`]ʭNg@B�(�1a�⌟~������aM�����/��r�����Bf ����갘��n�- �R�3��.Bf׍�%�)W}�!�-���[Uq� �	�b�ä��ǲ7�HA�=ӎϝ��R�q��OȮ���r퉥e�I~��Ğ�e����T���.$$�[s�uB�\6��j�Q�#,��O��y컾��� �Q=�W�v�ߔ9t�ǤKp�>�Rk��΍�4�E�[��W���9����y��Ni�^����&���&����6'���ӊ$|�5qy`$���VB>�ф���~:7b<ݍ�Cuf|��V����#�_��� }���u}X4oM�ͩt9UA��1U,����k̊�C��h0:�>����5���*b�gl�?PE���C����g��>a���~�+rlx�Ŭi���?ܚ��Q�&v�B����Y?��$P&b}*@O�X���!f����$��̋ѥu.�3��Vj�T���a���<lQȳ�5�7�<��h;�;�f(�J�k��)Y�͗��z� )?%��3�8�(#ŧ�7�A�+KD���\CX3ڠ)�Rw�,7r�!����z��<�4$ҫ��֋%t�}��td�k����f
�<��s�yc]r,A�x�j�y��s���.
~Q���i�PL70N��Ae0�%@ƉC�<X�)�?�[Gܜ-�}s�#�~ı�]ۤs�N�u�ު'���%���y�!T>�y䶾i��]J���h|���q��,�W����I��4��*2I�{�
���ȉE�]�vu���T�f��-=y!�bV�x�tv���	�;�5�7Ƀ���m(�˲<�q����b��uim��!wxY�Ŷ3o*D��1x�N!B=W��$M5�H|ϝq�{�1r3��׃��Rs���;2��e���OB�%=h�����3[�~�G�b՛���C��]�ɬ=�����
���$,�� �Ñ8�DpnD�I�a��p�2�<�s��lҭ}NX�XD2�Hs��X(b]�]�5tc��ƙ� '#饩�����w5�ӖX�c�%%��M�2g��D�U[��uO]�d�bL�5��� ���f�pي����[��t����b"���b��
�s��z̞S�����%y���6�w͌�84}4j�P�_�&��5W5'r�G��]Q�9'W^wL ��ϬC.j�U/wug�xE�զ���ly��'R�xBLg&�/5�U�Fŉw\u{���6���0kz�2����8�n��ɽ�<9Ш
�'����/_/���բ,��\zѵ�%M�]U4{7\���q��qP�@��<�ZUo��=�Y��O�dP�X��	����sG��cI-�?�0Åq�*�{[`<��c���0�^�%[�0����+��A�9�|2��sCWBP��Y)�S?U��sQ/ؗ8��:�1�jڃ_�j���g4��m�+q��7R�3$j����������X��=R�wx�N�p	�7�=��շ�WiƍJ[�`;nF=I���%�^�O�`#H��W��m�����Sͼ+�]��w��l�����ts ���Z.�[�f ז�5R�u��ʝr��K���_]<������T�{�>x�Ch�o2����ڊdL�`'T��&mDd=1���%�L5�/�������rX���2�y�E��$�:�q R���\5�S�'e������p���I��y��w���.=��#s�w^�I��U��ά��
�QKf+xN���Y���lޟ�rOH[�m#8������x�?�)�u�1@�{�2n����A�k� y�["�0^�ܴ�ڄ6���� �S���~�jf�õh8���o��ٹB+�ǝu�E�=�~m�A֫4�U���K�8�l�D�CvT��G�dչ[Y Ɯ�
�T^����"E�Q�%+�e����d>�ݚ_ڲ7���N$� � ��&v:��d�m�c�,�wW����tΖ2�_�PU�ߟ�_�"�G��Jp�Gտ��m�\-M�w��T��?k�ň�++���I��O�Yv���5s3��S��5ǁ�ԗDTr�?�Q��YA�?��3�ZC�ќ^s��/�5��H�FiY�d�������ݹu�;0�\��v;�ZVI�=G~�������]��;b@3�*�3NP6�Zp<#�j��u�Pg}*Z�,7p� <�����NFT�_Y�1�捖�eg�׶�9�c�mo��&� ����QR�l�H]�58z|��,��G��7H�D��VB����jsΕ��ş�F�H�CF�6���q{�'�'��2e��kf3"��8��Ʌ��������۽\s�������٢���e�$/�W�9'M��܆�.r'��	$ث�pڒ2��`~��� �����4^쑨�t�3�D����Yf���8��v�k���Sո���L�RD�N��
L�JQ1Am�֫)iw[0�gw?X=�G��v��B��Vn��9%���Fgjd�s	�6��۴ΰ=�C�֒&P(��Nlw��]@�&���	?K����.�[��C�3�d]g�i�����TOR_4���lN�O���C��shwެed��ѱF����n�{�c}DŇ5��]�9�F)�:ee�Vח�NP:���ޮn�g�~���4ݣ)��$c�*�*�1������� ٟQ=�c]�郺R�n4G���zgm�VFrT=�_����Ϝ�V�����n1o��[r��w�M:�ULb���ɋ9>[����)i=�_��3��TyH�T�k�,^4M��O�^����z�K
��K��Q��kģѰ.U�N�y B���4�8�zDr1�C����*ED��I4����W�p;-V�Z~ȢO�[���Ծ��Z�����8�yG�w�33�V�Ճ��^�jJ��P~Y�sz�E�CqSX�t�G�	������a���=H�П�>p��N/�5Ͼ|P�:��Ƨ:�M�4k}��`q�L�K��_�H�7�����x����;͔"�ҏe������ǃ��gc��M��Rs�S�_vvwtVlW�U�K�y���;��0_���V���-A�a���o������D���J͸�� �������6y�S�"�23��#���'��G�Ta��At$�.�Rgv��?�D�SZٯ�����àЊ�N��G��0��z@����	��q��ij�_7�9��u�����_�^��a����a�=Z��P��`7_�E�D�Z��ы�^yq�~Q|��A�"�~�ci�1M*eU�.�uC�r��^���4@��d�l%�}��/f�YQ�B WI�s�-pp�E�ȹB�����'��9���TbP��=M������4�-L�X.�%�����?k��z�_�-+.��Ց�g-i �xs�U4���$��u�+U5��Ʋ-%�R3��7C�����7r.}�{���k�z����M#�RQ��0��gV؁���o��j~�:�S�t��d�ӆ^qނ�f�cBvtIt��(��R�5���D+O��dE�--�~U3�w�cT�x}x�
*h�O�@|����KY(/�r{pH%-�~�PO|4o�.�qX\i:����g�k��6:g��GnH�S����9.��3�%9�w��5d��1��R�e��WvZ�1�i��s'i��R��o*hüe`�4�<�^YKmę	jD�����I���z�#�4f����s�=Q=j�)A.�0���!a~��H��X2�n�fԦg&��b��I/�L/�Y&�Q��B15	0���iy���,tc��ϟ*c�yD�����+<�z���/��M,]e���
C�r&0;�"�X6|���V]��͍�Wvχ^I�pԫ��A-�!8�E,���7afy�"�J�X"�5�u{���	iY;v u�Cc����Z����_����-κ��	�;���y�'Y�ᖔs����K�[���P���)c%�ۆl��,��V��q�m��!0djb�ے�ȅt��T~�h�FXn:l_�`c�s��텊���ז�^h�$�(�%��V_LH��]��3������v��>�m]8I;����Q��Nb�;���1_��9�Ga�ӓ�u?���wQ/L~;�qZm�9��F�EX�o\f-�p5��Ȅf����0Q�KMۋᴙ���>�����쫥▿E.J�(qW\��g��JĪV3��[�QQ�h�QeJ�����,��E����1�t(����g��8�9rv�N��@}��L�LYj�,۽14�ۑ%�{VlŮ%z[���A�3��w	����
ޖ���ofDo�����8#3��Mv ��*;�/���D���xW���h~��2Np �"z�$΁��P���lB:�C����Put��m<:�Ւ���?&��>�9��Ҽ�HOy*�2-Y{{?��[�c	�C�ʚ�_h�(� I�EC�n�x�Q����w~���.�F�M�5��F ��F*�0w�bsm9��\�'��u�/u1�T���(�S%�h���cE�z��-�����$%*}߀!��^7�n�<+MW��|cB��+��j�-��6��Ac��UwV�/�o���r���"$6�;z��� �5
\��Mh�3�#L2k1���k�;	�I����d:�ӂ!�r쭅XxQN���.���f~F��@���Ȇ��;(9$���Mr''Q��0$�n�6����N5jo�f��EW�`u7�0��\�}�� :���B�Nʅl+�f_��{z让�]�|J�!gW��	���~�д�ݽ���>ʪf���A��0�%9�Ftn��	�LLb�N��R�c��aN���K�%�6�
w�"]k�w)Nv���Y������/S����^\|k��P�|n��t���'�3�x�T�B%�	a�ML�Ok��J��ޑ�M��Q6�9h>߇�����Eqym�ZV5�x݆L�f�iV�E��Ɋ�Q��VW��h�+��S�>+K�w;�_�O��d��L�K4���:���ۖ	#�*��a3���1���{�H��.�����uΝLlo�/��l�w�9�T�G����?q�#�U	��Ug�nY�<��nbA"�N��A�L�5_#B��������C���zan���S�#x��h�y�| R v/O�1��}e(��]	�Zf+=��R�=�j���rC6)�`t��!�3��ƲB(�]���~5~�5���!�=������V!0Cm	�G������Oy��j�6�GN~�Q��
D�fxE/M�7���; ꞌR*��S��3p��b��nG��[WH<�Mx���a�Y�A����r�x���{�$:����~�[�sO��h
{U
���ɲ�fE��nN䨽��e,_h9��&F�Y�vc{���ĳ������	��,�(����uHL��Ċ��� H �}��И�0Z����IW�� �G�Z�.�\��o�R�r�����B�Cnp�l�x:��x��|ڼ{h���<J?�������#)�M�P�!Y�Kh��~B�wC���A.>���&l/�SY��?C*�x[�n�*>R�3���O��K��;�$(�n��鞒�Z{j�8V'B �oi����l$�Y�ZK������uI��hTR��@sx�v,�N^`%�q�=��L�)}����\Kmt�"Ys�sv'.u�Z���f�än�d��xQq��z�F1�mr|�wV)h����/�/f_���ta;�9�L��[?9�l\�)7pP��D�H
�Euİ�A�8�Q�6Q��ɕ�e��M�E���n���Y�*�T~f3��¯{��)zÅ5���\7�rC����=�T��K:U�w|Q z�,�a�q=���G�`���{�zim����e���h�<��9��Z����@��ǌ�#6��F��9c%��;~_���S���b��YHP^˷4��[ذ0�RSt��^�� �#O��I�@EE��5��i��g��Q�>8�W�'��T��S��OЦY�pt�޴��t���'ݜ������S;��U�\u��ޯ]FMB�B����B���~�r��g7��i͵5|j����"�æ��ǔ$���,�����5޵:0ګ^r����B)+m�CG@_����K8Y�+O k�*����?�GP����QH���	n��wM�	[����9���+�I�&̕m�J��P�z��L����;�Z-ڟ5Q]^��c7����8�9T�t\+X2�t���vAO�H6Q���h�9��rg] ���K�{���6S����k�/��Z���\�=�l�/*Kp�F��-���>�}=d�R�J��B�w����]d��O������*��}8�E�D��� ���is�7 JpwЌr%2���=��f)0��a�l59p��n�JusPV���N���G�y���Cnv�|���47ˏ��RP2+C���7ī��O���bu6�F�T��D!k��/�+[!-}j�4���Ε�
 T���8�WV�4Ċ��t[�5���r����w�#���Q�2��G�DHRC��l=�vT: %�Mͺv�Ku�8@р!��q�!�C��v�'���N�oM��A����e�������`�⊄���Z�M��k�9 ��o�W��M���k���Qה�/��� ��&�T�Q����(2>#\�iWEp^��Q
�z�Ԕn�Y�n|��`qy��㯗�Q8��_���C%�z#��3��ﭣp���*q���~�Mā�U�/�/��Y$�����[����?�cǪ	�i�.BD��.1�e��t9�(�_޿��A`3�גI�@����.ƀ�N(����_:C����w�i�t�#0v1����=S��;�n���Pń� 1�ʼ�-�2$p��h�B�؅�M~iyi��^�AIL�Ƥ���iq�ĊN=	��ݍ,��rm�ϋ��opLS���v /��t�;{���!H�~҉\6	c�y�yx��pa�n�Fx�M�H�ӽ2�;Ev#�s�E�Tw�i�M������oD!�b�A��$�v�+¡v���w\/�����Ф5t�LHj��k����3J+ޚJ����M�'���K�'.������i���2�UC(E	�,R���9�@��T�6�3�+r�Vޫ6$h��:DL.Q郧-U�y��ZQJV�ִ��à6���R�v�9��v-�\��e�Oڙ�gĄ�t}��̰���ÃT}RD���Š��6~8y!�e��WJ2N�(^D���Ǐ�="/�{�Ya3$���g0r��v+�$ч��)?{FO�C�I��������?���FȊ���t�r���ݕ�$�fG,�ko]Z�+9 �'y�S���@H�������9�]��X�K� ��I(@�	&����h�ˠ����y��U� �`�"�r�hn��<��֢"�$y�]x}6�Nt����3v,9��B{,�qmAp�?i�O����e�)'��4P�@�n��/����@���x��sc)+�,��ݘ8�)�������^��Q�=�I@� 3'��vO�ѻ?�Y���3E�s��6��X2x��?����r�Z�pf�8[��ؙ��b��[�d�M�k�����rt9Gg.�tT:��uym�%�w P-^���LG���\�Qn�ʲ�al�5��l��@!�4P���ɥ�z�r������ŻR4�٠���Z�Ճ�-^��"���s锥H�����e������ѳ�Xuq��%�ͬ���H��sC�_WC�-6`}Q[,G!���Nq�\�zR���;�h<�@������U�c�H�;�دS�L��u�����"hC��4֎za3P���=���آ�uL��[R״uP!���L.rǔB�r`|�������e��E���J��@�V�����V�|7�����4�ˎ�ƶ_3Q�&�f�z]��&�2~���.�?v����,"�����N%�?Ū� 5�L(����g��+=~"{_qpc�Kqf�����3�<�V�8��F�����=�6��$��.ٖv��h�Ѧ�p���,!ET�Yq��fW��4^d�Ƌ�ܒ�n��>a���W#ߟbG���~}���#oW�S�o������ a�=!W4@��YS���Z���9ؠ![���CXU7�#z�4(7��6�l��BbI��:���}f�7�2Z��I�0������5| ���V}��UHxֈ�����W!z4m���;r�5�Y3T+��m p�q�n�����~|N��ʺ�?��)J��Nd����ޒ6<��o.��Q)������; ��������U�Kb�<��MF�R��Y�����Ț�$F�؄�S9�aO+�JՑ���$ �$�7���Q	B$Va"��m�Q��#�J>�]j<�L��I�-]�h񞡤���k�}-�-D����53�^��h�{E�.A)�ġb�t8���Â,�4���N���-��3C�u���xvCY�Њh�Z#�#U�f�*0��}���|`�`�ޔCR���\U�/+�|i�SΌ'�ǈ��o�����ZX0��V��s~V�x�S����A�֤�Q�� �޼I~Ɇ�I��é��b��X3�AMe98��Y���A��m�g�?eM`nRJ��j`}k�
���m��N�Z��PpzV	0�����*�yc[�����a�2�&G�L�j�2o�.���h�}䩌R3�'�ȿ��7gK^�A�ߤGP�Qd�NFV�	@r�ǵ����y�Md1�@�|�y	�+�X��x!9qK��qi�����k�����<��ɔjƣ�å�����R�ޖ����C�FW2�[�h�e��n���L��We�gW)*�و.�S ��w�4��h�ޟ��G�X����1�v���Ym��6[ZϋBx�^�!/�e���PsU��弰 '��yш�7��Xb[�����Aq��F�(���%���b���p�* �s;$�����dz+ZK�4b��'o>v���VWJ0��c�q7fkpuʺ?$.�Q4��������f�"���Q�*:���Tr�	�b�����:��"��#x�d
)�e�Z;�m�L]�� ����ZC���pK��+`����mbD����v�ޱ`�L��?2�՛<5�`�!�,��8�b�[F٪-c��3�B�7�%]�$È~[w���+�IZ��O���*�g1�op��<��y%^I��t^.�q����3A%�;��kT��'>�&|<��	|���N�X��I)܆�Gd���c�xQ��#P%�`s'��g�c|�[f����5~$$��A¥�#�'��&|ו���B�d�E�k��]A42��?��vr(�[߹׭�n�=D��j�t�&���ɀ0"�	ʒ�ig�^jja����`i��@H�5�w��45�[u�]ia ���n �U�o���)=rE�\K�!ۀ'?X����53��!7��F�k�fV����"���1�iw���p��c�M0���%�\�9B�S��i뛆���ų��pi���?�o����A-�&dE	���*	���O�;��0��C :�N>F�b��/�L�SH�&�zs�:Ϊ �\GH2ОL����f��q�h����ұ�ڹ���)���ld5%W���U�4l^�zG׈S�dݾ���,�ʒ��ý1˝����m1��	�.4f�ژ����^ۇg�C?���y��=3��L}�:�tls;�)_1q�n�i����G��{"�/�fV.���+1}ii�:�-�Y|	c�N�!�z*32�p�H4r�/����D�X�l��8���מ����3�z�v���P;eI��oI|瘘��f�g��dd� )f"Q è��Cc���X"����q-􍇜�Rr�d������HB�z��k��j�|�6a򽣔�]v00���TV�+IBW��ɰ�<w����@�d�v
�tLq����04�s ?.H	�1�煟b�1�KW���A�u���}3�Y��W��ɣs�w�%j�e缻��'���O^xNI;-Ϭe~:�;չ����A7ׅ�$��a�y��:<l��ZI�g��ы�yKt,�(}#ʎ�{h�����D����AK��;�	�������8�0"�cl,