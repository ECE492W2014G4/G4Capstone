��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P��v�"<ߞ��&'��k%P碶�R�ӣ�sĞ������FY&�E������%	�����JO�Uv����0Z$?�`/W�ͫjP��{��Q�K����W�Y�\k�;�t$g���9�l��^t��(.GH^��%�N)�G��
�;��d�}<�Y�>�s��9��n��;�G_�X�Eg[4�s��4t�n�K�1{��(�����O��|�-��TRl��Kj+��a�o�G4S����NM��9�|0��dU���6I�Pe�;����l@ō�Q$�$�0��V��ڰ�ƾ]�h��7N�?���ǂ��]�"��b��'��?��O�������"�U�5�YT ��r)=��3=�Q�l-�O�%��K7���[�Q))Z	s��1}�~��_|�feCi=�es��桝��﹄��+1��at��&�ϒ5p�+A��Nn8�&�St��������43NN�����L�rF��)��Ku41�' �!��"��·a9�1Eq���k}�0�x}��g��v:A�{�cV("(��SK�����#��- (�/%^4���e9T(j=
-�5t�S������4�O����Mx�}K<���Z�ڸ��AE^Jsvz0)���5f��P�Rz��3i��@x���U��?;ֻ�ڇ���{Ʊ@�p�����Ph���Ք!�\-!�.�Ĥ_dw��%�<��E9{��Js�h��P�w΍J��/�Ab?Q�	D�K��?�)bu8j,�i5]��}\؁������|�J'4�C¢��3(�%�Z����G?���H�`ͅ��{5.L�w�UC��e� 1��YY���"};���@; �:�R\dҌ��B�7��c�<��ʧH����ב�%�r�2D����3�>+ňϖ�A�? 7��mȤ�3 ��PsX�h�D:�c�*��^���.�h��m����Ċ,��˽�
�#��H���AHv+������T@��h��S<��.�ޜ�޴��i-�E�|4��맙���j9ܔ"G]�0l��]蝗�lMw��(�ds[�����	�(.��\��:)�b��sy�6���m3ܩ�}�G�� �v����i3�� #���;��sH�A,�}�*ܰW���F��2�}�CF��E�7
�b��Ktm�u��>ܵ،&Y�%���wC`�}r1}W41�d���9Q'��x���~����z�MȦ�j!����U�_
��+��r=�74��o��@��hg�z���3����5J��3�XAP�r�w��S9�.w~�t�j��g��#(�}��5\GIm-�!/�Ȩ_��sB�?�@��	G�q&�y�͌8�tq��r�<��YWJ�MF&��{mQ~j�e����,��t�㋅��'l��\$�� <:���!��M��u��,��n�x�3FEڀ�Ҿ����@{Oy�'H�l���9����U�O�lE0�p�A���.��t�#���9��Cn����B��n?{�:��"�Wd(3~�?�1��9��c��Y�����j6�Ъ	k���$��NF�\�m�.��^l�+��4��+��b�Ll��&��tQ";�o��I���uO���|�<����|�]�sv�Z�#�����~�:����jk�2��=o��Vȓ?��WٯϞy�V�KǕ�	�` 2�IZ{�6gH����V;�1��狒��آ&'_���7Y�m�h���v0�*�59Y�5%������� 	�����B:��XT��7�(=ee�����q�	m�D����(ʊ!��x��촬ǝ��K��N(sk��;��e����&dF��@n��d��U8;�~lP�V��V
7��J{�HO)���L��J��a��4�Ur�%�5/���vj&A/��[ձnWɩ�^�T����V��Ӑ���p�R�t�޺DCMC��Ҡ-�ޕ���d�H�(He<��[$��s��W�\�o��[��_�����O�-kS��!�T�ݵC����qIW������Pf�8��M9~�J �&h�>��_K�-B�X1@f��zmiB�u����W�V�(q�3h��xh��}ڴ$盾��qZ�r����1����!�`_�G&��K�cru
v��P��؆��g(4f��$�'�3�[��N�v����s� ��uj�u(V���۷0�x)r 9���8�~�'bU2�]�	���vu̢l��'������_Z�_�pL�b�_Z��B"wũJ������=�P"��J�<�:�L�tI�^[��(�?:��2��N���যcr�pM`�5�]a����3b�"t�݃�]��fl�d׊9�O7����O�������8� N8D���wM��!u �8�R-�ќ7�y�j�Ki3Q���
ֻT�i�="�V1�;� �-����D��,�V[�mBz���E��Kq�&�1 ��P9���r�яbƐ�����:q��q�p�BA�32��e@>Jp��f�ҹ�!>�	����_c	[ǿ�T�|�i�c�l��Ȏ)v�><�I�v���t\�?=��#U�ob��M��ܛܯ�uTm�+e\�{ɏ����B��;I��*�b&a�̔Ed8}�Y~����"��D���@��[[ܛ��p�b5�"��ڊ��b˧�G�t��'#Q�C+���d�2���a�-�K�N�Y1�(���|#З�S��V�9�6+q����Ԩ�5xw��^��5�V��IF'!��dy��W�WT�|��hW�.n]��!�KK0�P1�����*+>_��D�.o;aY�e��فu�?�h|��w����hXn&��$�S!%v��IG���<�֒6���ے��->�rNw,�)�R����wQ����ywJ���?gc�;���;q��/�"�
e��\b9���L��-0u���F	�O�g��R��>����;����׊}��)2�P%܌�H�e)��K�q >�\N���b�L������z9~�D���;@Pn���)r�V�jǦa�AW�j�> �G+�X�F���W~{�+��Ma�0Gt�R!��ᨛ�֪4��=]Y�6�HuI���;��u�ѻz�:��K��#�ϙL甂����b�jkb ����<��Uv}�n����ZZ�i`'�
�ٯ��[�^�kM��1\�b��x߳q[Q��m��Sh�p���g�\�8�Ѽ��Cﱰ��7q�`cb�w,C|6� \0�{�2ԋ?5bY�Uڝ��~�0� b'�~�Lsx�e�b7���'�oP�������7*��={�0�p �"9Ԃ�����F\e]���x��@�g�.b��Q����p��L�/@��c|��0���mH����A������@>�3j#@3�Y�!v�޺*�_�o���!0�4�/�|���3��D�3����ԛ��Zrq��"��S�%Pr<���0rm�R�����V��9�Sp��k>��gy���賊�4|����ep-\��d2q�]�MN���3Ɔ=�}XyN8Z8z����*���E��R��+��5�����ɓΛ7��9���PP�k��ל��;Nm@,�$|�*�� �`m��|�l]����8+W�cm��	(��Y�ʬY�6���"�Q0j>i1�1LT�e�w暮OTOmOUt_-qɵ����a{;�!N�cgs��ݗ�H��H�����C�H�#
�u�����V#7�W��R�+Jve����(l�EO�SD_w��,���M����We�*�X���,���w�v$ߎ�R�������0�m?<�M�yT�C����tL$��fG*t��t��7��?L=��mw���^,.8g�R��5(����N���}��5*M��A�2�)5�<"i��x|������oBp��Nɸ��$4����b��P|`��8ILSLRn7���$4���]����cr+�zh��D+�bo� �o��Xʠچ_���ÍyH>��NO�]���I�rw��ML��D��P.i�}�̡8�5����y�h�s�n���m��BQ�tAS��sg�w���d�[O����_��[��/$6 K�t���Л���t ��ޖ
^�{��W�����ʳ���n�\�!鋉�f�Q�F�\?�]�Ê(\Ѐ;�ɺ#��7�,�ppB��ũ�*)���-K~������
�To'��9 H���C� e�H���8I��_ʩ
������B{�b_kco�:���9J��wi�����F'�z�bS���L	�=�_� �qc=�����3�e5��
�J�r�;���[�
p���I�ws:ϼ�4���Bm��u0-����0�,�`p�'�4p@���%�o$/�ҁ*�ܼ�w,-+�Y��� E�����HWJ:iV��Ȍ[��q�{Ib1���:��s����%,�uYw��X6��]�a�4jfr��{�e�j����{Q��������!~��xsV�#�I=���U��_������qTz!0nIzP0��Ŕ�L�E�%�'d�kLU��uL���W+U_3������I�`�$s�{D�l��+.�#�R�&��~f����1L���x�_� ���mo�B?K*=�4��S�s�+�b-��]5��N��#o;�5��#���7O=�}�oz�"���и�6�3�_W?Z�X�������^�����aI�8�V����"r�oB |!��!q4�,�iɅH�%y���4<�����