��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�"��F9s�`&���a�oq���F�g�O�]�<ݲ����eCL��D���{�5��8̝DFI��Zp\m|Q��
�}�6C���UnF:<�jΈ�2�����<����sf�k��,jڙ�����2��X��Ss�HL��	�������+g?���N�Ż�����|�v7�{M��VNB
��Rs�゙�Ld\��X�'��R :�J���^�����kMkx�Q���3!P}�e���Z�Y?.�U{�RP	�)��lI{tI(S
7ZF�W+h����@��	|.�0_�[D=?��\c����43�Eћ51�5�H�����v�0��%�͢,R�����i�[�I�Z�$r���H}Oԯx
B��~�R�ޞ�O'z�>8~�ݐ]���<1j�
J��L��{�S�E���A�v�Z�'���!`��$�%�_�]�鈺�Y���':����tx���Ɋ+TV#����7���V���%�l�gq�ۭ5���Ii�����9��̨,�d�(w��!�/��:��Ƚ��Q-����]`�����V�Hſ*��>��HK(4���hÑ`_�щ�`lL�q�$�Y5��+��jן܌X�S�9Fj�jU�)��I�ms)��Z]7��2��^�a(ZW�ՙMg���埏����}����o;��E�RpN�f�K>���t�d1�?�FqE5�Gep��hI2��O����[�>'�e;�_;Ǒ�K��X�o��v���p���6+c\���A�s�l_�� � ��q �ژP$v���=��rF���i����EA`�)��G�1_�(Q	Ɉ��qt]�̰��7B�dQU����������8%�b�{��-��9`OP������G��zE��v��$��=>���������|>����#��ɯrW^b蟯1_���z�/F9�f�����WG��Y�����)����&b�#Ɨ
󞈿��FE���>|�c{�䘄m(��F����YAz�y�.�c5M�A[��[uY�ؽ��Zi1�AW,�9��� 6�H}��Y�a�hwE9�'�|�nD��6!iƘ���VƊ��i 4��`f*%������3t�w�=�L#�"/z�R��L��G��HZ
8b���f��<�^q��K:��9�%�Iw�E�[L�U$X�-W��>9.@�AF-�����j�aT��[�"o�D6&�68�����3Yn~`�"fq��#����p��C��dgm�4��f3�1ot�*s}�g�����	��4`-P��.�4�I���L{?�(lx\Dh����t~�h򒄩c�ttS��]&ڙ����c9љ\c3�'�� �����H�"Q��#����R���'�c�?HVH�W��ʁt�l�=�ĺ6˱��[Hx`�1�TA�>Qbk+Ŵ�,w��a��%]�I�"�rJ8pj�Vz,���<�&�%�ve�xM�9O�O��Y��:��W���x}���~)�Ɨ�Yٝ��t��dS���D1��������E�x��O�2�!�J���[�@9��Y��U�Д�B���!�%YKhH�Y{�W8j z�����I�>ɯγ˄���4���j�5Ҝ��CU��>Y��vT����o���J��������]�h?ubQ��~)����SKWH�@��dZ���e����g ��B.�3AH��>�t7�/��-k�W��a��l��ϋ��UM�������s�}�
���-��7Ԧ��]�a��q?�ʕ���x�0��&���YG��5
��?���mG+��	�¹NE��x�O�w�y��A꒨�1���|l���n?�>��"I5��#�@��(��C@�L���X'��c\I�WyV[��}�b��|�O(k���B�,-	�VH3�O.&Aɐ��������=Y*�-��D�:�nw�4#����{]�"JQ�w����8��}���Ul�1�z_Ԯ��ɖZ]X�^*�@�ׯ.���eΧ�p���*l㹂m�]�����>Oe_*KC5n֚������ꮹy�z�D����ve�D6~�J��J�g��� z��-���;8�2����K���Ϯ��z|�)����X-����6%hfX��>��M���:�4U��u}�)V]�(j�����<�|�ʼ�b;/x`?=J�T�B�}��*D���F8~�,@�saZ�_�|�����|���S�7y*�plŠ<�O�z�����p������G��x,���X�_��uh��ܴ�$�[:'����Y��85O����\� �	|�ʟ�.. )zn�H��rzX8T��f>���ܯ��C)t��e+O��C1�vt�a���Ȫ6�`�����9l�#k�>`�3"x#�n0��kʻv����'d���R@i%�����4��yS�VW�b��z�]�H�-Ub��M������J�qnNw@�e�˒ʥ5�� ���3��n�u��ƦIZ�N��S�plIK�y=̥�p�q;j�>����H��5�y�SMd�o�겣
Bkw��pw�t��_U�8�nSƄ-B!�ɯ4vE�v>H߾���;�j�sfP�vF�ؚ�į��0f��/C����7�C���ֶ�W�����&�گj1%y���#�N�y�;�O-��G4h���ڍE�=�p�C,�0��A�j��V���~���6�+�r��vv!����*�����Ɲ����&�݁Lf#QN��n	A�\��̰�V�r�I&�f�y���z�.�5�D]�ݨ���Z�J�*�0%k�_�]`@����y�C�9B,F����
�S��N P��Y�×p���a.ؤ��-m����qt�7�i�j��L���)`t�#֔ɓ_�:�SO]���r=�⥾mX㵓��J�w�?L{	�Ȏ��C'�z�ZPhS��8��Q���0���d��a#�����|�;�R%"��wA�W	i�.X�D�7��Ռ,rךJa�%�A�+��9��o����%�fz�x2��a�]"U�!"#� �>2��*�k�������vx|W|c�z �Q����������w�|t�V^��WúҰ������F*���i�z�&��K�gb1U��7<'�Hx�b�w{�c[���H��F�6�QR�B�h,8L�8�E�S�?������/H����\o8��U��O 4��ٙ��7���:5Z��)�̶�����j���<���.�+�4�2��=:x����3��Ò����� ��Ǫƻ��냮c�`�X�[/Q/Y$�x1U�9#c'd��Kfp�M�o�Z�P����恔�f�%��G'�P�@��HH�u>�(�C3�T�f�y��Ԡ#ػ>��m���ĬQ��I�J��B\� �4g�fAY��z":��a�#)�,��_�|��~\��4B���[�����"�Dr-�P�s ,.��F�V�{l�Y�Y���<4����5۠d������@a�YZB\��5�e��b�/XS��C�����OX΁6@��>ۼR����h������b�.n���I9�){EY��3jH�q���>NCJ�6,:�Q}�A�B3ى(��"�W�b�˪����?h���+�S��"O��Pz�XȔňG/˥��a%���QZbK���\�!"�.0{��z�^�m�>r���䛇JxN{���{A�`?�߿���~��@�l�Ƽ�(d�9�D	��O��[���N�"�_5	,|��٬�L_bT���J��>`R�f��V~:�׊�7�3���G>�Jz����x�n���=^8:���(JQm� %k4>���]�`�j���3I�3^�����4��E�f(�>I�����l�}�����&1���썧�_'d9ɝ*�LoQҭ���d��+D�w�<3�HQ����>m�$#C���BٖCj*����(��L2X>���'~h�� )��p����۸��p�ͦ�x#t�Z(�-��f@����ǫi���XF��b�YU�r�;�Dc��΂��`"��w�����f�Q�"��&"l*��Y���&�\'�M`�:Ҳ���˿c������4�n�&P�[����I�����>���
��m5��ƠY��
3pC����ޱ>�/jԧ;c��"rl^iɫ���xH��g`p�_��D#���x��TH ͅ>�e��|�S�-��ғ��v�V���=�v�%9�uʊ9$؃o�W,�c�g��n�b��ڗ��
ZqY`�-��!��/���:��Y��q:\<�TH�C��#�v8��wD���yr!�+�%{c�p'+X����@i�P<���q~�ѿ���QCc~p�W�xׂ����2�̕�9��ڎ\�
ЉȾm��GW�Da�a}bݳ�y? �ƿf��PH�4k'�q�5X� _���?�@��g�[��#�v-r�!�VR���BO-���gI^*S�N�QoV��k��ú��K^����lAD�&`Z��{+�Wm�����[��l�����(�
Oۿno?�-O����e.�C�h��������W�?e�M^L������8�E�/�~���\��j教BVCi��xh�Z��e��7b�WPyy�
�}���o��f���].����cGV�=��ԄS��X�B�	��3,���6B���Lo���Չ�k���&�p>o_?{�ڋ^d��t���OcKk`6a��MՀ���n����ۣ��[à����O�F�ap^�hK}���[+�����������m?"�>��L���&�C�H�bvb�d��<H1��$v��ކRVZ��.���<�0�	u
���2r�<�֢���';���t�Nujc�@�7�N%� ��v�ֿ��lL��<�EY�ɱE�D��s��d~!�8�x�t,�5�����uUFq5���9�+������, Ѹ��kB�e��C�~�c
:iŲ(d � �U��+\�:2x����]�z�6��θ����O�"�V]%d~�3��,�d�X1�j�k2��qM�1[=X�.z��Ȼ´��p=���T�J���I2���"���6��#D,��Y9g�.hJ�Wx�����^�)ң���ע�)��J���a�+}��`������B[�]�v��V>��K��zt�GT�m�TI�:��h`/S,֚K;�@�u:/�nw��-��X��q��(fb���a��	�ő}�Ԯ7����vJrʥ����X�����t�D�����G���u!P�B�=��^rZds<�t��1q�C.t��~l- _���`�p�q���������ؐ����KUvZ���r$��O��&�o�Qgڟ�|Vd����-��		˲C�p�0�{C�ҫ�pq�t�����C�0�)���Se������FW�ʰ?�[AoRh��4�*>ê2�Ɲq��A���)�����g�ـo+��'nڅ(��xý��� Z L��ބ��1t�'	�Į��/nJG��>(�ӯ��!a�<_�e	G�DSd6aG Td8�Ű�iU��2��j8&r=�[�=<CP�3��������9~���|0?A��%)v��D!�.�yٜ\丕
��S_c�k3�-��6�h@*�&N̜a;/K> e�yJ��r_Nu���iw\Q���#{@��:���1p?��F��N�e�g�Qt��K <��:ԟL�T/G���hjUv�@Y6)�����p]��p�)/&Bwc9�" �SKL�S���لy��HK#UeM#�2dv�?uI 0�n,��wi��mOi|t�ON��ͳW�w}�C��?o�.p��v���	�n�{/�e�j"���Q��� �a���Lpʹ����(�xD��S�ԒŊ)��R��a��Rcta
�z����Gi&wD�{�F�����ϴ<7e$�2�Ua��\^���x��{QyY��k[�v2o�df�v�փ�F���שּׁ����]jr��b��
�(D�]�Z�~��Ư��R"�Pf�d�$��ֿ` ���&6=l�7��s4�K���V+^�BhJ��ۡg�m2�&�������N��[4K�s���r���Ә��j��ƍZQQ1Dm�i�}yU�J�%�_�^��ƙ��c\�?�O�ߤ�X��V�*x�d	g1�}��IV�to�%L�8��*2J��F�����|f8~��ލ��X+����p�hMx5c��=���
��bX@D�9��3u��(������if�������TT�"��yH�M����c��x�K���O�7:1(��@����-X�����O��A.�N�x5	��#>�����m���k�I����1x�.�L��,��ʎF��h;�0b�b'D����o;�N3pu��E��s�c�����\#�P<�Я5�w��_gf��ݒ�fзhk��%�v�2�~UQh��J�G+l�P�h��Щ�=����9�!Ʈ�:X�Oˠ}$����'b�6�8J�5<T�m�<�X��������H�������J��j�p���[�S�N��q|%͆G��@��� �����,c�Dҳ�Q��kg�
sn1�t ��U�_8;&��?;�!����k�iF�������A�&0�����v��[x$�+�G�n�z������k���&�J�ܑ}��d�ΐV����h��
Qo�J�:�|#��J����"`}V�_�<
Xyt�dSh�f� �pK"f������� b�O����[�]-�Z�_N*5�
x�M�!�%�2ԯ����|f`�|�@�>3(������h~���w{B�ը~F��o<�`���~�B�j�N�3"�C�D�=\k���$%!$�h!F���f6���̈p����*M�mѐ �O��Q�Brą��K=�`1p׀�g�)T��!��2�.\��?�s�L��(��ڀhg��=|t+���Nd��`
�CV��J-��Roք�����fD���4P�\�yj�o����k��#v�l�-�e���C����4�.�X��I� �ݥw�|06a�����P����,t�
����O���\	��S����y��F��_�Ԟ���Vn�7���f<�w��(`�#�f�����n��(��%��<B�r ��{�^x Ep���Q�����E��:t	P��A#�ɭ-�n~+m������� �M�n��³�%g8�@�2Y��Hj�mc�rz����ц,ԠQ�jwrŴ�m'{��)�`ּUUsުI�p2$��b:���~�S
��rF��_�^m��)���&��;�׍ЧN#_H �m�=F�pG%(�6�ֲ�,��\v��ߖ]A�`9+_�j�ȗ�[�r`��c- �2`+-��_��6�}':�N*$妣C	ڑ7ݒQ��)5���$����@����s�~�F��0�#d&��,O]��_z��]�7���P~���74��
y���l�[�F8��+�����ڱ���h����3�œ�������cR1��M�����S�:� �V
�5u�8��$t�m!/)�k��Fi���d}��.O�ޮ�!�9,�4|���A[y$%�����&'OEn�m(�����ۋ����֎��nd]���X�Dj�a���)��ro���d��

�;F�?L���
���:	�HP�e�{�����p�T2WG�am�ȍ�\��g��������Lp��V���	ר��5,j=Pw;>m^���u��}�?��h��:tp~��La+0�R��,�{>Gt���-&#�@�d�e�J@�,��c���! ��d�8�(�
!9�#n&0���}#�> [��긝o��������B��&V��j}ٽ=��o��V�N#��;̋Ubւl�'+���*!���4�N"�j�7��DՓj��N)=�vl���v�5r.�L�����=��I�@=���Bk\�h���"U�,BW���*c�\�q�֓cPq*Vؓ�~N�Q�nQ�BwRq����b�)��y������g/IP�W?��<�f/�*�5�;S[�,� O���Y�4y�"�^IG!�O�"�r
đcq8��xw�o�+�T-_�0q �-�f��no�O��^� 8[X�}��j[��Մ6�Z�E���5�S���K�Y�1$�����7pB��Ð�;j�ؑ�'9�/��Ee�ވ�IooM��)Lb'���ǐ-���%"@�����X�}�o}�!f��o�e�|�p�c���ж�*Gsb�������5�Y�T{a�o�X�\�_3K��w.��=4����%�6�� ���
F��fe��FT1l|l�VP��Ean�>��L�Ɣӕ<�*a.�-}G��2^R����;L���K����)@�nҮ�	���̳>��dk鏔z�V]H�NǻTEFoӰ��k�q�p��Ȳ���+g?pʲOk|�b�"���4�~����Ɩ��{~�w��ED����	��v��/d(�>����]܄ kaBF�o;R����ńi�1��i��Ge�5����=r(]6m�A>�<�G(�ƣ����
��ޣ+p�+�	 �;��'��3�O]uNmu�a�'/؝u8���H\>�}BP3F���{����ev�KF�WG�kzC��1v��=�ꞥ�=�c3 �n�v-{��QD�6�:������*j#%LֺZl�(�lݒ���f�ƈLH;#f�G�q?�?ILН���F�]�0'I
�Pca�=��T�\�lω�W���Q�������8������ �<�w3^��b��C ������e�*U�Q?�"�4Qթ�8�%0��S�חķ���D�*�����2���R��]�"�O����F�5S��J`�p���	���K$~>�Z �R\e��́b+B<BZ�EU|�ys
��-�B�m��$hy�/VO�N��3�Ƹ�s�	�
���mh�a`�P$�t{��>�#�̐^���Q�o}e�;����� �D��"#l�?�����_�a�8���ԅ��ć<ą8oTx�J��͘ ��X���v�ϴT-|w�\{���e�c>��iY)ದ�2k�Oiʢ��rFW���I7�����.�KRE������ì��W~��}W����a0Zy���+�.+����V�PdWqмfKQ�&w����R�Bf��!̕�)���m(�"cVY<
S�?23l���ߺ���<.�M�R�s�NW�]=��5 7 ��>�T>����aN�7'� ��K���ej�&CH�z�b�w5 ���iTJ��ٺ����,,U]VF-�ȂlJP�8���e��1�ʥPv+^}���km��GF#A�i�D�3�R!��y�d�.{�Ɛ�2����'�h�g�x�$^i�6�slH�%�֍G�*O~�Y`B�W�\�O�Dq������7��x�,����-#+͈�3�� ��
���u֥�d�u��M�|��벦ol,��.�N�ń��E|�ge�c�g�ZOB�&gE�f� ��n3ۙ�Ƃ����u���>� O6���0=����R�U���f��]һz�ق�%QS�#N2t��|�L�<��b1ػ�"E��_�L�+���ԣF���n��E"������	��)<�_�8��$ �""
�*��p��	(�TV!��u ���kZ�8RL�&Ϫ�5�Mf[��Ӄ�s�����<�t6�`�Y-��F�eu���N�✰=Hvk����}h .!�~�|TT$�'R�[鸼+���Ԉ���&Oi�C9kݺw��<�
���b�^Z�`�B0K����QD��+��>��}���z>O=����r���SV�R��Z��cj2l�ҙ�؃��Bf�%���=U�(������z\ S�����S��bY9��"}P?��g[/�G���m_�˃��]�O�-���`	�� ��m�S#pMrk0��j?�_p�,]} ���"��S�@�vN��o=�K���*�Ѫ,3 �P��Wp�'[�W/�Y�f�9^�d��{������5ނt��E�*z���w��/*�p�gh�!=�/+����\U��$�c�E�'�'2;��z*R��u�bT�%B�mG%�wX�Ж̴�r������9�A��2�ng��El��\jv9�>k���Z���H!2 ?�<�!�ޕ�l�L�������puV��l�pL��NM�O��h��F��%H�X�.��{#Z�{瞰`��l�t���qDA��U��~vV�2iV��sTA���?���/��^*�$��b� Gv���H�fb	aHEE��Zj�zu@.����MO�G�>dv��^�;$_���ǿ=|V��cݽ����Џ�Эj�z�0]^�9G��GN#��d���Nc��H�$�;��{V��dȈA�F��
zvX$Ii1�!��*�g��p-�!P#�|��>&�J�x�D��K��S�&Qu�<kUɣ��Z�C��2���H��+:�q��W����
~O�gg�W�����1X�?7�TJK<�&��BAI�y��i6�[�Z}��끺����7�3�����(��}an&]]�)����3��1�ddW֋d7���ÜsL�)o\%t�X���2�t�x'G�O��RP�
m�l�%�p�����&��Sj��g��Y_�}�T ;fem*�S�ʭ�ʹ�ÑH�U�����p��S��>O$;�GK�眞�M��e���c��仠,��f�6�D�r8�|�S�XZ6�j��M��(���F�i\.���J���X��e3%�c�F����K�����M~��P����I���W`�wi^�n��%�> ��X���3LI&Րgȴf�hT�dx�M���$���B�k���� l���G��9ܩX0p?�@B4C�º5(����#��#�*$97�+�����?���I��a�{�����j�`^*^Ij�*�l$�9��σ�'�^�>$��{�-����rTʤ��g���e+gv��E�[V3��hڮ�W+V>
�@��OcY*�8��-ϴ�kX�3<-߬�#�J9��.�T�Cn8`�%0U0,�.D�Kn߳) �UѼ�p;E*9a�&�l~�;�@�Y�����ٵ굈�n�l�q�'�W(0�[:����d� ��}СQJ	�fӿi\�W>����#�
k�����*�XY]�K.��<��>-/��Aصl������&��MY�� ��͒��Ȧ��~0|���؅�n�.Ѥ*^�=��~��}�c4��{���Hl�( ��?`j9}���Jb�#���,� ����Ջ�E�f�Ά$h��WB!�5��M{s?��t`f{����mF���t����+����L-R��x�h�T`�;�k�7N�6��R;�x�:3�_;���4���7i~,"���.��.���r�_/KE�b�2�*�w��C�<�K�%����e���A���r����="ǻb�W�Bp�U�T���'�14�k��Y_	��+41t��H8D����*_-[w��dƙEd}�d�o	ng�7�u�zRP+*�z'0�zU�8G���ϱD� h�PVQ�%�ĻwE�#^�PuG��֨�{*�����/��Q$���t͡���G\�*�MD�4��ݔ��h'�}m<$�
�J�h���-�J�[���F�$���w(sC��[����by�6i NK�+��d�0|A����|��s��g�M�33�m�j-���()�D�C!����-��S"��x��1����@Y�:$`x#p��]� #�D��?j��&M1�1`��)J-���TH��=N(Oc���J���)�h<�|�a��zIu�^:zߕ`�@f�]T���SN�
�S�����ǎ�-�Ҍ�_���i�'G���Gٓ�B�����G���	`tf��p1� l]Ұ3���G�����U����ܬ�E��9n{-'�w>�Fb�*Էʾ���SX�F�f4ˀ��f�z��>4�]HuD��h98���"�*8F��z��:n,�k�ؽ�$�����A��6�-5�j{*ќ�_��(������[Ÿ�c���2Q��Ѷ���[H0/�S��*R�vD�� ��g�*���^.ڒ��Q��P9�8�i��ݻW0f�֬<�>u��0|�;�nDI�XC�}����H�=���j��������|���tDKb���}zʨf�r��Y+h��z�\:XO���RsEk�M	Z`[�� k q�}q{WOs���Ĵg�*�ó�i4�J(x;��"<GN�/C�U��!f���Y/�w�!�<���^�'���יx��S9�"e]��듁T�Le��
ށ�d�>.\��>Dq?�'z�b�α��h���q�B�cqS�[�H�;my9�f I�wq��&�i����߇W�(�T���LD=	���+vÈp�°}$�G����9/�km��7��3&7�W���m���TCzH�x���b_jW�b��C%m�a[��,�k2_�� l"�R���<8X!����{��e���� =1�3#����n�K� �9��k˻��������E�ז<�-C���3��$n�����Z;����7%����%��1)@�S�"Yl���TY{��&@���1����\�H�ʗ��M�90A�>��{�|�	�'ʇ���R3(;��uu9k�i�DΑ_��-·�
�vm��1���#ut�c7���|x.-��e�e�t��S�S�fፍk�>1�Cu1U:�.�Ոʭ���uI�¨agVj��,ϓ���e�D��E/����_$5Og������I�B͐V�1�Y[��͜��}��\�΢��t�*U�	 b�BR�ܜ���@"Ch�����7W���g
Y�����U��t>g���(X䦔.�s��c��xw[�Et��J���`��|7��y��u(��,�(�����{�	M	Z4Q�����N�O�ץ\�U�G#�Y���=��j�-�J�g�Ԉ�#��ص�M]o�c��M�4'�������0?����b6w�C��u���vQxi�T
�4My2�a�ZY1,9��F��\��h�<\�-�h>���2g�����yÅ���(�X�x�O��9��Yw���c%���} ��l���@�c1��U�Of�P�vq��;�m {�!Ms8p�����Q����-uN���zVb��c_����yŚ�/[k�d���`��}�����?X�db̭�1dg��sM��B*��U�*��DHg���� �5?�,�rlyyG��W?���գE~��C8[�߸�>.�+�:��%��sUH����]�z�&61�ڟN'�9��j,���T=)�g��6Ymѵ./%�mS�S�95�Z���m����&�J��̾�3E�s^v�-�>�v����̚�v�Ȉ��c~�͛�m�{0@LHw:k	CW�ʌT6t�yL�~�d���H��z=g�v6ͺ+�y�[��Ei�h�6�Z�ϱ{t�Fޝ�	J�7�DAs�4��.��{/O��Lc������3�E�s�J��Op�F�R���.���<�h�6��@y,s�3��s�_�S-����bU �w:nAsʜ��~�E�&��Swb�:h.�����J���=�&���Q �ueT��X�IR�ג��a���!?,�9��j��.����<�K�	+;R�qmy���KZ�Nk���z!��tD�W�g��*�f� ��B�������vnЂ��a`N�kZF�噥?X-�R�oEu�\�Q�^5��J��)�b��q�]�i�]aY�~vuCҰ�C�Z;"I�^P�F#=2F���]����Ҥϸj�
��o*.�B3��J~?g�/��'��sOTIS5����
�7�o�ՠ�c�*M��W;�8��QY�ڋ\?I���w��3�%!`\t|�x���`�}�q��5�Ώr'mJ�� <XY��ֱ����Ŷ�mk?	�,�8��	��^�����	��|\7��wGhsؘ�GZt�5�,�e*�g��v,�Q�L�-�t����W�GJyػ&��]�pSY�wɼ�?���d��4��;�/-����6��V�>�B�2��='��L������VB���iR廬�~�t�A�ԑz����< [P��ꔩ�̺��U���oS,��}��އ�ƃ�����������ϱ1	q��zL{���Ns�����>ϕ��=�~���n=���>M��=�B�ァ;������E��cw��O3�D�<��F�$_o�O3� 
��kM�G�g�Q#�B/�h���?�CL�b�n�d ��w����"���3٥�r-��׎:t��	��l�Wd�Ao���\>\ӑ�&A��'��y�Oن��&��8��eჾkd�U���C�Y�Cjw�ٯ��?�y���C�HU��>�E��Y䵕�N���?�����WXdf���PF��\�5��h]����ޑL��Cܡn\�T#���e�ĸ��XUؤ�L�INң�5I��hք�t�Ɠ�j:��!U�K�=:v���|�u��ش�9���I~;��+0�Iv����A�R4~�ESUɟ˷<3��+ s&)8�м��s�MnҰ'D�5�U��O�����*,UHT��i ݾX`���I��`��k7x�k<E��i|5���^�O�H� yw��e?˸�������$��O�M���e�� }C*���S��tH�/�c#�7�в"r�8BY����]�����N��Ù�r(vz~&���ihg�}�HI��	�xEJ|�i������b����y����}��m�=^���d>�Qs��	<�x�H6X��� 
F�E��yt\���ל����/K
��ש�qi|�b�Z��z�V�#L���M���:.)d\��x$�)�8}�!N�r@xWB�ռ}�V{
YA>��8
6H� �9ڪ�e�����1F��M�hz�Q���mB�̢f2�l~R6|�A�O�\H&$� t�� X�x��_[3Q9�X"ރiڜ�N˓Sl�퀾֓�kB6�42Q�2���A�g��#��������5��x����F~��bp���9 ��_G$��5%O|������+e	: �t2�V�l]�����}~�j���澿�T�'�~/���H(p��Gj:�Ba��G���ox��M�pϭ�����PE*�m\.���4(2J3ƽ��������ˢ�L���UGTE�w��nC�V��3�Z{@^7�{�!<��b�����!f�aj�,(��a�Ğ�m��~�.]�EcSC�U��>�h	�Bd-�P��{����Q�=�I[erO�:"O���;��q��u̝���]2��i��&jX��|�Y冤0�FJڎ���F�������?Nn���=�CZf�C��1Y:_�+��`	S@4��Z�������"i.�)�������2 .��XaQk$@�G�E;��f�����D�a>�T��BRLYH�y��R�^���*��(ӓ�F��21u�����r��6b[8�DZ87��U.�Y�� �ipwq��ؖ7b�g~����?`��ę4(��Xۖ�)_�����t���P��dؖJ�mA�?�>r����o$������K�ן"g�q#�?d��v�ǧ/?7U�����eS?aB�rS�g䰤5Mw��N6@	��B�g�ޙ@�\q��K���t��	SI��Z'� �F�����s�.^hF2!4���4G�5�;��5�����j]�Q���0��Y��x�}9\��Z闻�Rb=5��>"9�C��zi���Ŝ+�n���X�e�L�^Ŗ�\�g�V��O��]��$�6���C@4��N/�h�a�M�1����6��T.K[��+�h�w4e`;e6B�R�����!�+�/XS��P|P�gX��)lK��
���B�z�[&�5���*�x��*]`�[�[�@] �t��4z#=��ە".������햂o��X�H���!Y��g8 !S�
E,�I ӂ��؂����k��y]�W�:^ߩ��]��9�·(����e���xc��Cq��FDP����i��J�V�bcU�:��m��Q9�C\ڧ^[�/����X@1B��jv������i)����!t�A:O����q����3��l]�=�?䴏�B��.q�ȉ��6�M�ʒJZ���v �F�8���'�=�˛�k1�:�R����Q9-��+���u�Ka���L��-EG�!l�2��91r��	j���QÂ���)��TJqe=<u����:i�."=�xQ��C)�����I����H��EUC��0s���-/��nv�	���R�0�G���\�H�<fYO����5�+�r�7so�	�qו`g��d��g�lRa��D�s��� �\" �C[�eu�R<d]Ӣ�U'�&)���XX�>�W��bf"�gɼXL��GΔ�J���'���������}ӌ�3N2D�E�X5?��5��*v�ڹ�(��$��	X6��;�O���~7b�Ct��8�(ڰE'^1�mB�`u��?��D��Ϭ7Zf�>`���j�==m�����D>�n��0k��������!������>���u��#��Q���i��Wa�yf��N��Ͽq��$0��$Z�����p�"֪)�M}q*��U�L�|��&�B�aJN#���vs;Gd; �;<M&�����t�S�!N!6�.� H�,0�M�m~W�e|�	�6�� �][Cn�]�?[�啼_/�X�7$h�@�[��Ư��\j56�tE����콊���e)�JL������2+�w���.���-?�@�o g�v�n�v:��4�k1���&oSOI���Sڍꇌj�dW�5
Fb�;b[QJ�NTO�;l����>A���%l�; ��2�ƚ���i��?Q`�:�]�8*�]\0�g�oU���@)b'��᥵��(CR�4Ej�3��#�us��J�Vp�<<o-i�IA��[^��_���l�H%C��g�l�E	���
L��A^!r�ZQ -�6�VY�Z�#E靈\��yŪ5H����n$�q�1(�d��
U{�}I��6e�7�D~IQ��y�"�z�כ
7�&�`W��h'���R��ZsϾ,q��m���Omr?e���(�ȳ_������o��AF6�;�3����l�K�j��uq�N�����2zӧH�DW�a;;��������6����8{x!���h���/~��ȳ(��Q����4��M�Z���2��q�j�/\;������a�Ҡe�!�8�5��x�P����vsS�X�C�y�K�J�(��jF�I�v|D�%��be��Փѱ-L��ci ��ܤujF0���,��=�7��*۝�"�-��qN��o�T6��01,��gKT3w�oɬj ���mhM�[�;�4]��]Zxg`{�a���.^�8R&��qKhc�'>@�bmhcI���Xj����c�V�}����I�|�%1}�!�7!\ܮP���_)�W'%�<�'��P�8;�h�#a�`4p�o��.�'���;{/���02�Ţi�I;l���4�.���k Q�<�@ڞu|�۳���r@��O.f�l����lo�ʽ�q�+�$�ʌ֖�|�.oC�ú�$�m�b��O�.>W;�v{xt=|�U+ò�N��՜�m�c�9dn������d6�G��BdM�y�(+ǐ�%�YR�1������H{�A��y�� /��� ���a2
s]O���D֔����U�����{��jp�����V�L��`֢�Y ��x���=<E��R):;�YP���uۄЎ�W�~Sx�H�eL.�&��.w��Ӵ"������S����0&y�p���|�����M^�d꥝b�ý�ZP�Z���n�p��]&ܵ��D�0q�^',��8�0֌V�L���r�'G!a)�k�֒Ԡ�U�����CsX�w.�m���9�m|��A���L,'�XBn��S=6����P�� ����j�R�*Q]�E���ѹVy�+"3c\�<͙���Pi��Ϝ*BZ8�`�(0���ɍ���`�����Ｊ��J0�-�^C&�сV��_2(Oi{�N���:aUo0(���Yt�\~D=#�������i#� C�Y��a	zϻz�Cl܉ ,]�1:� Y�!p��s�$�kt&՛*��	%5V���G��u#5��o?���=�aѣ�ͨT�}�.�j��J���H^��%�B��x( �٩u�W0�(K��	�w�y�͊Cs#sʒ��)���>�D��/i���Gx͎m�
C(�z�ze��Fr�����v���d�Kˌ�Z:Bf�$(`1��uE�%�����ꓺH�uU���q��Q�+�Q�|H��+�jEC;^� ]�u��ܥ���)ϝ*��1.\g$�V��G��E<��f�P�Q�k�/~k�IQ��2d�8�Q� �k���i�܈8(�EK��R�2���CNήjڴE���|��u|�^�L�Ҁ_�üI��|�8j���T�@�Bwp<��,��͹C�T��P�0�W�aޣTmm+�'G��D��gZ�.�jra	f�����ŸfNQHs^��x�U�`��	'��<�B�����r:�k�TQA\�����#�<���̹���05;�o������f�Y���l]=C�A%�@n�����e�a��O�ϳ�Ugm �*[�ߟ����U�$�Bz�TF��?���;�l��{�_�/4R�xV�մ��/��Uv�IQ�+_�W�s���^��tI��C�)��p0��o�J����݇��f��-�8�/H��D���؆w�Y!��u'ޖ\�b\(�_b��B[��� �M��ܐC`9#b�Ti�܍~���r�#׍�-ۻ��|S���|Ag��=w�S];}SQ�)O:��ZZac���S\B��ʋ�A���i���K��B�Yӳ�v�0���qU�v��aeCg��.���j��Wz@�xbd�\=f%����ranⱲG�K��/���?�9f$(�f7'�"%bIR��1������e��}LC8�-���p�O&��k�r�I��qN��iu��?�7����5n��3>����,�4�R� �2�c��'m�n������k��sep��3}'�͞}q�L�ā��MQ�NH鳪��
@}�i���x����@���-^C��9� ?�+CK
��iEN;V:��z��m$k_�#߄X�UC2�k��#���m�|��)�}գkf�9'�X�)�L��k��g��í����s�e���Ku�8���>n�U�ѯ�O��C e2\�yG������e@�o~�aB\<�	�HR�
�Ka	~��:���eX�b[�0�\x o~��/�!��!�pA���a"��g���S[8����ǵ�J��>8���z�&츹o�j[FP��1<�GE�>�t,3��ۊ����B�����FN(I��`q�����'���6A���y��~&�=G�hV���u��MUTq2�&5�ϗs'��7��e{���ɧ����4T�����Aw� �a��@��Ms}E�;��kmi�KUxSz9��`nʯ �R����Y�Q_���F� ��G�`q9���}��c�zw��X��MX�Sb'Fͭs����N�ǧ,�����-�h����u=&��	@y��L(KzX|�S�H��;��T���΂���O����M�`� �l�D����Yk}������r{�U���I��G� �x�]mT��Szg7i� ��kef~�M	����x�p$�]�fc����L��gk�s捫wǦN�v��PF_�T\i�����+����Ź�~q��.&'�l�|����Kp���#E��u���JYUJeC˞�>N��^~?�a�4ک����d_�g�?������Iڻ�^)V�B�A��i�r�W4ͽqmN�����E��&���Aa]����V����/��jәh�s�������pw�:�lE�5�b�N�f<���%Ϟ��4�=b
��r6�m׼s!~��}���P��oC"_w$$>U�n]b�R偘w{���|_{������Mю�:�{4g��1��
�AT�f�&����؜g��6;����%���NE�L��=M-��ʒ�/ӝF�{���+���j'XAV,zB"��ګh� A�g�����c��H0&�Kd�W����pJ��#�m���T���J�`�9H��^��~8?��H"�w+�t��~��	i������uIj�q�f X	 3-T{�!�-6����ӯ��lD���(��V�3�3����-{+=2)���nԭ�tP�gMR=���$�7��F�E9��z�eL/e��@<Ӑ
�ލ;�7��L�mЍ�r����P0s^��1��;`(������8:!��ϰ�{�B4S'�J}D�S-��B.�O��Z�f,B�p�w�[ {O��V'����d��ɥC±��,�|��Dr�))�ҶM��FX|7пj�/�%}�R/��i��T��2$�)//݅�T9@���w��o�Nv���D6�Mf0o 3F,};Hχ�(��0n�X�Ck}�f�I�RX�f3���D�G+)(�zzy��w��	�2���Fɶ\���+�<#�b���ö����JÏ  73���>�!��8�I���Z�h����<V�/U"Y�6���7�;��~q.� H��.�H������q�.�ж�#By%�2<I���B��݆:����=��%tE�Gt����CƵ %}ɀ�et����>����=�p��"�k�K>���zz��Q�Ԝ�z����d/�J��ա��:vG�j�m[�\V(BVX:I���e���e�Q�� �'|)��y��qb}����g�Y0�C�D3"?"L�eE�`&�90i�M���۟�Ϛ�1Ir|�y�Z��N��N=��\����}�tt��"�>|���'�̥�fj:ml�æ[�R���7X�Ц���8D�0�$������}��A���X�|T�ۥ�*�:��"��G��AXy ��>�nwIeD@тğ��"T'<]�qIȽ�
��.�^�R�s���[m��w}�k�����Lt{(YW�����1L+�P[A0���"�>�7�s3@��=EM�rԯ=��[��b�I*0���䓪�sI�Ŕ�;��^��b&E�g�Z�+�G#����?���?N�1!!���S<���2�@�g�O��`�ڗTXq�e9�dq�*6;V����k���GW���8�ꠘ�x����p�l�׌>E�,�6[�(/1_\�yY�(
���承W�I�~q\OARR�����@k<�����(J�Y��ܻ���?��,��x�!ޜ��
��K!,�s`�&�z�#(���\�"���@�#u��ZuΪܑ�����`]�Ϫ�E�g���G�f���RIe��~\��$ͺ�(p����p������1UF��	������������D�ᓷ1��G#ιݻ�ӲX�D� �G^a�}ZQCHÆ�(���!�6"��z8�2$�� �6��a3�Sܯ��:.0D��d��ȡ��bBY?��f�8����$S�D1n*f
/}��[�_�l��|d��=���5��4b��;\�;��4���DR���r@��<�{7�B���I^���|~F���������<�<���~��/DpD�ɜ�oD��J�q��~�[�#�v���?�f��6�E���5�l�a\�\\#�k��V]>��O�c��Z���͂��l�?2���`s����D�'/��Rm�vK0%�7 �q���B{WԪW�\�r̎n���}�#H�k�R\��E�p���amE^���i���)۴����=5�O`cO�W��@Wt�;\p��zw�G�NT�y�4W�e�JȮ�9QQ�f;1�?��:-�*�9;3�$43�Զ"#�,2�[�W)\��xM*��m�|�,�`v
���2V�����7�א�-�S"��x�[^�B�4	��9��n~���/`~�8�g1��WDJ���N��W�5��j�s6��٫JA�w`z��6�;PLw���<�s��)����]�Tzl�e���v=u����#�㛉�Q4�d)�M�����L�
y x{�;���5�͞H�E镟�K�vM(�4m��>?23um�ܼ��I�#b)SPUMCs���"A�ǟ\��8|�7��pwYH��y�li�ǍR_wP¸�7�\��pn�/�S�����ZI�������&������6����'�&]�x�PI�ì��Pŝ�)����ɩG��9�g\�;@ʈ��0��:�Z���G�?~�7i��]J�=b���=��%�����_}7q� ��~}8�H�wW�i0�1rV|Z͕�ąЏ����>fSk�m�l���\>�� 
	�;3���D�%
{p-���Ѧ���ۄ�o�C���O���㐂 9a���"�7��8z��P<���U�|b��y��P�̖� °��m��>0nzBb6�X�x?��cQn{C����'|N�`�c�����Uord	����rX�C���=��Ӵ�BɊ�l.~��$�7��D#��ҫ9����+����i�\΁!�~��m��dƤ�)��5�;�u�#�S�-_5�3�(�]cB��3�m�Wب+��:Q�"gYم�w���������Tg����j�D�]SMB��k�?$ފκ�d*�̘��!l�x|�������>(�?۶��Jn��t�=�o�o},��8,G�Ь�Ǉ�2��5�M�6F�FƭS�2�!U��S��lc�A�q���ᄱ`Qj��>
EK/M���j6)_��mOˑ��t-���v��V^���q=�w$˚�Y,٢�vJ�$C���TZ�H%�:�g���$�yo$?�`�x�U�M����[���ʄ���hX]Ϳ��@a\W��ŕ��Z5�|�a�C̀�ٴ�p���y9�ݔi���{@��.�	��%-H�\��|ɷV�ud���% &�>])�S��*��!M+�/6Ѐ=Β�;�B��J[�����F�鏠E8W�%��H��%:�|����� 7��ڐ�6�Ir�\��v�zf���ߗ����Y���ǥ�F+I�d1�F�/9i��A���ϩ��i02j@�@$N���(�0_ o�����K����	;9Ɨ�%��d9ue�Kx��ڥM���� �7��	p�#�������(�'�.z�}��S(�PCypCvU�P&p�h|ٳ�RHx�O*r��b?�(mUC͇B����r�$�)q������]��r9�p>���5a������t���$���� �u��#��U��s�ͤ�Gł���1d�M�����e�����Z�r���dT��&iiAn�M��E����e~�.7)����Q{l��e��r�1�,1y�������F����?�CZ����'�s�B�P�ҍe"�a{���bݐ{)��۹&a�����ˠ5I6��4�����3�P����i\�>�/�j蹠�[�a,)�Ĥ
�f��e݉��q�_v�f ��ɕ��2���)N=��=�'�o�_x��	��5G�>�W�����A���һ�kK�Lm�}��4��� �q.����s�X�zRy���f���Q��&r�K7n�|y�c.��H�Z����@}����Ę6)z�G�ܹ�}��	� �=Y���߶xd���T�e�Y/�J�������t���8G��;�����.A�̸7�` ,Ny|�]"�4��6MI�?���KT��E����%�h�0�'��Y���tI���
@D����Ș���'RA�i[�CX"y�Q�	+M(Y��(�^?g8�ۄȪ��*T^Ɓ���6��o~��|}{��{IlhF�x�j�ۮ�	%���p`���~
$�H�ߊ���R�o��x+�^����uD|��U�_���<� b�u^�	=�l}�r�4W�j�'8;,���V���D�r�C-pw�a|y�m�e��^J�"%}\���Z�
e��鞕�)����*��p#V1j����?�$���c��� �~���!8�e�x����q뫭���=Ŀle:&V�|�~f&W���ѱWa8�����혵4�����i�+Ŧ2.zZ�p!\��\�T�E�Y�i�d3%��z��[?J��~��O�Q�
}��g���	�|P�3���i�������vwGp�$qIص��_�-��۟��4i�߫^�
S$V���2��Y�
s9��=��N]RP���Hvњ�&��^!�[*4��i��K�/!���!�x}WGs����R�ᬑ��p��'�O�A�DǕ2�`[�{�*!���Ϫ���Le���o�Mn���d5
��q	ڬ���4Q�4|:Z�*�:h��C٪݃�s�O������pt��jV�`���/�����d�z���޴�J��MX�P�4]�գ�a����,��~5�x�<R���m\p��S� ���=.����GG�-s͋�D�ȇ��7��Lq:�)�#v�F����1�OJ��z@�y�`������;�/Qj�d��\���Ĭ��wH����8է{)w�%���"��JV��x[�-��˻1^z�u�q>�A	�G#S˭2gx�9�@�7�(ԇ��3�:
�����n&����x�f]߳pt�n�>C�@����2�P�8��,0���WZ�@���+\��T;F�Fug����ݰ�<�gm'���V.��?�T(ϡ��~!dv���/��=���/�| ����U>�HᾺdV�[��-s^��4i'��l#�y����dF	���19�-C^�5x�n��%�F�J�{=2!@�k��J������F�}�:&O%쳣��Vjp)��Q��fR�{���kqO�zR�y�mYv�+RΤ]�,���Xz�kbuj���$%{�m׃�D�O����N_�0�A�à�~�d#:߲�V�$H��	2��4n0J"���(L��z%�Q�J�A���Q?q^�(:�E�	��@L!����L�i��7�-��IMG|4�������(!�3��-�$��Rp=�>�ŢpH����Rnq��p�����N�F����.^~F/�C���iILx�� �'d�2���D���z��rV�_Kh<vO\)�/�����}�o?dw?��FU���(佅�"��wo�,x��}?�L� �B���h����;Z�sW!?jm�D�*��6wF,LFct����gN����Th׉�8�������	1�]�#2�1�5�̢��Ze����J�G�'1=7���Y�ʦok��9�R����IJ:�w�N���3����?��4���(TJb|���bM2F���Ol6s�3�1�� 1�ꅠ�O�1~��;���.�(Gvݛ{�y�4�
Ro,�rH��
�c���)���m���V����a�l-���{�Ǫ�B(Z>](�������%�E���Z�6K�T�<ĕ��~��%��Ԅ�1
�bkދ���~%,t���b��?�j ��bB�`G�.���XZ�KX�h�;VBDp�>쳆����`rxK\ʧz��沮�OHp�eb���\D��8D~���všoi�oq:R�ۅ2W��M5)��4d3���n?#���X�:r�E4A�A����{�]e��|�u
mKׅ?�v�$-�<��e���e�T719B Iz���o�r��Aҽ��Yא ��Fc��N���w�~���O$_��w��c���
-`�PQ��0��1M�[���fl��l{�1QTO�Bѷ�#j��R�h[���kD�7���ٰ�ś�[�;&�
�_�?B�(J��"�3*��5Urh?=iT�ҵ��@����}�	*�f�u�ab�r��$�����/h��j�����PD�\�ovR��iHL���k���'ޙ��uGl���k�2�_�H6iFe[!5(���u���R'h],�ou�&s�7��옐��E�$�;�l�K\3��u�s�v�T[� ; �(F��x���/,C�K��]fk���*>"��h,
��I;�]��� aV����9��}�ߚ%
��{�dQ�q^Uy~��RU��.�Sk᫷����C�\�5>�hoҠ`̥�B�|)m�Ͳ��߅�&	�6�Q���b���c��Ym�l����d��v���,O��C�5���>�����]�:���c#����(CE@o� y���]L�I`�S�(z	!�|����\��ʷ	�����a�L�ȴ���gǫ�8L*��e
uǽ4�=�c`�<�.>I�D�;��PL����VPJe��'�]ǘ�Y)�$Q�L�7+��m��K�U���ɿL��;;�c͈I�c<�$
-���l��E@(JEis�z���(�O���j�����R�
�Y��%�s��n$N|S��f��4�wJ̲����M�z��@m�.�x̣r��$//Go߫�cki�b�~j�޾A0��h�f$�@zV_4�����n��+��u{���� ��	�n�I�&��ߡ^@z��t�\emrj��o\WW�r`�Z��^2�Er���#�'�ԝ{��,���d�]9Ʀ��㒜�f��/ô�$^��N'�-ݾuZțQ�3~���]�a�G]b&A!J�
�^Y Č �B�ݖύ���0���p���
U���<P�=]O�}ۊ��G�E��~�w�E��V�5.WP5��� �� 4���ql7�C݀_�4��:D��q��7m`������
�'6�4h�A31��b2A��м���R�}]?�}b&�����c��DD�G�ᖮ��>�L\/��Cv�(NJ#~*�[��j쒻`n�F?�Y$L��{�&{����0�*��˦�W��Rd��]�Kr�0U+�;�����cyK<�Rb�F#o9R�ࣲM��\�4�	,+��Q��������BĻ�+S���`���sh|;D�bybnlW��Øċ�h�92�����*�� 8(����=K����}��ݢZ�UmR����|�]>��~{�L�Ӥӏ��_���R���`�-5��~I�8��F�B�`��U��/�:C$a�a��**
E�4��U��`�T���vp�;����V�~��ve#X��iv�>
��5z�㺣v�v(L��x��������f���������x�o����Ù�?�Ȧp�Ƕ����A��ͯ�l�W�L�Y�,�;��	�Ԏ][�-��YvJ0Օe*S��J���Ї0�'y�Xjq�֎����	�b+�H�j�ϝ��	x�&#,S�|fTp-xu�"���?i�ߐ���Yإ�{�iy�x{�2�Jwɳw�\�����w�n>g;��p��m�o�B����d"�ֈ�s�A�c龩N��m�R 	b��'K9���.R���I	Rj�=:����\�>N�	��l����T��L(Ja���΃�YF�mnYf�ꓒ%�Ь9b�����eP[L���a'RwX1��e8]Q�?,�S��*#��D֫M����^��{�����C�Fu�t�m|���~�.S��W�n~斅<S}��ҧ�=�����+��Wm���-TH���/j*����[�ѡ(}���5u
�y�[(�'SU���gŉt{2[�WjC�����)�K�C�N��M��3�J�_|[mc)�s�8��J�; �V���|������,<���KM�Jp�'@l��^�_�j�[�p�3���5J^U�!��l;+���� 1������"��BM;1q���r+��7Y�<S�N�v��V��)���xP\a�S�ǡ�N�kM�;36�2����6�t��V/�~wa�3Ͱ='����:�6 ��2��lY�^m��	�ښ����f����34�sV�.�����,E������\�ӡ�Erz�
?T$��?���mm�V�4L����t+��s����{�6v���d�ad��s���x��E�C����tsJ+�H
g��I^dZ�!�i3\��#����j�=���l;�1��̭��p-�N�s1���s]O�7=l1���咉�����C �+�*��3&)��/��%9�_w��qIU�ϵ
]���{J�A��v��k���k��g<P�倱����d��;1���+�	{�^ -՚�kLƛ7��� Ӱf�ca��"#�i�p����ĉt"q0�R`�7����S��Ǿ�W���=����{O�gl8Z�ךa�$�V��r6��+-�2��o��#��@TO��6زTgѿ��N���Ż�'U�Q���������0)�9[zpGE�D��e쥾��,д
�%)�4�3)���4n\��{�ј��H�@���+f���j���\��C�u��A��K>�D6Ɓ*�.�ޚ��1�$V7���r���qӞ�L���(8(���v!�{aUYo��Q�� �i��!���
��C�HlO�+�DQ�=7Z�Ov�������#,6wl��<��&�e�R�����%��Y�AJ!���Qޞ|�ܻ3�ar�#�+Z�W�u����j;o���OߌU1����L4q�S�RxJ�b?������Zv&��?[~'ݯy{��d�a��4���rD,Y=FaEE�%6�~0�VvC%�|�t�v|����a���{l+��$A�J�-�O�� ��f�v��,Yݻ��Tb������M��ձ���k�(��/r$fJ��o��6����a	5Tm�)�Q A�3��],�7���� �D�ei�2wq$_���8��Q՟%��oUFI��b���B�Z���!܃���}	aN_�?�(�$�D�gʡm�m��z�O@~.`��#zFZ [<�L��KgFb1��/��ʄ6T@�SGPĹ���|Gb2��$���^Frc���r�C�_�iC�JÏĸ7���	N el�aıԶS��{��T�M%��[-�ج����=B�W�Eob6b��h��_h:G�N���Ƿ4A�H5�����ͣVŜ���>��_,�e�O����Bb�;7��߾+|J??���N:�o�B�z���#���*�g<D"�L����a���Aٞaf�%��j�DN�)Wa#ݏ�%<�l�Г�Qĉ�0se����Q2A�b�������XF�j���q���ufu��	X-�S�oL���Fd[$�囼/E~�����vb�bLJ�/2^D݅=~yh!���g�!N�bNpq�k栠~m�c���0{����KsY�����;�����"=O�k�R��'�}�"�`��j3(�(,���GK���)R����
�O��:	��H��-7,�4���=����S"�CC�t*o5k�����8��=��uVe��F@�:�K���q3��E14��p��7���e��v�6�?���=�S�^�u-���ىx�H(�=k�A�|�A��fq����0����\p]�IiP��vec��5rE��5�M9� )Q�J���FE<M���׆�h� ������ ���Ͷy!q&wOs7�2Z�7	���t�z�{^��B��?u��m,J8��_�'�@����w�ުDH}@�i�L;�������a�=�_��$���9�[m=A���Ƃ�>� �8Ѻ�q8�X����4��� �)6u��م��T�6�X<�Y�����'_Tn[�f?��fn$�3��C��!W��;2�/��$h{lkЎ/Jz�:����g���;ef��u7K���f��+���� �~o�$�"h9G��Z�to�����=�<�]��nq��+	�����
Ds�.o���=7}���O�p{��C$�Q�:u�W.�x��O!az+J��G�0�JH᫮Ԕ@�̺�<��Р-���
~f�F�Q���'q��qPqb��5�^�X�Du=�vO������+�ɒ�~��*m����*S��X��=S��_Kh��}����r��y�1��"z\�����{�t��!ŎHD�j���զ�z�
���c8��/e:�����^��Mk�عA�2�5��(���Hp��[R<��O��Z��dt��sCW����)_+��:`�E����/�͇�$F�[��cӋ�cUgP��1��T�!j!�Q�lF�EW���];/B�Na�n�Y���G��bH.��4�N�K�hv�9V�(���_�Oo&ǹ�����kI���o"92(A8n�-�t�S�O{:s�X�iR�E챸�0[0Ky�W���p`���DZ�����U'-���2+�|3C�ϕ�vkm}��8W�(Q5�IOW�˷܅��|2J@��a	;w &q�
ּr��wm�/�,cqİ�л!��JP�җ�1$d�����20.|+��.�Ρؚz�F7Fˢ�ױ9K��dd�c�c�$�k2��7����F}s�c���*�'��5��78���Lq��>O�����]V�����ѨL��]o�S
���+��C�y�m�3��2�6ٍ?�-��#��Xט8���N!~��ap�%�_�*��Oj�����
�E�#��n����T��@�H:��26<-�t�G��2�-�-D�&�#6aK�q��o\�_���9L�WR%A��y��hBo%/��X
�F�Ea=�­>�|���A@t���)<�Gu�����='��Ȟ��TvYc��OH����P�3�Ը�u�J����E�"B��4���Jڈ�I�n�����/b�&�.Fx`;m���Y[!�>�(���X8����\� k���{��u�`�пH��5®=W�c��jXo-����`wf�X�@�����|@O�I��W:����*��t��];9+�َx@�h�"6 �e��\.�������;P�_�<��{ƣ��Rz&�������@H ��?�=$ȸ�O��d����H�z���jX|'��q���!��q���\�[S�==�P�����i��=C�0$yᶤ�F�QrV��lM�=��_�1�B���wC�:���࡫��Ӈ
X����EEPۼ��F�xZ�n>2����ԣ�(�b�Ar�=�����4��68֗���]�����p�:��\�*�w������w��K4�2�I�;h6���M�g$������°���Sk2�&��b���3���7�Z��i�֐��D�H�Cm:�U���G������ifg�@M��B��q
�J0� hn��Z}�7N���{�Wm��y�R�~�#��.R�m�]]���ZI�WA�-V�u��CHo7��� ��^���	�����8�Ok�޽���zD�.�\�x�L��@�LJ���yGS�8�	V%�EylP�D���kעj�h�6��RGM_Z�|=45k˄�1��D�4�qlȉhؽeJ�$���6ܻXD�n����k�-3e����Bگ	��{r�������e謹vVƄn|2y� ��&���*��K{�1��s���(��$Dt�gơm�u7Oz�旅Ji���x�Ա�:��ui��L��(�(��!�W�fH�@��&	�ZmF�| 4�ަf��>H�r���&���7ʂX6�`i����	�v����	�n�aUbt���*�
�"Z��:N���w=.�y��)��@p�U��%t��i�8Ϫ��>�F�.���*+m)]�Z9
)/��F�n���+|7��9��$<����$��h���Y�-�%�u�Y3$stu�R����Ӟ����.F���!��C����M��p-�eL�-ђ���-�*�ÎO;��v`R�I��1��I��0�c�ؾ�4j�Q2T|]���5�a�B����{ۻ"�H)��G�6�˞��d���">)Ć}j_7�	.�|6��A��6{���«�6����gŇ)T(~Ij���#�;��>�k� |����D���&'�a�]��=>����QXC�b6ޯ���������㹵a�%�
G%�Ȍ�<�s�TOC����O�����/t��N���>k��Z�U��ጨa���qYƦ��Z��0�m���P�
@��u��6Z�k�a�Uv�~�d<X�G�E�Q��gf�����B%�x��/�EL4��zFX�0p�6?p��>茾��Am��1�����jD����O�K2|M�Fа��8s#b���`w*�k����Z�ɂy3�Q�]�m�5Q�P!0@=�����$��M���V7��޶s���<*\�zC3L�����D<]�Fd��ոB�U>���S0C_�<����sI\W?� �c��TbsT7�.X��i^_o��&�UD��P"6F�џB��Ů�USִ�1�����T�_�.��fזA�'�������lڶz���1�:�Y݁�[1&��~��o�o���89�{R�0M�|�5��3���_�M;[3���`U*�U�R\k%��$�ٕ����������~��++�F�@�8��^&-��g�kI��V50y ��jGpx5��̓J��ͲC�D�0����b|���f��>��.l��VR[���ۈ�C�)�>�$����c =j��y+���]���������g��G��GY(��ϛw��Z�Cx���M�p�r鍮ɗ�R"��u�����B�É�~�<o����El�wOod�<՗v�}k��ٟ(1�mC������jS�^�]�:h���*X��_���}NsU$�c:��ʆ�t��S
�޵^��c�al���B"7K��XX�u�-.�/��xy��T���7f�?����Z7�^F����|�BD,%�bb�����ܚ��̚�� E�.۵ �4q�:�0PQc���y.���ϴ�x;E��}kv`wܭ�pR$���2^�4��N��ܬ.�-3u��5%|�a�:�Q�3��k��_��$./?�jbT���y���4^�q����bY��x
�����{_�l(�H�Q|*Uɏ�ԣb�c�5�КJ�JCb]�n_4�_b�͘�X�e	���j�N�#󨵊�<�����T�ʢ�ި��>�� S�co  <�Kr5�a�~�}��͔�9M���pG��X�'BJ����
�x�7�����I��!�Tic;��ME
���6��cSu�vSwS]�jL�\iH��m�NOA_j'29�B����=���:#PaK�|�(A�4[[�|�_4������9@�ݰ�*��+;��G{�^E$GI�k���~+1���QG_1��g+���U�?�H�ca���;�>���^W*�������f�d�⠰+n���Qz%^̰�J����3#�>����<e���8𔼌�O�	��wӉK��I	�H=��*��)qf�.�'�鳭l�0g36c�&۔�-\��F�Edc�|I�%��R�k�V�������%�5#bPEe'��b��p%�g����Za :�L�nF�t�9y��k��[��+�b�%��^z���
�N����xZ������kk)�=��s�V��"``�a1��ϋ�6�B�mN2N�<`��'?7��$����D�����G�o�u��/#x#0���B��x�D�0
1Z���위R���sH��vD��`ޫ���µ��?��.n ���^�����Si������ه�y�����-�g�g��?���-��}�h�ʦžT�_�0�!�&ꪕ�����~9�˨�~��5��nH<]�ٵ�
2����Y� i��j�4qs��x������F�}�!�'��L6����[�YlP��Rc'�m�ՖT��i��!a�\�77�G$�X�q%���,���;�����R��62y���W�DR-O�%
6��� 0�r�h�@$������d���;�ը׃��[L;��;����gBK����p���9w��r+1A>�6W� ��l.*X������3|]E�7xեHZR�BB�#̓t�ˤ��/�����BR�΀�Ͱ�T9��v{`�P�R�~=T������U{u��HW�t�dq��B��r�r��Ob��gM�LGc�#�����y��y��J�h'm B"���$��'�@îr3~�@K	Vz*�0����7�8�Z����p�aZ8��l�rþ�Q>=W�-j�1=��j�!��<�ɷ�C3��AԶM뵧��+'D��G6��Y�m0�%�`�;�H� ����E��.J��J���S��ᩆE+��hk���9����	e������Z!������Orkb�c3����M���n�\����ا�	���`��=H����ҥ����#�y� �7E�Q�mb:��f�t!��0;M�-b䖁	��}#4evA��C���!�;�G[c7Z�;��Y�HEc�ˊh�@�D����
��ӊP���9m|������֮n�1Q�f��o)��ŀ�pхr��u�UL���K�@�5�L��{���\j�Eҙ�t˲=�����\�z�x�\[6#���6�IdA��s"����*Gu����錱��C���"����[�|�/�%ᮝ�����l�q�?oV�&j/d��+ĴC�ؠ�>����`(Z�4��!���������F0�o/0 ����MӱЙ)C�Y�x�����ܫ����(WSN���[�]xivqa�K��/��Y�H̵�Ĝc�Ygϥ�g������t6�{˚��U]A���ě�ٲ�i���"h�V>uL�(��6FM'nP�1�HQr�ij2v^k]w�� ���y\��sN�M��ϼw,�l��V��ʷ�'�ݫ�Y&|V*�Os0��Xo�����d �)��e<�H��K��C���ݒ�k|�;�:c�;��[X����fV
X�ʥ6c��:~J���p��d ���f�+{s�y��Xع���
B��Y!\G��v�3��W��Ά=��x��4��#�K������Ux����fA8����x�F�h�ަq#.{�XF�1�'rN��6ˋ�~�;�i�F��J=��[��^�V5�|_d!�c�K���� �c�-��`i��&��ds
�g��G�F.� ������0����~���ĥm��hv��nÛh�7FZ�*�KU�Ŀ��/�j��͙wd˨�9��u��R&��U�@��.��/��/��hq<����(΅���glXz|����Ϳ���g���ţ��g�� ����rJmw����YV����>�]t��!c�dAΨ|Jk/6$��ݦi�>���-־��*IS^�����t��|�,!��Nh]�c�]�`S��sd�%����D�D��(�7s\�9aTi��S��}:���_i�?B��n��s.��.����lJޙ|��,!�o�7�����b���cf})ڒ1��	�%*HM6�z��ΐ-º��st��n4+��.��>�;^�=W`�AC��(���`؍���LԵ�ip�d]@�گ�`�F�I�x ��N�3��H<j �+V���S���a&���w�";��!�����J3�2I�N�`�HF.�D��6]DD��VVU�-m�π)�=�\��n����L|�|CbD��jw��쉝0nOPY�}ͯ�iY�c�ߒ����ޤ�S�т��Jdk��oyD�>�<��\ł�L�	����W����/�4T�����y[m��E���h��~<�	*�v����H�/65���5m�֕gT�)Q�'p�:�?�eƑl���4�q�,o]�g9)���X���yv���`��?%5���Oo��7�!�O�f ��Q���x�O�E.�]�\"����B>�vLW�V�|��ye����ʖ�oN���� d"�֦��1O����ા�+��R��d���vt��$*��">�L!��ϗ�7H�N��ОΝ����L�&��u�r��N�M^>�X1y J|�׷[%X����G�VJ뇂�����v���J;��f+����Z�Z�����&�S:��e�*�����~]�d��oـ�L#Iov&*ɀ�&����9��'&�=�H��V�������v�0]�F�@��7��G�8�q��%2v1��i�[�Q9N11�)�k3���ټ鄙=M���0�*�a�g tV�.���y�{�P7b�\ޅ;��;R�_'m8kƪ3X*�9�W7�o�2j�|�+Yǘ���*��q��͑_K��aw_�ALD{�GR6���1��U�
3���������Y�,��P��oE�n� h�v�ۈ����F�2����c;{�o"���H�F�Ȝ���,\nJ��'{����ES�X�����pݓ�t]��HW�#�2tn� 8���7�1n5&��A���2��0�-�y���c�	�}^�c�'���:��:�\k��Z�_l�>!��<6����bb�t����1�u$��R���z���?*���y ��F��B�������w%,�:�B�r��~א�<��Ĉ��Ӻys�7������\>����X/^w�Vw��5�5�Hb���oD�_e�n�Dv4�9��׊{WY0���r(�{�S)u4��g�^��#m�~5��� F��(��?X����k;�CB��G��q�����p%�N�WC5�--�����>�exp_0}�o�b+�h?'$;a ń� �1ZלQE���k��g����4u��y�eVwd�y������ݢ���4ӈ�+��)t���-,�Ő�:��T>1�E�g��Cl���|�FDD�0�#�(��!�S�r��h%?,0�/��UP����P��<�$T�r�/�U�j����y�Q���m�ǽ!�dc�s�,���M���G�SP����mFs�U3� �ﾻ�-O`��&}�a{W�гD��{��J� �I�m_,g��N[��ڙܵ���u8�/���m�����U��3{x|rCs������TQ�zЊ�N�>9y���N�������ú�>�)�b���V�c�*5�iD��˪��	_5�����A��*���9�Vϡ-P�*��� �Lm�X��k��/�@�U�� �:t��!�DIY�m�uRc�7rhL��Ŋ�1��L4����w�c����\�s��c���'GCs���A�1��0� +�<r0&̭�3 ������g���!�b��K�"w�HLj�k�������Qhˊƪ�
�)��M�Ԗq6�E����V;��H��@����/uxg��p����떹9St�1���A(]�>:f8Cʆ'��O�ۧ��^+N�g��ā��Z�ڀ��Zqە�-�IBI)@tk���[�Pc�,�4˨�B�Ή���H�cv�CĆ=�5�z]w�yL�^��8O�4>�����	��U�\-�8�����v��k�ƴVi?���&����)igG�tO�
s*���A�����	_�w�A��}H�D:6�9;�8s�~��e~/E�xq��t�f�z�ͩ���m�bM%>{'`w�� (u~s�Ws����x�b r''N��gS�����������g��~�iU����?i�5��ԃa����N�#�X�S���)ί<���Ä�Uޫ�$n��.����k̥�avX��A�~��2S��QQ�JL��8⵻��<�dv����͟,Wε�͊c�ǫu�Ce��("X��a�d'�nޔ&-�1�&���[׌��C�gF	m:>>������O��c�y�.L
�)|_b����%�Ϡe��0H�tS^HN0YM������<(ެrI3�j������D�B�FbJ�Iu�Uނ���jEo��&�����TT���B�7C<�N9 � �(�0�@�H����a�&'�
b<�M7�YbT�����\��i?��BB���A2w�����c=�E�.��T��0Hev��C�Q���)��J�z�Tzh:��u�(�������z��h����yj`Lb�|#$n3�d����F$�I��=�F�Cz0��;�t�-u�bc��d���s^�?2�k1�5�Օ#osx4������������k�N	cg@�%�,7۠͟�T|��ȟ���aF�Wu&I!s-U��\y5z`�!�V���Y���l:]AM�]��{��z{�?�����E��$کmD[�Q�����J��֮X�f��X۷IC֧yd�,��\���((�'�|�'.XdN��D����{9p���z�D��J'�'���vJCR��g�(��~jM�Z��Y:�\dl*�E ��o]�.e7G�F��B���D�o�7�:�-�4��l�y�?zp��'�/C��L������ȵq	ku%xZ��&�OОQ�ܼ�?��%`��<�_��lg��ͽ� �Cq��Q��M�t�	��۾�mo<BVEt#�$KW�.�i8 ���]aĚP!ޟx���g3�+��v�}�����?p�(���B�x� �y���6���������6嫺�v}h�s7̠�t�عC����noc^7@��֢8?.Y�l=�2q� ���1��ٖ�iڏ϶��@���,T��x�f&/J��]�Ԩ�n0�k�s`PQ��IG�@�ɬ8اC�I�k+�]����w�ܧ�Y!����jܔ�M�,���B�*U�Cb/;���o��=�Ŧ��g
D��<|��D�7�~ _^5��x�U�g^"���/��`�Q{ʖ����l�tɃ�:_�̖�1�����2��mb/9�f7��[$��Xcn]�Z��A��b��2�;����c��n����{,z�O�z<,�Ip`���g��1'P�֜;Q�@}�b�o�����	r�$k�%V�~�:�U	OE�1���bx>�Y������!E�
���T��n��E��~.^��U�c=�1�/�)u�t�Y��Q�j�3��ȋ'���Lr��3�t�n0�͹�􆨷ݔ�,�@��0��' �Q6��@D�ث$́�o���j�T����r�����8��M7��˒.�E����rH��ߦ��<6 -y�8D )b+���"��^9Y?�󓭵9l���� ,�5z4���4��<ao���9[[.�$��T����~�������4<�&i�#��ZlĿXmu.�+1�����?A��c�������A-���k!���1�6���Z�G�����l�vmUU(��H�7���<)�g�deKC5���&�rK�DG���F���R{�[��+Vp>hr@6Z8��OӗohIP��K��=���#2��S�R�� &���8���O>�'��T���r����H��鋁+P�a="�
	ȗ-�8�獎��3�|���r��{��:"	5�)���2R䇁�����X��鞳eqC���|�>;sX�"����#��-���>��C��aS�خ:�&,��]L+��;��'�ް�f�}��j�H3c���+�\�}ȵ�l�����p�z�x�J���~���Y[J
����}%�S��n������Aa#� �Y�a����#ά9��@�y������n�sw�0��k�8J09�L�v�DC� ��@�MA�A��ۊ'l�6nH���6w ��X��1�Ka	Ơ>���k�sd�}�@�p�C�\`�f�5tm�S�6hw��a�J6F/��xylmE�,���j�xh�xcb�	�fA�4��WuR��ܡs.��L���:=���Ҹ�����{V���2THsf�$۞�z�灟+��F�Ēdj�Ow7��Y��_bb���?������� �PH�kڣ�%��*Q �Xw3ƾI�crsa&q
a�S]�~ͶD,'l%ߋ�Q�NP���J|��(�"�$#Q�pf���3�zO���%#����(KM>�d �.�>��}yl�)���wz˃�Y8k�57�n�x�@�ya�@���Ј�[
g�n�(��Ah&~ѐ���O���g���FNꡖհ;��*�|��f�*��z�[��W�@�h7�Z���]ѡ�G~��1q���E$�j�~,J���}�i�1G!d��F��V�U�;	�Is�__��@yuel3ݰe��$r
"���%�/k�׌�O�-�F��ͧi���߰��$��q6fd�	փ��W�-K�抗�uD{��i@�ǌ�"��=�R��3�j�-��CM�ӿ1�����7ţ�x� ) � �D%
�7��U�F�«>�nA!�y�r�/F䙞���^�I8}����P��Rmؗ�X����P6��<����s)`��֫6u����>�2b�/ī�/���C杛FG�$�{皅mM\z$w`���p�ӄ �`�Z�v�a4lC����,��������b�(�zF,o��pN�JF=F��֡�q���iSǵ��v�$zF��I��ƳlF��ɶ�`�ڢ��<L�o�vK+�F�@��a�r
e�)x���vOh�)�"�� W�����Q)9?լ��Wh�U���D����AS?��Bd8#`KG
̶�<Oe�[d���-��ƌ�EP�r9��b�F�Q��>���s�q��N3���^��b� s��'�8�lf"��f"�5���4|'-��݁����^�A�VB��=�Uf�́ʷ�hJ�������M��,iTH��рk���'߅.�&��>xPi���ɍ9#�Ȍ�� �H�d6Si{����i���NF���7�,��tU��T"*�u4J�� �-x��-U�,B�	@�V�į�N� 0��h��1q7`UL�FJ".-!��h:�lz`��:6��}����xV�ٗ�a���҈
��N���O���1�pZL�2�cc�~����T�C����4�sׂ`���bߕb�P`�±����%�tJ2�]�� ��t�[��4h����_�20U���~�Lt���Э-1��]m�;=
���������JԪ����)�@j�����Pĉ!�+��d���	:��T���Z@�`	Y��A0�S���ɿ����' @k԰Rg��*��;Ei����|�|�s,��ji�7��_t �3��ܰ��
���g@$�����@�?0ͬ�?D{)��Y�S�
~/�N$]�6��T�'%>��M۷$�3�a	�����M�cW�D�Y(���o*�BKڔo[��~��ʄd<���$��5�^��k>�\���t!)�%J������d��n�2I6�%�lX�%���,&���\4���ZA!2�GzPrB�^\��ځ�q���/�8f� AT�������mo��&ޠ���Σ�\rJaB�-�W��N�eٞ�Ш�oGj��Re���N?��F����CD�������!�����\g����J��̪���IE9�OH1|1��^�>J�d8Z����㡷 ��6����y�9�i^�����^��i��;�b���u	b�x�l�>ɢ5�f����R��k�3��@���UC��C#sj�{���<�f@�
�_�?QF��^��V8Ծ�������Rn����/f�C;[�c���Lz�"	ex7y�bz����c�����A�R��0y��d%9E1�8���r�h��/s����^�l��������8�����8�W�˂�b"�ƛo�+a�����e �+"3H�:Oq����/���y'}�uS���R�J1�H�������,ޥ~��w�]Rw>����/�\�ߪ��K:�U�]��S�'h QO���& ��	��g&�kȪ�V��]FTEmZ��ɇ�,us�#���1�� �����g�����k+{w1�Y6��1a$yu�"�H���ʺ�ݮy���	f��6"���T(����rH���jh|��� n��ʯ������>~5 ����S��ހUd��Aֹ^���埣G�"め���N�%��3��V��t�y�l���#;�`�$��g
)�r5�:��ǀ�-����? �y��#�������啪V�@��S� �TG��Y�Ǔ�	�!H�V��r	��h���O��j�{��n�+��/�ug���I&2+
��y/�f���P����[���=��g{dj�h9���y[�;H`��9�^���\Q�H]�������nc����F��){����
���Kd��4��?�p�O;xGy��Tq3mk���a�V��?<�ϏL�-����I�c�I��M�bq �\"�
m�Z>�C�ăM4�d���c�Q�즵�lﬡ��ż���^W�#��<��JT{���8�WU�<��${��Q���ŭ)���������j�t�ϗ��'������3H�JHN�#k]X$,Yص��<N�φY����Kn�v����bQ!�k���x��/X�XYk�ژ�ߩi �멲#�I�]�;* �ф�l��s �gir�X�t/2��[U��^������V�/wg����by��wf�Գ�F��͇�USD�ɛoni�z��n��? �K�B"��Z��C��+sFf��mXd+�蠕D��ב���T��t@CtP�*U���|rKW��Ё %	����bOC�.<q��в�6a��+���k?֫���*'�Gr+q�8��V��)Pk+K�0o{ �#��7�W����Kb��mY���-J�7eހ��R4Z��a|��>f�$a�^&����k��y��֕T�sA�ϸ��� ����[����1H�
^g�
ip0��3r#3��*��d�
��_N��ja���e�fObe�[�L�1�����	7_���_Ƣ�P�C��L]���9�3�4ϑ0a!�|���#鄢(eu�AcO��������*���\��yջf��c�_ T�;���Ms@�{�«���7��]�����)ۘջ�鍤"TKU����r�����@�q^�f�K��&K�\�����<?1�2��,��M�d�(�*�ϩ��48�lއ/p5���B2�i�+��-	�N�7C,7vX�NR�W�Z��*���p��ѿRpy���7�ndP�.Ā�彧�ANDcBL!��:de�����s(UJR*�q�cv?QŁ�H/j��k5O*��׬O�I3��dL	��UQ��� ��;���$�F��[NՖ[B{���y#����0H��e�J�������t�ߊ��=�Þu����L
��rpj�Ћ܇!C���"�F�ȼ#��E��O�:��zl����X[ע�\ٔP-�Q�6�V'B������'�ᥔ�#�se�I~���	ͥ�#N�� �*֏��Jt���*0_w�|�fD��d�G�k�f�u(v�o�����g�L�Sdk���EN�"�}gxn�;��u����=��ǜT�-�p���S�ܢ��Ћ&��Q��	�����'��1��u��M%�����kx�p�)3�1y��+����`�]5��᫇����0LE���IA�U���8��n�FM�X?^8ޛ�[�U�n���d'�;�[�9�yf( �"4���
o;��[ώ�OS��2*�wXv���K0���A�E,�_�{��.܏�ue�s�wq&��&�} M�+����]��9Ʒ�J}����m8ը������$����
ן�̝l��r���^��g���|e�7�����)@gD B����ρV�Q2�{>2�B��bKM�4�tk/ۺ�G�^��m��^j״����I��DK}��L���nƾ�Du<�A$�ԃ��>�Q�(:xLeA�䣁$=��	���[�}H�M�W�0W�R���т����Ø%��aU.B#�ڴ^�6�̗��T��c�C�e��s4��3S|�ߜ1�@�HLmT�(��%�m�௿ݧ�q�͢�s�ۤ��I���6MOO�� 5��ϓ]wӂ<����f�E(k{FZ�D����n��;jzX~v�I� ��U�M����6�jL.�V˖y���;��_�.x��"��_f'Y�ڄX�a�";N	a������J�b�fٟ�p�*A���A�t/�ðY9�Q���W��$RO�zK2:�ƾk�J�!�A*�c�1����w�v��/�,����l��N����9���ʃ�Nou�۶�����y�^�Z7�幈g{%=c�؉S�� �g���¦���[S>X�QTpN6"X�MR����1�Q6�ڥ��P��L�G#���;�Q#�?����W��Mz@��M��>P~����0Ϋ۔1�#u��v���,p�n���Q�J���q���'jd�v��)a@Q>K����^�[x}�dG�����Ü�_�V�T�1�Y���O52o�6�JDIFb˪�&(1{�I ҋ���ځ�q_�I�u�vl��}h�m��1!C��&��/��+}h������]U8�ٰ��)��um=FJ�x��*�Yj3M�l�=֠]��r�D�!7F���g���SR�(m>;���>�h9'�J��G�+��>._�Ղ b+E_�\�b|���D�#�FU��H�V�&�AK x�~�w����L��7�QIB��z��s7�RĪ��d:��C��S���N����)�����)�X�+oVBӥ!�8��
x!sPGɒf���ɖ�X*��MJ��a��?3STrfw�S(%r:X�.O���$pkf8ҁCҤj��8`.'��p-3���j�ߏ�#5e����dH�ĝ��W�S�Ut��4<�'/s�-ě��.�����#`�4��� �G&����躂�aޗ5a����I�Ey�f�t�lu ˵���}������7b�d�J&DL�Z.�8h#��)V�}̒�|a�J�Y*��܏����2����>�6!)(�İ;ay�l}��s�S�Q:`]"86�|�����k����ۖ������Pg:1�f�
Q�i�����k�}�H�ۯ����XD��,׃2����7B
q�`�>�~YqWqOՋw�C0@Yz��[g��#��M�*���+s��GY����[�A���C{�9����}1 oyk2jn�A��3�`>V'�NLJ�����=�7�ek�gp/�Q�2�g $6����3�����}�1PC�q-r��$a���c���}Y��R�F[�o\@<�|���xI"ax��\�<����]A&�������y^�������Ysj�z�UաP�~��&�}	��+���GI���Pf�w롌�f(���n�Q9{�7��jz��mO8[W��2�M�e�2�V��H&���Af�"87�6� �P�U�0U�b���,h9�����j<p*6�7�h�W�1�t����yr)%|�$uӢ�p�2��|�B\�ʂ2�$�!��em�^}��q"^%c~�7�1�1���P)�x$A.��S��F�vӐ�#��P.UǸ	���C���`�p�I#�h��0c.�3\-�U���o>�\��M��lz�)ZE��g����;)��A�*�lg�xP�y$�3�ҤaL������qvnf��u�{ɗ���$B~�f|2|�D뼆KTz'��s��,����5���ʶ�+�~���%��a@/V��W)���=�!}�ajWUX�nr_\��������w���p
@io����ب��k@&������6��|O��@��&�4�5V�q��QG��g$6�?+;���{���'*T��5teӝxK�Y.�Cu�Yv4"�v_w@0��_����(c�)�x�/s�v���ӑ���Qq�]�m�V���4E�a�%=���?q�u�w���.y������{z�GF&���H��c��-�����4�hɱ�ZI�Q�e�`TA=x)ɼ_�"g'�	��Ԑ1�y����s��iv�c��1ϜO�O[q.Z�1X����2~�ʨ2���
R�3��!��:<X��f�������Y��,>v�+�i���8������ 	���i􎅙k�����6�����>�>�n�X��5��鱋�F�י4g�m��J��u��EH~��⹦r����+�$��v�,1Hfko}Q.�W��ܠ�icdよ�P�``k�4y����j�����s�ݦ"��P{�X�:�F��Ҷ{?����n���o��=���I�4�+i����ߖ79eV6[U�lZ���� ���ȳTct��M`�� �Ӭ����d�Z}�����U���ay�l��+��&�١��>G�&b�2��iO�/�sH��ơR���I��LBJ��b~�Lp�Om���x�,MJ��*�/#�i-�	�5�nbР���DQ��1([�'p� HU��h��`1�2�{�tp���Z@zd��cq�*AӉ��!"�a����Y�͡�W�����P�Įm�Y�s��bL)���i��t���e��=�CZ�0��5��v�y���"���S�}�� �c቟�#(E��
�mnM3��>g�W�t�{pEZ� �O�NU_�aZ��ˆ�D`,�"NA����X�C�|���.���Vi�)�
'crY�h�$�e�FLi��o�� y�y��-gƇ>�yc!,A��92�i�N'�(}X����?ѡ�z��!K��&{�b� ���>�G�k�ڊ"B��e�����%�P�5c:"����P�e>���=A�!e;��B)*�2�&�g���-��g�����<ml���R������`;Z3�)�C�v����7^�0?�`b�ᮡt�1۝�%�+rk�b��[�໗;���ֻd<ܻ[0;�}36�E��{j��^V�Ң�f���<f�
^A����L�MW݆����W��\\ ��F+�[���~݉�-1�N�H�p���X��R0�x���pn~�S���B���)	$�B�	�G�\D��	s��m�G��9<�'<]�GP��nt���h��9�:����'�d�7^�x�r�AW�XgZ҈]�:x���]�e�	�2�c��aUN/�Wľ�>!��@�:lK��:̢5\L]���a쁴nsE�k4�M;:��h0sT���B�h����d�=��Q���>Q��%���~��W���E���;l[z�/ҷF���;��O~����W{��������r���������#��SY��	�F���FȽ�]�h&Dd���O���wyd�u���-70e�[_�z����w�.��&�@� ��@�(��b��8��Kڗ�X^ӥy$6�`|�
�n=�m����Y�B$��l�/�<ydH<�Ԡ��,O\R��J�B̃ )���!��pu�I\���!���L�0�����P����D��B:le���|��ו[�>�*�Le���[8oO�x��p0�Q��[�~��rH� �pU΋�pO)S,�W�u�v"�\���C��qyi��Z�d;/@kc��w�Α��C�&����C��l������Sۋ��Y�� �Q�N{ɘ(̓CsPRN�+{i�ʅ�T�-M�X]kOHh����P���q%q�7-+�:�iY^�&0��e]V�t}���S;D
��Ҍ��0%�%���%`����i�1�[6�r_�,4i���e��17.v�?�7c�%d}�Y�
�����%��Wg����������m�4h��{�o��S�eq�6tc��k׷��# �M�� �>,"�a-��d�O~���������J�A���X�`KԉE6"�|�Âa���(�qBK�e��������zb�f3[2bMX�B �1A�*�4��`��5��r�~�MP3o��c	m�	|��6~oo����O5����ʂ�+\��������p]-��~�����"r�n,��8�7��_<>�[P��GE�k(4t�N��h�\����L!����)z��D��c�]���[%5i:wV֪˲�F+�\� 5"h� �=��Bn�D0���54�"������tJ�ʈ'���EX{�s�O�а���Q1�Uț��Q?Yu�sɁv�O�/�r�������AM}n����&���	y���-��R/|M�\ؽ=�7!���÷�i�Η�3y��}�X$���|NO�԰�(mr9*tR�R�+S ��ds _I������mL�$���2z��;EAք�y5ڍkc~��9�<��/����T�
)f>�7�gs�8�p�N] ����mF�ݼ`�S$�����Ćq�:����Qs2VF�C�Q{YS�Ty�f�rGP���G4�XR�K��v�#�X�ENOՠ������;x]3�R�w�f�u���}�����+����7�.��<vৃ�l�]�9�1�H����r]	V��4�kx������Bd��$�^O�����}"(�����.�L��f��g0>G�(�w�\_޳S_��/�CJ��|��S9c�[D��`wx^֠��l,w��4���dgkB��4�O�?z��l@�[���A{������(}����I�D�m5�O����:E,h��û�6t�p���K	���+<;�Xe���2b��Ô�y��W ������f!��[��}���Q��p͚#Qb&�l���0¾�8�P�K�B���H]&�" ��]VÆƫ��,��ly�U�)�|�>�P�����NVz���q��*�Y��b����n�����O~�f)��� ����6D�UV��:5�5/O�L����~��[\e9 ��B[�d��]�#�N��/�֏}�`����5�tbb�c~t�(P0h�;��L��q�H������d"��Lt,xlnbUu��"om�g_�����b�y�bۓ�P�3���~��me��es��ٝ�C
��&�'���=U��/�~��޵߈e�n��,w��y?) � H����ɔ�=�u�B`�+u�z'�-1uS1p�"O(,$��B�k�8��_BL`-КrN�	�ۀ����N��nnC!�m>WM��H��i���b5��n�_)(���u��(l��E�?DRJ�	���'ǯ�t��,�g��	����n�G�;3�u���	ۂm�w18��y�I"v"�C�T��l�f�ѯ��կ����9���"G��WUB% 7qW&�[O������qD�O���y�1�%�D=�,㬎/`f\�A�d���:Tg�%��
���k8pCruC�Y�n��;���ACϯV. ����sU��6���)~lWw��5i��#�K����.�x��V]׆yA�(����|�r����X��&hY�]�\]s�>�YY{źP��-W��J�v��W)���L��2�:zZ�ϧ%6��Q�As�h|�D��������E�X"C?31l��9��
�n�&q%�K
�Fߩ�3���ް<I���:�bĕ���ٕm'D[<a�jX�@1�}����y�s^��tu�٧t���M�er)K.;f�!�-��=砣�δ���]�|f}�M���d������F&6�"�$	�#�<�e`��"�����ȥ�0���Ќ��x���ȡcpq�akA�c.�QJO�|�+�=���2�qX5����S[������H�"��\*�΅���~I���3�Y����A7t&���I�a�_#�]��(���:W�b�T�R���ρ��۸��-�����-�kÖ�@o����^8ɐ��n!��cS��ܾ:�1�	��L� vY�wp��+��J:^��C<O����VB�'[�A>�Y�C�wj_���e�+r���ڋ���N�X�b�d����!7�2N2� �D!bq,:��K>$�:'>E�!�I�?((�8��Ӄ�c���k#I�o��0;[7�{�N�c�R�$U?���D�:Oq�)R�r`��#\�_ͯ��vq6��W���r�E�e%��p=K��|��=!t�9�狯��a���g�������x��BOizqS����Vᙹ�/O�h����T���k0r<¡n�a�aNs�}��E�&����Co��:\� ���I}˖���>H��~,m����~�^���;�X��p�0��E�uW�(k{�E���,�Z�8T��ފ�r�[� V8qq-8�~��J��L�+�$]
�l��v�鞤����IU����Й6>����WL�
`� vV���\�K��Hp��gֻL����Nm�a`"�ů"¡
'�X�A����U�(,��&�3y�q$x�aR�������si�һ]��{˺��*o��1E5
Z�� e������f��ԯ�eB��6P��og|�^�4�[5����K*�9驵���VHF�ns~�;C��/* �Z�h�r�������o�EKy�2)������)N�n��j��<>��6����X�*����|�Cr9��+�|Q��o��G��P����x�0jR`Wȵc�,w=�ɬ��>�[�'.2��o���q5y���J{U��dp��%n=-(���¿t��ܓ)�/Uȗ�,�M�T�>,��A���(�H��*���khL�is\C=�૫mJJ^�R�+uF`u��$u8��O(땙u�=|�W]��\e��Z? ��Txo����ʙΌ�=GЧ��^ �L7�v��?G�έܧ��4=f��FT�a;d>T����*��}M�D��7�j���u�*���V.��hp3��~s%��%	���ܘtU|��5H_�B���gS[�u��xҚg��C4����A:����6�9<�ه�-d�
����e�$1��ۛ�E��ֶ	�l��+{���^w����t;�A{�F���ߜ��b�3n��g��,���z3��W�c�2�$�Z�Bށ�@ܽ.��Y|�h��آ�J��Lժv����zy{����
	���� �n�A�p�*�����X�2�}���5l�ꝵH'`�rl�
��j�+���=��*�����*#�Fe�kS����yfN"�����.�ݝKk�D��d�؆a�p~��5H�yډ�<�`{�H��B~R������=�G�ٲ]F�p����}��F��_�ޓ��z`(�h
?�Y>#NҠ�N�On���Yf�O���tYM�h�=� t+j樧G���ͶH�u�3&3���C���8����t��`��+?�*P�
� �������O��W�����Ǭ�%��)Y�lAMvƍ�!dj��^�����5J�?�밒"�6%qg�0�r�E��r����C���/x�� ����g�z����j�^��W-'��r�� �g4���z��K�7�MQʋ3�$�X�������uD��.kC1tp�.���s����V�f�CŦVū��L�awa��ۮ{şk���b�*���	���x�A��.��`���t�1aw�Z�L�����v���D��HĂsk�_�Q��H�������˃����/��>� ����`�oub`━�+�P��V��������x6'�Mni����&ek��R��Bd���<S)��`���z��iԪ�LJok��i�+g���Eve������উ.�Swnge-�p)�߾��?��@ R@π�6�b�4[uC�9!z?������P�|kd��)n��|����!�N��v���@̘M"��l�%UD��1?�0���B~<��]z����f�zr�h�	M�ҩbg5�����%	���̴cvvS�5�}���b���T97Y��1[a]�YZ��x�K��5��	#j1(��[�Q����Nb�@��twm6�[s3`�􃃾��!���b�������k]��҆{��v�ֲf���8��,z_s���wz�?p�ȧ�O��{,���p �yR������p�����{��B�^��U���L�o�������}�^��0�X�o�@M#)��$�3���&GH����B������T�s@��791{>ަ�1���`c���m����Ƃ��Q�*y �W�[w��J�E�ܕєs�Kt;��0�96�oO#�L��`���c�s�I�{��%M�-�wfI��g{X/�n�8��2;�P(# +��ĹIN�G��4:`���&����c���d2�=tT�.��a"<����4c���:�1]�f����
�i�>�g�R��ǉO�������w�}�,�3/l�X�Ór9�=�V>��	<�ָ͎��+�[ȶ��/��{�*G�3��'��q�)ۗ���H�c�*0\�B���̶���m��T�;i	�]�һ�8mM�p��~�Qf��I���QGPbQ���Pi�7���YO��e}_�#7��[]ltKq��K���>�aN���4�^�\�Q�	`]��� �Y�S�-�H�X�3����|��"��q4��|�h���lY�[���MF[z�֞oo]/�����������%�z72w���F��@9fGfc7~��P7�R�}&5	�S���1��85�)z݃�S�0��B�"�Yc�_D��33%Et%Cv�FCL���=1����_�3�0^���τ�7�RR�k��|��~T�
�ח��V��[N��h��iN���2.f��Qc�#���M���ƥ Z#BP�2�kd�F
�Q�nB�P(ɖX��$��'�
��j	8��R���u�h;�$�n�oHlQC�:�u��m8�EG���@�Z�8��|ǹU���q��1��<�y������9�KA����S�&v�s�b3�vz$������s�l8��L�9sm�f�{3��20�����9:SS�ƛ:�т|e�W��-6�Q�=��L��[�I:G��7��Q0
f_��w$�U+�~�k46d����y��d�MmȆӊ��S�;/Ӛ*�Vz�w<�C�?�w�������x9
��_��6���D{�,��p_L�޺J8D�s��N�����)�L9���Ε`\^��}?��E�?�!�`��0LZ�q���6⋨ �Xt))����.��Wj�x&�y�A�!y���̌��a����C��ey+�����m���Q6�g4�P�o&�������!Bǆ_g�.��F�!�S������f%EۓN" ��y1����q�,<�a4?!�!1B��Ki"�1'�t~|(ƕEU��:�ox �No�,����xb���6��woR-s�AF�v#�2��uR�[��vŜ��A��R�m��~&����鼡�x�Y�����u���D�����]�}�����Ɔ�̌˺y�8=D]
+~]M�$�4�ck-rE�M�%ݻ��T���L�J�ewrKJ$$'u�`�,i�_Y�5*ن�SR�%L���Q=�����2j��]�Z�و�\u��Rc\��UvPf�~1���7��V�-�q��۩��ls�b %@š���,�/2`_
(�d1��_�����}�ui��U�����xcJ�X[{M�v��6�\8��Z����K� u���j���FWP�r������C�C>}��S,RKM�O�@�v$��Wΰ-��+���y�N�����
��r�tQ<C�,����*U#1�N
V�9#����ǻٔ�p^0�n\��94V.�mȳ,	�!������~�a�M�Z���+�x�J�a�}�1
������77����Y�0k�ϕzU��n��{��nV:�}��xbx�Z�iU
�;SA^�)غ�H"5�{0>������n�=��
u�G��-��"�oQ ��}��3i�����Z�һ�����Pżb!ӂ̤����+�?��o2q&�@ e���%���U�xGȿx�呜�&CL��饩�ݚW�;6!=5V�Y�K�~���X�X��
��.�)٦+�R=P�Dx��]��ĥ%��jI/���j[ұ���^Q��<.셸�x�A�*G�tW�D��K������e��V�4��J9�q��I���p����!��;C9���4!<ݕ���A�6�����K�;�@|�5zY�oc<�!*��!��WOm�cVn���2����I���T�7��b*Hx�5���ه5';Q7���ժ�#�&s$*��Z�O�2�E�}��Z����\:��T�8dz��`�Ll2��FN	����_�(����m�'zM5�5��!�^ϼ�R)��y��[}�eN�1K0\~'��n*��'eA�x����W1�����jω�*��+�0?��pު�A��Q�F�y�pM����r�/�d�3���p�a�b��y�����I�~��O�xs�u6��\�9	W�$q���9��Ac�M����,i��G=�:*IJ0�:�z֖���ҹJ���ZL��n$�UJ�3�}���u6t7�:%�׌�S�&"��3ۍ;���Jdw�}��}��|��f��?6����!1������\�{�X!�7n�n���X3-��^�)+�h��L�T�մ���6�ݢB��{�DWF��Y�RG�p�<Y��sO�C;u+�����n]���Dk�#A�k@��E�".}g]�j_�9��5��J Pţ:
|T��_���>�@Q��Y�ug��T�I�x��g�Oܱ�j<��M����u�"EU,Z���|q�?e��X��,�)�o?�s`�է��'E�uѩlnn��?;���3����sB��VS���Ӊ!$��iU��ׄΠ��Ǧ����u`��'"�Pd
��U������s�S���8l�n!��4�|-9�M'��wT�5��:0�Nj���"�gO	�J�J26)x��#�0�i,Qx�d��i
��y| �ߪ^�
��P܎�{��
�ّ�8.~���~�,��F�n,������N����Z�\��>O�,������M|1d�-t��?��jo���D���|��]�(Ӝ�/Z>�s6d�V�c��{g�<���`C��̔($��bU;`Q��v�ae�1FZ��c���~A1��Q!>8DǮ�;�{���\o�b�)��G����۵UxI�1�����~���a6��K܆����@���:^���vO�7������Z�If�~8�f9 [\�jծ�a�`�B-���<qh�����S�<�7��e���o���o����wo^iNԱ�U���Wެ1�D/TOz(���CgZ؍<����O�}Gv�g�����
��
�DjNY�ڗ�ьNJ ��׌�*��s~T�'r}m�ch �2t��p��>�q��S�������X�#�WJ��'��0��Tj���fx-<��\����6���j���M�í�Lx�;%�,�v	0`����'oA�o#��ADPP&ZN{6o)ޥ�OV��@�Mg	Η�o��/f(����N �G~�$�H����m��{�����)=��E3x���2(�.D��5��IŽ*�V���n��wZ��Ȉ�PK��ж����n�:���}���x�r��c�э�������Y�ڊ���s\�Oq{�N;��ZP�3�z�U�;���\�055����[�]�\�@��F.�ی!3�+<哒����0ȇ�2���t�3��^���Ձ�4��]�
�_JK_����9~��n���]��7P�1Q�jӨ��-��#<�jW^.�u͵�\�� V�5���"����z���@]hP�)�&�P����6�L��O��,�K�|A�K�'�ٳ�y�`sN1?pu�t��� nH�X��O@ @(J���xS��� �țt"E�X�� �>
���7���I+{�^��$��AҢ�Q�)P�|�壬�i��rD��r���Sxd�Ur����]�t��CĜr,j�Q��D��m���$�R��_UΔ+_]P�n������)&Շ�a��7U�a��J{;#wv|��ac�6�x4bX���r�9U��h�(���l��������G~'�%�����{�;O�Y¥�gQr�Uu|V-/�I�Q��Q��4|uUx@��S6Y3�9���`�����#��2SL� P�s��LҚ����^W��T���jE�Js%p��_;�&�U�Ap�2m^mS�R乥���~���N��^R|+�<�7���<3b�)fh=�ύ�A�?hK��H�w$6�Iy�p�Dg[�i������ٱ*�~�0��8�<�z��d
�����ƅҿ-��)^��ˍD�׆-$�	����UQ�r�A���q?���T��'g9;*��\�)�>�eiC�L��I{mx�ê�ܜ��Ќ`�X�wH�-����V@�GY5��&��?��A��0��1�ɟ��?ٮ:��[Iyk�C�x�"K��8hIxk.:�s��:ŕ��Cr	Њ"��.=�-9����<8z��	���$=�ښ���ŧ�u�}(�Ujf�ݭ%�}<s�l۫=�
�0��G�C��][UaoA߇|�N��lKfRͣh�!�A������OiƧc�y��t}$O1�TB12i_����I[^���5�����y�\3圊x��^�4T�_y;&�\K^f���wR�=�ʜ^h�//>"G�r���y@xy�-M=�jCRG��Q>Cr��Ҡ��v��@���ݴ�Ƚs�P���Ve�`o)�=��?���L2�iyZ�j^&�(3. M�5n�<G����.�����/�8R�F[�Z�˨u@���}�$TOo��Մ�s�GxZ�oU+O$�7��\u�
z����*�~� 5td��``�أ��/�Q���,�j���3���0�Z�淰j�H�n+�L�}o��Z������T�����e����s؄Ɵ#"�y�������������Tj���KZ�};y�2�6��]����������4�o�M��oz|P�o䋮u����u��}|�ʭ(���I��a; 1�Ŭu�hM�P������W�D������!w�f�h�p��F.e���X1 ��D�Yq�Ꮂ*���5�g�����6w:�[��2�I��7��O�VW�r����^oQ���@ݭ""�c����5��0����0���§�� 9�Bئ`�)�M��~�tA��˛���#b�&�l\l�J�H�0G.?s�]�o,~uJ�酎�ۜ�v_zB%�C�Sk�h���_$�Ƌ��ˌˑi�G$�\�V|;V���}Q�vtT' \X;�c�x�߫s,1�<H>]䍞��]�Ȭ1�Z�F�}�$
���bx�m�N����������z1o�.�D���^*
�"d�"Dδ�u4Zږ^TϹ$�תIc/Rqq�fJ�"��Ĳ���m�	U���d�Ky��)�=U���B_�� ��*9�����,�59U�g�~���_��H�4��8W㢆�G/c�"�DU����(z2��z����ɝ�ސ�	F����Å�_X��J�4���ӕi`?R���q�8C�C�5��Dm鮲+[�>u�s����g��1����EW-d��we���g䗹f��b�L.��p��	�4�{^�ȩ��	�s�>����I��-A>�lk���ݘ�k�0��P��T�8[,��D��L���"�c������N���5�#EU�tWk3�J�%j��I��86���A��߁@Q���pQ�]����Ya�٫�t\��N�^�v��/0�]Y�)��uH|sޖ��dpx�Qm�e�����ʲu�>Vq��S�!2����>F��̆�[��A'�Ǖ\�R�kaQZ�:4-����vP7����j�*��R;m��
��\�!�hB�>W�b�����آXky]B��}�&�m)s���)���S�l�ڤh��-DXc�圱�{zjG� '�>:�L���b�:X��#�L]��Z%��R��O\��E,F��%�~7j�Y��<��s�=cQw���q9(�?jkJ�@��XeO@��Z4�ɼA F�<j
�j54O˧#D�`9���s�U]'�aN��˂0�v[3Y1��R���P|���՘���6�@L�Y�s��>�Z�_�?5l�3'�8�]݋wW��;8G-K��t���^�X]�F}Ԏ=%t���ڠ��2�^�q��x��>�ߧ�j#�n����I��f)=%�X�}�?͛�/���ǒs�+��O��-�Qfc�Tk?=f!N����½�����\�i�`���m���J�`���|�f�C�4�;���C�1QC?6�-�&0�8���-��{��3=�PQ �ĕ�"t|�9u��f6��Y[���XH������ ˗GP�W��;w(ɍ�17#m���f.��r62��=׷g�c�T>�H�L��U�^]'�g��r�W�3A��frՁL��n��N�n��*��#	-�<��46RA���w~[���&��ؙ���`b�(	��g�)0K���o��)���u�y�OuTT��?W	1q��6u@j�<�j�
��M�f��:��ޫtI����-�ڕ���E��l�uk�3A#@Տ��+�#������-�E�))#?����{�i�X�цz�S9)}�*O���/��s���O��ضi��}�7�y�h��N���'��Im�y�\�|w�T�q;�r���b��ו�+�V�*�ӌ�b5C-eL%�H����P1�z�U���1?n:��f����Ҧ�Cwo��q$���z��QO-Y�5��O_
̒��2A�*�M�Xs���X��Q��ƥ9y��u܅������"g_"Kn)}g��~(s��bv\�jh�~Q)h@������C�^6��S�����2f�v�t��c�l�Db世D�@#D�����
w���P�q����ͥ��)ݟɐ)I�ET�����ɒ���� �>Dj!' [L#>�X�ʱ���L��d�����(�\O��������_�Zꗫ�#o���\���s�n��wN.��n��[`$M��	��"Sr�2�	�D��Q ʏRc�I�d,8����L$��P���!|Nֶ��*�"�l���p���l<��OI1=�:Cs�K�(r^6�;j**g,H�UoOA���$���[�w�"f+��L� ݌T���*e{��eu��E�$���|ɾz9	=n����5�AB�u�xQxE���G�hx�_�ӧ�Pݎ]R���a��.���*���v�̐�'�M;D�`ٷ���	'��xsB����CM<])�:�_�Г3K\��4�v�Up��N���������(95G�d�V���q���Bɩƅ�֠N���+\\�m\ ^QŢ��3,Y��f��)�6I�243d�A����8%��_��	(Tg����I��3���� �ˊXކ(�A%@j6�
��V1�-aׇ���!�Jn�S�s��^8x�>Z�p5�?8E����'�������L����Y�>�SE��������$����0U�|�~^�:*¨�� )QD����'���0�y�W�2�$��l�
��P��SF��'p(Uu�"����wC�6�;�Ctg�>^��&��d��ڤ�V���g��o{|���N��i�!�\�&��=��v�g	҂慠W�ͣ�+�� �ۙ�<j��,�v?��ۤ����oW{7ҽ���A�����ܽ^y� @��N4L�$�LF�{Bh�u4�]���*i��d�ʞ9E�;`v���ʧI�:�ǩDjd�<��R���%�HP��Nvk�90�0���
/p�՜�<��r�}#�]���d�V v)H�7Qi��O�%�cXӅ(W�V-� y�DX-�]~��/�O�� ��J)H$u� H���a������^c)�������ଯ�pD��WA��C�P�m��æo��oa6G�/���Z��zo^kq
�`�:!Ib;̻�w�f��1U컮�z�%w��Տ	�A؋=�Ou5�+*��������u�ۤ�>$�|J��7Q3��tf��;�mWݿn�����{|2aa��B���K�eXN����y�W�Z��f�ƥe�HI�Bhߚ�,?�U�����T���� h��p�`PO��f�<����Rj�;I*�5/:kz�As*��u堵FK{b20HoF�����ᑮ~Ձ��y�����b
F:u���������V�++�z�����K������9(���*#��	�ԑ󠔪�)�P-	m�,�������}i�c������5���f�m� ��RE��읨��+U��q�&tKf�*N���]3�Y٧1�-���v#��%V����lD�5@a�y�yN�ӿ�O��#���@.befXϔG��>���n��7�֩ś�"\�L��3&L x'�p0;Q[m�ӓ�«+Tj]P������Q�^r����w��K,J�U�{�KK�M�������� �հ�ɅD��3��b@���6�_b$�#�
'� ��`���b�"�����(t�4�ͥ��`h��Rp�H�W^=r��d^�숵�����/�/V_���O�:��YoL��˪~-Ӛ��q���i���1�>��h�,°��jn4�Qp�E�G�6һ3���`To��+.ej�j�{����9��^c�F����{[ˆ�e�:�9���*e \,9
j�eܥ�Ӛ8Y�=�	�B���'�Y���JߴĹ� ^𯸂��0����q�_6#P�K�flu��u2_w�kP��Ѝs��:���1Re��W�堡�E	��,5f	�5��0֨7�z�e0|n�\�S#�aU!G��v�np����]�uqn���_mW���� ��U~��m��jҧn���!�ǂ�����������m,S���Rݭ��0�,�����4S��q4� 9b��+��jнHT�1���R�~��2��3h<�w�g�2�$媝Ƒ����y3{i,�|�ة"�6��&����a+	Z�'��|�#R�< v�X֭d��rb�XX=T\54�����о�����l`����d�W0��Kp�|x���ȍ�����`�T�;6
	Ҁ�)Mm�p������5�Ě�BY�J�����Gc���8Ї��w�.e�AKh�7�s���;Iy��=cl��L��ǕC������
�p󜫅=��I���D�ɍQ��>9T)~ �|�{�3ZJ�=ϰ���WW���f>�蝢��G��x&��R�R�0=!�)[�c��V&�)�#WVu���_����84�܉^��ϣ�=�w��X���zw�-�s��d��G��w�.����_��ʪ��e�MGљ�%�b:a?���J��(zL�
�ۇ��9��X�M�H8����g�9���
kG��	�5��j+���@�a��jlC	Z�x��BNޟ1��W��@���	��`����L݈T�T"m_3����Q�YEy������r�a1g3?��WhV9u[Ġ[ �kpcm[g=[�m�d_��do`��rI�Q���l�8�xn�D&*vt�'�1yG��l��{�M�%2L���7�.�c�K` �Ig�Xg��=h��c�*LFw#�1���ڶp ��Q8��^0t5$S����fP�!��ͶH�G�̯�8 ����\i&��9���֠��M�E	���6��hY��%�!R�uE�/����qd�� r�.fe)��MZ�SCCI����)R<)}����n����|;���Q�;�AnH��$����C�Gw~F��Zu����8T���ib�8`y�����p��m�ш�2(�%���E�C�t(Cc���� �B��z?G��S�p����.�R�y*��!�������O3�ed�}�p�cF�?B���{o� z���n�׃�:Ŝw�O�L���P��giJA.k�"��y$�©�&0mi'��\=�'����T.�emio0��V��!�]���b��a��*cOa�j�`�ű���t��0��]7bE��<r;QГ�"�����4��<�0�hA��� /�jG-r?����Ķ?��=�`�a��-n�(}�l2D�U��X�ҩH8�/��'�ao������`�d� j� :�'p��e��$��x��:U:�#�� ���j����PRC)P��RX�p��)��m�T�O�H6P:�%�]�T=g���InhT	R^f��Od�o-6� 
bZP��%�u'Qx��p{�Z�vk3�v���v6���i;ǘ��%-�������HR@�#�~GC�A��t�,��4].�B�.��y�*-��~�;$�C��V�P��{�/Xg�w3�[���<��1��9����@��j�m����ꚢ��@%���7�@ g���h��M�f��L�93�-�4fb�3h��o�ː��t�����#}�:�1�q0FS�9r������CJY��׆�;"XT�n$Y�埾<��"��St��=S�����IG�J��w��W�l�2�1�"��;�k��Zߓb���R�K7%�8*��ܢ6����9Ybh|�*�r�:���"���9�{��s���>�C����$`�(�֩8���m���V�����ajE'��ߘ熪HQNIm&zsO�	���s�Y�|߆SFu��aS�,1�N�?� ��"�dc��|�}��J�`���b`PZ.�j���6ݠ�t<�ǒ�-������Q�>@_Z�2��Q`ä۪���QFp��������:�6��\ź9�V�]�gN�`q6$��;�6y��|�	5d޻b;���r3���z���k^�W3L�T�fJ�ԅ�1l73��8�;;�I5Ȅ���!��V%}��ς_H��ݺ-��M�7��v�E��Q�-�-�,z������R�ǧ[ũ�����(�?'9�D�\v!O�{�������(v�~Β��%�A���6�9
��(��o���K2&��gf&ߜ�5 aI���f ��gЋJ���M�5����|}�VEA�6�:�=c�h�k8/rh��Cօ��6�Y#,vP�'�/�l���	fV�KYP]�,/'8�7�k.�>�ݑ(�K��|�l�>?�z�w�1�C�d��>\��qa�Q���g�A��p����P�c!���;Ŕ,�\�y�4+Kl��M�@�����zQ���,ʎt��|ѵc���T�ʿ}�� �pU���w�ܨ������Kz��u�_g������K��HKL���Yg+�G~�颇/1���jA%R.�l7���|��'W	gJ���7��ׯ�'�+ ��
w�^�l�I���'J⼺�i}�;�9�vx�<$K%���}�`ï�j������<��h��#��B��LQ9��ʙ����b ��)WUV-���e�r3����iJTI��m�OX� �'��y��dWbR	?����OY��w"m<�/��T��s��c��������7�]����:G�f"���K���E@;�kyf1�\�~;i��IP�S�5$(��1�ho��#�
�Y<��ş��J��� T���C�։�0��?���B���4<.[ -�W	�B� 7�+��ȗo��+�bs�j��7��+����	��%|}/�/��,�F(� ��JCM�0��q��������𝌊<�Ēi�����8�폣�t�/
�=�c"ݽVu�a��w�٨1������T����8^|����J0!g��� ŦW�Q�����L*��m/V����l��� �p&����%�3ļ������6mF?�錦b/���K��k�J9��~2��4Wx��W���M4?�>\��,T=�;���4���1$�Za��&�������oWj<������{ߐ�����l��Ls<ĵ���#5�h[J��a;d:��B���~+5C�M�J;�y'a�eb�{�%ug�`#Nw�-���`��$�n.��[LU�/w<�٪��ˤ6STg�;�-_ȭ�F���VX�:�r�h�"~���ђ>���[T8�����Ҵ�<f4�@[����uFJ��z���]�D�5��J�
O�z�'b8k��̲�ӎ\n�V��;���ei0��+���r��u�2��!��8+.�ݯ�t��  ���xh|�ٕ���G�Axڍ�Z���:�wG<P�������/�$S� �HK�Օ��	lW½��hBe6�;�9:�������^_жt2���{�A~�p�'�,r��{DId\�#���gy�9acS�˥�4F�����Ql[�����|E��#��a�p@��W�
<r��a�Wr�-�R`�8X�O��5r7g�Q�K�8�QEG���@u�����}U��dd��I����*2��EN3�	�lP��QKe*>+Z���W��r����'���;�����5~'�y;��6��L�$~n���U��p��BSd�j|#���XM4Z��*bʿ�[=���bXY7)�!]��ǇCtց�[�j�Ի�!6��K3.�s
�U�G���l鯜�=���u�}۬�M��\��6(�� �8S�6Л��O�9�8�BH5!���������\�P�G��9����g�hVem!��� iA��~.A�B�U���r��p��~MӸ:��2���8�\U�hX����	v�!#ji��&��q��T��m�ե)9~�����u��Ue=�%v{x I>*�ʱP��7���C��(\�F��q���08vr�&������������Κ��j�����	c�;�ڣ�p����
��������ط%�'~��[�gi�2���y
�nfh	�t)u�M�5�6�v�t3T�qN޼	�IbI˖�Y,[l>�暈<�M��`�m�ۓ�2S$L�o�;=;�!)CK�^�������b��ix�ܨ�z��;*SCs�A�E������m��tಝ��NBf�{�}�3䒹��U���&�����̃�e�B:�����{v��̓�E1sb��$h��6�n�!�)~�]L�}w.����/v�j|oO^S\��*"�{��L@~���f�хlTb�s7<�6�T`���y֟�������#[&nDnɮh�����s�ǌۘ��wR��!��y4��'$ӣ�؀Y��:u������ű�ŝKo*v��t�+y��ٮ"�,�WOg�@��n�UM�Gu��T��1-�ՠ��7�rb[Y(��Es�`�!Sͷ5�)�87`����� �ҹLE��7�kv�������?�pL���q"�y�ȇ��j�>�Fi�-�^�+���q(�_[���`�LX�^$�P��׷!{u�'�9m���qO�'5ɴs#�nm�YŸNx����p:2�jz� L#��W>7q��^F;Z��{�(U�3�j��6��s~���x^~@RP��-���pE�`���Z4�D�F��ϫx;��ܤU�f�Y��x'��y�����,��8L�:�dl��	[He�<H
���ʷ?��b��к�{9^ۂ�Z:Ea홒g;G�tp%}�.cw.Zv!]�0p�?0�*"�Ѵ+^;���):�� s��<l���:7����!u/GZG�\Cv��«@K��$�5���Q�p4��u&�/�=�1���t�\���x���	��3a
E�ź���.Z@^Ը��:5���k���l��0�O��В��Z66P$d�-��Z���)T<�r��o@���|�Ɉ����@�rDG�� )17=K�C�{���e��ZZ6�j�:�{�_j�g5�������{N_M7��WxЩa�0���aх��?!1H�M|�-2���/���?K<�1-� w��o`C0)�O>�)T
14%x�U�҈���6��M/�ܭ��P	��P�/���+��E��~4s햵�W�z@O�$Z$?�3��j�X�|P�RR}�e�JA�I���$�����g�V�fT�����f���'16i3�7l���>��6�ʤ�	$�A%�܄p�Z�`<ä�'T������%��N8��κ��� �%��X�y��шޤ�=z�I�jEA�_r'Rp+&r�>����Qɂd�bL�mg�J�yݭQ��<��� �t�ڙ��XU�I����v�����R�m����Íj`��?(��CL&tg|z��v�rmN�&��_�3�8K�vI�f^�$$���\�����j5!� ��iHyD.�P7���2��G��4ݹW��!E���R���2ê3v�&#ђ')��M����G�����sw�Mv��C��ڊX�a���J�s#��ɔ��]�v��A��roE���F	#��Ze�a>D����,�J����=\�(�ͥ��k��~&��_����,��ڍe��"Y2��[���dx����!�<��cq�%�d�
Պ�g\�3��)�R���Ж�fU/#o��3�L��+���GhķV�.zL2J�<��m���)��/"���L߄�2��uj����g/�K��x)����S�w%�:l��_X�0�|9o��{(�Tx	�S_o�\��s(����$��PvW��F��e!�7�{7�q*"�����"�����@��M���0�j���,�){����x���ٰ^�+�|��H�g��m���ڬ���Y�MQ�'�B����!���|��H*&73����aTg����>ٺRF��vAX1�}\f��taS�h�w�h���X�Y�vq��Yx�-�'��m���m���#���x����;�2���OC�!�\<��������]���y�+Iϥr��0�r�������6�:F�|p{�i���l^j��&����[V�w�uj)��r�nb1��/��W�q]	d(�d�1�C�$ϴ!E4<��(�p�"k)�(�(��m�.�3�J�a0�iz͆�A�'�^��T�C���>-�Q�r�Hk�;��ؿR6�Pt̹w
\_2CH�����S��!0�}!�����lܾ��[9�D?����^�f5E'��=ޒcDM�;�x��A����Z�xsr�=5Ҽ:�]i��EN\5��?P��`�7\R��h�u��1��������a��JM�L��>~o�8�A Pz���L8�=L)�`�H��ja����V=S����M�L���mv�=��H%|����}W�ye}����ؑ�rG�"�@�V�ݼ�����kR��s[�Ns��1�
d���I��W��O�JJ`�X�^�-c*����TN& �#��y���������5���?��<BOF�bCG5GV�}I���W��<�+��LY2`��$�0���FqTZ��w���Ct%��I���KraW�(��r�8V[�-��{G�k��9a�o���@��]�I���A��W��>�� �OOW�F��>e&f��p�C Nơ����YOzAF�(�gL�g�B��B����_��bܗ��܌�ǎs|�T=��IL˾��
y���=�Ѳ�%�m�
c��d��Mf�ѭ|FB7��*}����'|����@�&�l��(��/V�,d*�R?��Eѳ��N���z��]DНW�̢U19���{I��;�[�M#G+yK^������K�(D��3V�,j�UX_�*�О��f��f=sl���W�ށ�6�+ʅ~�T_d���s����HػE�j4S��mW���:jL��(+�Z֔-X,��l��rg�!�)��3Zp�'GHN^۷��8�,���w�B�\l�DO(F�3\��>?,��ַ%� �=H�����@��eR�}cbH�Ո��DHB��9`	�,�o��F�F���ʡ�#k�v̞��fj3�[���"Z"G�;�dt���e����ʙ~q�~��qV��x�H��2o����H�z->A�C5煯�	i~�|I���L�T�d�]����Xm��£� ,W��� ���E՟/���:�6��������n�ý4��/Vx�og�&����N���;1���z�/D]1=�a]M#?�t���ȢQ��}j�7��m����`,�9L7��:��)�&�Y��^�M��%�K�,}��X95^H����\\i3C�>u�?-�e}�|;AN'�-�� �1�Rh'���z�w�E�q�U��p�s�Xtܶ���I|<50��[�9��c荙i=C���#��U3�Vڜ��?K��(����a��O��;��yl���Ơ��:�X�x"N�u�P{sl�q0g���o��$�Ƿ{���M�W�qK̪<��V^����HU+u`�Zs,��>�s���P/W�mB��8f��/�24K��D�L����@�FHZ�,R�c��d/�
� c^�6
/���t�mk��)#�}��m���ư�C4u��
LJx�����P#�m�!Ϩ�`�[�;�	�T�0���7K���K��q2��>9g��K����.oU*Z_'����Mqe53�e��[�@{��y�l/�y�n���&K�G�ˊ&\�W�-J��\�W��k0�	���V[.���azH��+�s��O;7e�(`��Wen��%`_�QL�avX�MWj@7����^�Q����+7��:ǭ�����Ff��l	3B�A/c����������p�(O�v&���S������ϛ���E�4{�`���!4����x�Kr��L��Z����M����V��p��hR|k��W���UWJ)�#b{��&kC5L=�D�h}�,VY�@��Bo����)��b���{$۷�R�)�S_4g���a�0B�9%�>�G��e���L�l%������5 ���(>v�Z���s�j�1����C�o�}�8�Ⱥ�u���d#O�b��O��p2Y��T��eP�9m��4IV��)Y�Vhj��DS�[��ʺ�Fl��6U�Q/M��J�4u�"���ڰvCL�j�g����3�is��o�X^��#xs���
�_*dG��1�"Ym����7ѭ�&9��9T�|AF>IHL��d���]�U@�)9"�M�ȻL9���W�YS��XZ�[pJ�Җ����2��w����ч����}���~��ͻ�FJ�W��R ��}9��\�R������(V�>����T���v�#X�|�m�Q�U7�����nc��vMѓt��<.�.6��8���@�����8嗜�IC��Kr����+�;�WZ@/�yͶ��V2v^f�!o��4���̦����Z�_�qv<�������Χ���
�� �R"dEo��̕VLpV�v0���$��)0z��R�r�Q���t�����`h��d��y���q��e� �����{��cǛ/:�K�Ջ��ȋ)(c��(�,���ƚ�v`�'9X׶�e�uY�.��O�DٟKM��A��J�c
�q}��2,��lΒ�i��|��ߑ���&�YV���[бC�^����S�^�b�b�<�zb�{A)rEC]��R���
��mĚ/��E�;B/}'�I`�|B%�+����w7p����������g�9����[C�+�ג#"��s�t&�/� >kۂz5�n�Oo��y�dH�:�>Y{��f��fL�YG5P�d��4���]%`O�F��|ƳM�X |�C�M\�b�2R��6@3~�n�1��s���TW�d85Ά�%-9'~�N�
j.��I�jD?%���N$���Ef܃VD�L��>��#�A���֪�WƼ���9�B�U3�eX�6[;��^Fρ��:�.u_�X��)��=H�uz�]��C��Օ�jj�$��h-"�!CH:+3�+EH)V��V��W)-���ۂ_H��/��P��k-��s��uR�?�+����P H/���V^b���~`uk���W��]<�	���7�-C����חe�����&�ј��7�i�&v�i�2����n1|M���H��k˵��$�ED�y��=�r�"n�>hq�ؽ��ڜ������ƶ�t2�5q/�孰�E�{�i��Ad���w��_<���Q��.��f�|�5����5(�#��|���w��
֤�Ъ��#��H��($�CT���2�9�\�>0�%�	M�^�P��T�l;�*�@)���]�z��mK��� :,�"��y��eRf� ;�9|��6�S.�G�sД�.�r������#�J�G!P�3v��̜N��O״�^*��żo��r��ll{K�/;ji�Z�#k�BR�Ƒ��c�H�h�S��z'+��9��ܔ)� $1��g�U%!3�W�@��£���m�ޅwQ�cEY��0e�F�55H�@y'&
z�68�sY���#�ڈ�o͉5���[(�X�R���檑#_ rE�_�RF��7���)�|z���J�'��z82:�O�I�=V���_~��N�y�Ķ{��=���tL�\����s�(����v����5�O�lh�Pn��GA�n�1�h����OO,Dl��$�]jJ���WJ�J�ֶ��9����?o4�ZgzA`�f�Kg^/���q�������=�]�0U�8�&3XE�A��J�nN�z��<�D������a�������n��Fzut��O�tJ'��P��?����LE@�&�f)�e���ď��"P�J}�5Xȕ/{�V�ஂ�Z��J��j�ĻBg�?�k�۝�F��%9����q�Ղ�[�	G2Y�sP1}��[������[�$|�Di�'���횉�RX�v��ȱ8�o�\Uސ_��PB5����I�v�����S����OM���,10��e;/ŗw)���J���TZcU�*&ٖ��)]g�XoD���D���  ��o���[�aQ<�?�`�j|�y���E�D-������^f�o�6�|�-6�L`l%�U�-��� Z����d�8��� ��a�P,��\��&���;X܎H����8ֱ�S2	4s}W�@y���ˀ�i�w�ǡ��
��~ZOn3qҰ�N�>|՚Swv���W"�!�U������pv����
i6H�ED�p�MdE��W�.Gc�O-�Ck)�M�C�%~�"[S�0a�
�����Q�O6�(V��D����0 ,�YI� ��x}\�T��9���v�3r�8�=J�x�Y`��Z���m��+�%�0=���+�h���0�Pvh��YZ	J~p��A�Ƹ�ǖO�Z���nd��#Q$U��W����,OR[�{Ff5�&�T��!#�x���F��/%9D���TM�`��ټY�'�䏱�5
���?'dh�JL���E�4L9n���ѝ=ڞy��?,�el'�*ѽ���Y�;�!:-��*R��^�[)�l?�������:.Q���[��c.#h��޳(΃{���Y�$$�ɡS[5-hY�B�4b�/X;QKEM�%%������V�~_`q��{Ʋ���m�5�ju��4iI�
�/�GTE�`���?07�.���=]71#Q�i�/�Z��ű� �,g�#����k��;?�� �#"��]&���V!�@G�(�?�e���o�h����{�v#�|�Wڔ�,���t��D��i<Am�Qc���J~����*$��8�l�떱�_��U�o�'`��v �	��
L:H$܃ܥ9;yk�a�%�n���N�ۭbƟ;͵������ir��Kc���u����� ��ٗu��c��l~�|Ҏ��͓�^4|����ML(���2��� Fl��h��_�O�':��H脮t���6��Y~9�D��]R(�kJ`��'�$�H�g�]^�(��*�O���7�\�ւԥJ�����m��M�����GD�ڡ�ƅ>0>�5�]�n9�[)��E q��!U.z�- ��T���3%��9�3J�d�F@b��2� ��-hoz��'~)v���0{u�|Ay�)����r��ks3��T����.h1�d��7���I��L~�6.ܿ��J�V�m������F�✇���q�v��+��'�Kz~�9(D5�5�cO%T��;�A��x"������L�x(Dʦj#K	`T��S�`;���s���!��.�a,����"h,7yӠ~����XfVS?><�[��@�����d�ȱF$h���U�
��|w`To����Z�r�"���������]y�f��X`�'^&��QofV
{~�~ۺv�~�6����w��b���ءb�ר�.
J4O6��٢Q��M�-�Ƣ��ѯj�=<g^QI����B�7���&pT��#Ǐ_y�d�]����
O��_$��r���N-���t�� ����]�@b��Iq�[dOW�~,�zMj�	G ��A�f�`5���+����jЄv�y���1���H�3��'��3�s��8̒��q%	XQ�C|�^����"�	��|�M�Oy�GtT��>f�!w;�F�_���/��e�&�ނ�P��:7��49�I�`��Ơ�<MC�P���q�˨��ұ $t�����(d6��;h"�}��z�]w�Jm��:��m#S&o�#�,ꆜ@�����Kg��oB�]�� ��d�Eet�T�T�T���O��,�%X�:�b�|ǘ�qu�M�Z�5V	GG��S�n9�lؠ!�s���;��\ٔ�r5�`�f���Ig�!�M�e����C��n�Y?�_���^���~).��S��F�3<a���-�ܮ�`�d	�D��X��Yr�����iX�U���J�^T^�Iu �t�R���_O`�_t���LM�<�ق�z�o�h���)�>}~u���U���w8�~��Wɺor��}�k����O��:]����{�-F�/|C�JUJ�m��U�LM�c^{]����딚��~���N;kF���t��AåA|�� 5q�|-uc�0>�1>k�͵�^����у��yW��10�6��J8�CT���B����M.� �~H�?�� վ����$�= �����iܿY��I�T����1ǩ^+�*"��0���B/�UU�_��>D��Nm��4k� F�A��
*G�x�l_�<?�؉�ڒ���xH%:��k#3�*= ��zr�ĉ���n����8	���u5D���b"}��6l�P��N�N�	�&��T��@��6e)j�����o�ďɛ�=N�V���u
�cM�>��5��}ȍo�#�� ���H��C���� �^�
[ȸC�w ����z]i4k	,�����Ym����O�\��ؙ'�'���x"ϥh�����m6�0�k�Y��j���AH�y�ɪ�(z�Y�!\˺52��}.��]30��_^�>�׀��ҽ�����@��5ϟr������p���^x���4�_(��d��'vP=���:>mʬ�s��d������f��E���3NU�����.�e}VL(��l�j�~C76�&�R�T���7v��F�h���"��a,��
�_�M��1��.ҹ37�����3AĘW�s?�e����R������7���������;zm*� �%�� �k4��~�ԟ5F=n���)H_��Z�LV��'�4���T ;9�[�=�����͋��AfB��V�J�5P���3�0I�df{�W^XKVM��8V�exV�DW��;���C��bm���Ϧ�w,W��J"��1[Ax{�_���-{�o�rj�/��ΒȦ�Ԍ0�(>�Z��S�J�ӪjTO�u�Hm3RirEMN��5��L�#���`�+�{��9#��DYS7�%���<b�z9�}҆�+j]�W^�r��;��7�w��Ў��d������?H�i1[���L��I̡D�+6�3_SH�ʅa��,d���hmփ|,���ን�h F?jk3QQo,e=C+��x�����V��U"�L&��T��?����$��g9��I�H&b޵H5�N�~t��k^�k�>Eޢt�N�V����)�Q��|�kh�U#���q���/_1p�^1�rdQg��{�tJR���%*,k����_LJ��}�*��%�L�뎥Gyy�u�73���� $	~�����
����Pi�1п�S9��ȯ�܁Ri�l5�����WcG~���Y��H�;@5ʌ�.U(MJ�PYE��j�['�;)M�X.P��
9ٜ�t��A,kЊ��5���*΃�[w���`���M�����5���
�2�^��Mvڶ�K8eSA��.�Cf���jC����B�Q�Nn����&g��3B��4m9��}�d|)��َ��F0C�$�f�x��k��S�@Rݽ/N�{; �$� {̺�3��@��)k��Ss�z-G��*5#b�����Z7D��ُ�.aJ�*Fks��S�g4����(7�oE�f_}�	��m����˻�wՠ�DW�������|�돲:��U�����U�I�3rq���PA�u���kӰ�A�	EeA���ܻ�����/?�9y��-�$�p�<֖��,LV����|�[�{��rA�
 �+/T���P�n��V��gv"��)F6/�k�FY�ʖ߃��:�xns��]��Iؤڎ�6��_�	�^֠��6��:PX�E���>I��x.j� ��-]��L_
����n�㠜!4K������Y7"�K�Қ)f�,�È�E�����}U|ț0\g9��Ex�!�+R��-���aG����z�?7���Y龀-7A��/W/�O�_�8��.d\\2KshA)l��QQ�@���������i+P��;��fn�O`�a�6�ĀR�Τ��2i<�U��vY�A(L���y�}ޘl?���k� 
�%1��i8��X‱�E�R@��)�������|�������AtP`xe��HG�/�FϦd�ZG�S��YKHO�T��{�#:�]%�G�♺~�o�ˆ ����l<4G[Ɖ5X�LଃB�|��e��]X��Z���kw�'�&��ݥ��/�L�:/�2QYt=���t�7�Bn�J�b{�z����]5T=��>�	�����i��[a�������	?���+�b��#5_C��Ҟ�Ɋ�禸J��'�\����{8�Ug'���i�rR�2��$7�ŕT�@�j1��{�A,%��RA��	T��6o�B�6g���+�Uc�tPoלh�6�pn��kx�6'nd��n��V�UZK�^�C,��|��0�(x�u����Ki���n{�_}��4̟��PMY�g�+$������%P�\��%���2�n�T���=�<<!�239�ӓ����D=@�H�q�#<��K:���Q
�'��\C}���u��uݐ���_򿪻���ឍ�U������Z�B�a�w ��I{��%���t������hw�zq[ݧ�~�s���'�*�L[�f� ����u�<��ЭgU���g�CO0�����+������/���&�t���|']4�3vE+�4J�N=��c���/}=��O͒M��~o�<����00]�ȶ?ݫ�����la"��&I�u��4hl�Ki�Rd��Aw�]� @GH]\i.�4$Z�[�V�m�>g����=����6���l)P}`n�>��ʊ�?�E�H�t�YʺV	\�#�&�b}��7�˴�y�F���A�Wl�����E�8SA�`����9�u�A�(&�E6���#�V�ZM�,�(����޿&���i��H����N,�䁥(zt����Ԅ�R 
���ˏ�x��y�[�#BV"NM��&|O�l�����ڽ��%��^w��qx���n1FJ��8+��"�ŕo�ƟN��G���J��>����e6������ ��J�bR�듮#R�����߭?�3| ��^����n���n��S�d(!���G���?�PaO����?�$J�4�o�U&I�x�/]�j�Ӑ�*�m2R����~r�L�o]�-�+2q�%�7�t����u?�lti�? V6�<U�x����[��	��^BF�K��_o8���'�V�MQ�E1U�S�o4��Cy(PP�̖l�J���2�;�<��%��J�<��I !�!�w1��I�l�_P#G:�(z�y�$�Ld��\���qVz�B��ɉ�j�Bm�ŻU>Y��O��*��3���71�>�u�P��^u��ϠJ;ڊ�=�2Fv�|ު�]�PĦ�n�s������+2�+Gf�9�cU��b�\�y���Y7`n ����=L����[/�s������>��|�e8��_r�L!�j��,B*}J=��2���<�L��Z�1·t��k*�� ��,%̂ �x[L�\�'i���Ӓ��.3�ߞuww�(I뻮?��LP�U��zYO�0�t��X���/�S��j��^s�����HJwM�a�{���9��2К���&N?O
���:�d t���,���TMdG��JFE���qr��KUo��i��yW�tLz@��
.���K䆳�4L��OjU/;���E��}�i���am{)��Ԃ�"��	��x�\���uEs�^��&��̉��K�8��p�GAİ�ổ"bĬ7�S�j#�
s�*c3 ]_Y�7�ZF�A,�w�����vb=l������_ �U�Z��W�\ E��ub3f�"�]����w"����n�j#��|l�r��$�h���%&8O����������k>�e�:78ٝ�^��h�- ��Z�Q�my�Y?�+]�i 9�o����@�@�%����g+�3��IlФ��q�?���*���-
�,��m��SK��|���`�y�[z��՛~�*�"�Y��F1�8��^�>�dJ0�k�R�E������C�m�J�g�qJ˼u�c�5�ז ����9IX��0�r��ʈ^�	���Kf�b��N�C���*euE�R��Rc%V���k�8��mu�d,��\~�=�:*\I:�G_�ix=:�e���NL��G��q�{4�p_c���k�UZ�S}��<��_&D'[��5�VIel��q`m�ǅ��4ŉ+F�H����;�H_�U��@t3���+��C���E&o!B­Є+o(R�f��|⳪�������~�Ź5�+V���rҳ=I*g��_6;� ��w���)�e&�C�ԡ��E��d�7�_xƃKkKQ"���@�r���7���=[�U̧+�L�Os�1iS�AA��~d�}r�,[��S���Kn3ߕ.^1u~]���p����U����p-���K%k�|���	1�Eq��3fp����W�� ����g�`vW����6ԜW�(;$>���ž�xx������n��D����N��薍u��� '�m���F�3u�j�L4���.9��Z�eR����c���{���^�'q&�� k{��o���^f��vT���+*�<���A2 ~�*Q{����U<�l�J������8C�i���1��p���|8�K%r�)��=G�>�1]���ຂ*�ޚ���@�z.C?��:�D~G"��;�S)?�^L�4�5ib��Oq�m�#S�rGŗ�aV�LC�6��E`J�;OOu����u���;�m�:�.�%���X��*�����2���bb^n���rɩg,�0�G6w% cV��|��$�Q�ޤ��&+QO�&ׅ�]�|R��|�o8�� �5��qT���Y�PR���t�]�� ���1I1�2#�)�EOw����d�W����5,j�s_$����t/�ӐV�Z�l\�SS W<"����p�y{Y�Ҝb��xW�9�E�q�5���34���@����@��`��� �w�kF���+G틉�
<s�')'�@�i�o�	��5ր�v�G�?�q����r�kie�ݙa�~\y�3���$)�����<N�$�C�vf��bk�uLh��1�'y���B���r�+	n� sEJ�qI	%��Hw�B� ,��`�B]��͐�>�5Q��|/�-SL�7[i�� ���j�D��j���U�4	��e�*� �Z@����逻qE�Pz"��o�7%9W�2Q�ة����Pۤw�i#�rۉ�Os��J;2�$d��<�g-����]����̳q>K�G��f�ƙ4��_=q-�ؿR�m�O"��`�Y��D�!�L�:�i�%(t:W�܍2>m��|��
�ܡ8�:`��G�q�#�)�� tjT:ٮ���B3̀ņ`���(9���7^�30�
��*\�4�~��L����o�PP��]�kD�*���8#ԭ���!����r�qTфW��:f�7Hͳ�ى.����J<��뢮��w��j	��rX[�/�)=7���Uq�gs4p΢H<dh���q�Ǆ%R����Lܕ���k?������Y��RK;�*ۀ��찎�m۠���"^)i�wx�u'̋�!Kڶ�� oW��-�<g��c9�b(���Y�:�ȪL<It�[���7JԻ���g���΅��,4����n�j�p��D>q��^=Y���d6�������ւ�9�"�\1�(w%��b�{��q�;n��;v	�Z	ǯ�0�z�Lh6�U�ѱ`��-bgnu���t�[�g�/�Jh7˲�	�n�s� ֱV�g����&��7��|++����2a�!f��B�>����^��yuҥ������Lɯ�yEe<��yڨZ�1:�}��+Ho�@��h5%İ���#qU e�DP[��F�P��XI�M��`�7��j��@O3����U�<w���b寅ꕜ\{��T�Y��&�K�q�)��M�\dU+�÷�}��&�b�Sy�t�M#xY��X0�ȓ�؋�8��|���P�Fm�����T�����Tg�5r�o<1`|v�����x4��a���3[]�X�C�d��;��O�W��b�#�En}];�5�<����0��l�9,�	�Ǉ��y��[�^���%�BI_?�"��
Ҹ�H��.XO�u��csaIbŎ�ـD\�g?Y��`ͨD/��t��/6uN�a��EA(���%S��GyD�����	�+^ד�\�@�5m=UG���KnFW�j��\)� q��q��P���Sي� ������o�����neH��:��E��KWz�����E��".���O��9"mD�o��=ס������j�Gq鵼��V��g;Z�kkB��]3T@�N���.N�j+��Vd������8~O��=�K�������,1��Wkw;5&Y��	Cf�+B�~ҒÀ�O�0�ڵ3Di]X�A��Kf�_�`s~�>`v
�`A���W�6���!��J7���w��CK�-�{Y��$خ�k�g'I��A6��uF�S�ܖ�2�v�zw)��G�2�
�V��:V���}��_Zq����cڠ:V�4��V<�h���l�zC� �OQ������i�σ)2�,7`z>����
���˚u��<����KyCP�?2�*ӊ�bq:?w&��J��[����S- �������\k��W��{n���X�@5�������U��y�N�.��c�Z:8�a����-Q�ö�"�M���f~]��Gy��f�6���oͲ���з]��♰%"mZeӯ7xFm���Q*�"x<C�����`�:n��o�F\U|����a>	>�8�B�@e�u�`���,��O���o�71�!�h����.��q�����rs�+r㸎���a�8���
"U:F0��F���w>c��á
o�FZ���B�gm6�X[
&��6��'��/�9$�ճ^�8)d����79�B|~3��{������B��&f](���;o��R�%u��{7_*�+����ϩ�J�{d�X�}����,�ڢ����ܩ��!���[���o˞.s�s*�B�c����@k�2�Ϋ�u���B54�9���Up�Ss_��?%�0&�,o�=�u}t� 'ɴAޭZŻ<���f����"0{LF>��js������<z�N��	��w���U"��q9�擴�����	��\�J3i�mk�:�-�#Tűv?����
uN�9hv�D��K��6�+��Y1ߞ��#&5_�bm���R=@8�5�:��͞IL��*Y���=ī��oW��Hvy?���&4�=�L��p�ZQ��Ý�S?-���S%Z�:��Ͳ�
l0�,YdZ�� sfB�T2VU�i�?���������|��2�H�Bl��]$\��`���3+�R}	�by�d�ߝ�y��MX0"����s���n؝��\����ly�*��wPKS��+�Q���l-��1��'�v��-#��
"�(]��ʦs�=`^=���[+e3Ȓ���־>�,~��
b�7����Ĩ�{X<�Ƕ�}�v�.�.A�pW܏B�09�]	.-��JS�6�y �[�ۀC*H0���iv)�̵=�4�\ײ�m+�݂A.ί��֬� E�� ��=�1�_��ՇF�0	�h��:�l�qm����Z|x�O��']��K���V+@�$RL4��_���)1�t4��n��W��_�.Q&��]�-���cbC�QC�k
�i��X�a�9��'��f�m33L���$yr�o-_XG��[�Y�-Y�f�v���X��PNh;��]�]��K�v!��L �����͒����^=&��4���`�Ż�X,����^��I珻Z��I��H� �(u�yn��HӲ�\�Ư��mL���Mfm�!ݖG�e�>*=O#e4t�7��<�)�^}��r{����¿Dc9����^N	Aa� ��
W+^m���t���'l���F�1u.J�zO���=�L򧠪L�-glL����l>s<M�~?����f'��s!0�b���h�ɠ����,��K�-��܅{�����Re;w���8�jQ�̊��@H�^��f$�vR�E8V�tA�C����'AR��7^g	F�mܛi|�XA@�i�$��12f���>RTL$��4Y�T�
�lQ�Y����?�P�
q*���ۈ��+n�V�3�d��"��8�[%eJ
�NJ\q9bPC���f�P�Y�u�M���A���Z�`�)�s[@)���n��Ӧ���� �S�1��bt�H�v�ןXj���� �ӱu#�S�1�K=�sj�z/�L�	&�;&��8�>��bЦVK&ыy_��+����Ƶ~��c5�i�+v!����!�s��V�8�5�M㒦�],�ܥ�`�[~񡅏4�˨}n�����9Iy.����ސ!�X���'�tGPp4�`�8S�6�=�cd0B��qf�W-�g~Y�s������~�f2�I�ANhN�ȑ�L)�x&)����sg�����^h��S�/�v�#9}���l
���C?v�>�>]'13��� C���Ϣ)�`5~�!��NWO$��;������ц��g�Ц*f^�}�&7Ӧ�\��7�4k�ⴺk-��g�
,E1Xz`e�	�`5���� ���cM��#Գ(+F�[�;>�rД����Z"X�r���ћ=�~XzY��+aܠ_�Y&����V�Ժש���4�@�-Hy���*h�ԫ�N�`�����ES$3\7J
��7Kc+�b��]h�����e,c���5�2�v�=4�.;��o���YH́�^�B�#�a�� ��OYEmǿw �㵰�\gI�u���� I��g��I=�@�F�od!�A���	.�0��c�^����B�3�*E=`�6�@x�ؽZr���ݲ�����Ei*:j�;�e�T�0�?硁���
"�-@���������jY
�ʓ_VU����`�K�67$Io@���=�Df6���������e���LK2��(����Rl���;D���V����l�E�8D�Dn�U�8��'�]�so"P�����{��Ke��6^8���e�ԎAF�|�dE�.��O�dJ��C�ׯ�!�&��2+�m<B��mۦ�|s��C̦�QC�Atba��'����hð�����V�)�Ρ��ha]G�I�PC'��g��l�su6�Z�ش�U�;AD�1f���^�r�<e�Qd���,���A>�Rw�n�����]�\�1�Z=������R)P�g� ���g�wq����P4��9��c�#3�u����0��Js$'�_�ۻ.��&^i�t��S�N���U��d�0�T\Y��^���	�N����<����4�b�U`�0�����f�F�6����}�đ?�8�A�7��"-�𱉅�ܱQg����_čȣ��_Sz� x���E��o��Zx����*+��.bl�q�9PJńG����g�д��;H\�%��P`�hsQ���[$��&�ZG�J�"Ʃ��,f�﫬5	���9�p[�s���(^��aP��b�s	;	6�M�ۢ�sF˅�ea0$��II�n�C:�H�n4�S�o�̢�b}R�`�7�s)G`m�����6{R| #��_�KP]3��hbN���zx����t���)q�3ysF��yۨkY;'~���V��g@��7�\�s�?:NS)t�ra���%���<��J�>/>n(��Q{���{�Xn�h������#	���UO-/�Y����{DZ0[��������σ��9�J��Ƨ��Y8IM@j�j�r�4��Z�Rɲ�j�>�9��t:(��A;�\Cє��Y�ʙ��>pr��J\F����!�7� }��RP!���1K�F�ޟre����2H���ʱf���>U<ߥ&����Od9�����rw:	G:'�E<�m�rE6I���^_%��I��d�bu�]{�j�C�O�ƛ�]5˂X��H�|�	L���G����(x�-f��W!�Q