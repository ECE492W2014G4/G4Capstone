��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P��v�"<ߞ��&'��k%P碶�R�ӣ�sĞ������FY&�S�~�p)oZ��٤bG��$=���^�I�Ύ��f�cX�O��S�!|��a(9r�7�A=����CQ�j��;5Jd�g�+�*.4j�Z�7�d�����OQ��3+xt�lK듂=���̛��7�)a4]k�Wq��u��hZ�����h�	Y����Z4E���DY��=�C8	t�QeTM`ۋ��#��}������٥��e�+41
�{�,��:�s��
-�\`�1�A (���{S{ۇa��W�?r�q���k������)_�B��� ��S�=^����%�
ċ�\�`C�'���Q��J�P�N2���@��W\ԉr�ۓ`�Z��g���^�-G���X��2�m�t���T�Y��*�'�^���ӳ������]̴����30A�i���	Ĵ�Ժ5���1V]Ь�N�8z1��*5��k��NZ���q(�I�5OB/����f`�^G/�QÕ^j葧��z%h���sQr�Ȟ���zg�x!v��L�ns�.YF)2=G�y�MP�=�X��Tw��"7���DJX�q<��G;�"L�d�f8֧���O_ �'w����:~Ï�����/S���ܝr[�Ou���(�d�mB��u���D>�l[Mf��M�Ĩ�.�;�
/90�{��p}���w�OO���#���7�O`B���(��*��(��}�c��m�s�0j�ܮ&0��Ld�kHtb{wڜZ`դ�|m�F���3�r�b
���:����K��}�B���//5綨e�A���9�j4n�bu:ph���_��)��D{b��;�xk��X/-��P;]�� �y�ݽ2I�3�皸:~�o.Z1Y%s-@�G[b�NR�ۖM�9۞ۺi.μ��^� 	�'`Ub=�	�Hr���9�����c��\5���]�7N,I,Y[t�����\S�~��iJ�z��ҬG��T텬@a�����/�����2�X��j[�������s�"&W:8����j�[.��U�w�b�������o��������8q.NpT]�"?�a�˪���8��j1��x �?�H1��V8�8i����}�b�ޝb,\A��H��� Qa�	9=��UA	�5�G(�=aV��>6����]oo��K���i[��;�ٽ��Sp0409�%�Zl���(t�Piva�"����n�BL8->*:D�uy/KW-��w?,}W�?lͭT�1ziF�K8D�l�d���M�� gm�B_|x��LXx<��#�|�2�Y]D�c+(�m2�:��~�0�S��Dۢ�T�H�+�)t����Zc�J�k�#� /���'v���i��p�+'+��!�:�!�aQ +=uD�e����O��{���l�Ɨ�ؖx��	��H��2j��%J�Hndh�*��`���^��Bi6�(���(���F{���`���;I��!�h�l��dF�W�fŌ^`@;=TV6�Sk%����S�֢)`V�t�Z����{��|Y���Ͳ�l{�:���i��ד���^��-