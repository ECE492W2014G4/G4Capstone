��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P��v�"<ߞ��&'��k%P碶�R�ӣ�sĞ������FY& �c�]��bh_��I��T�i����K�SH��s��S*�i/���!l�,�D��R�	�+�7�t(���n&�/�dqּ+F�l�	;;?OH9Z���o�v�����n����->��U�^/�+`6�$	V�I�p���l�&�	�M�2��s�(�,~��k*�<?нyD��X�k�E�"\+tt���zbU���Q��{^n���]���**����rґ�h���L뒆k�����3$�:0։q��V�]g$��vB|��fN\D��>�0H3X���68\Pɮ\��w����w�e�ZBQ7��E���\�#�zQɜ�
  m \R���~���RF�ңD�9�z[�ݪG����D��H�N�	.�	O�j�~t7�]�1+��$7���6�(���(�ݿ�?�'!����g�lW�\N�A�ЇW�0=`A��tc�I2���s*ր�0�>����gH�Z]�D�q���5o�+Y��p١6٣��$��[��W�ٽ�1��D�"�+��e�!�C���ͺn�C O�1B�ĒN�G����2�� �%X^����x�j����ltg��"`��"Ƒ�=���E}��g���So|�SJW��)�*V�:qm�v�f!B̯׊u_�N�@Kk�<]�'~��+��a��+��w(�CL���X;�0[@U>e4]԰$~���A���ר�G-�	���1S�:�W����{]o���bG�|&�x�t���ԣډ�pM�P�����뀳���;��0�	.m�G�ts*�X�w�]_�O?g�5u�Q��~��h�qm�/Ns"��>��I�B��T�iգ�x���5�wrX ���KL�����c�8���efB)8��)T�I�)�_���F�3ͮIK�M�ֺPO�}��A�� �F���|�!+���Yl%]�Z�Y�'�dE����X�.���vG^�-9�1�����]�oҞ����b���Ҩ���f��x�a1�+�K�r�(��0ڠT2�(����_�8���wV��G��9���aK��&8�������yaBW�h�M����N�0�Rho2�G��Հk�43�B�� �6�VP����%�6:�29u���V}Öp��yx���M@;p
��|GәY8y���B�C����v�u¾��|F���x�bg�`�[�8-�2T��?�4��6�ɐd?��t�y��/�
�C��P�����
���	�����E�Q�E=|#�T[3��k�8oݎsp�V
�0%��%ר����ڛ|��Չ8��l�,<s���p����U�XU����ѡx)�3��� �[*#7�X�W(���Er�.��ʴ���U3���@H6�hQql�?�j���P�8L��3�>^�{N��������P����z�Ņȹǅ����ئ���fG��=U�Nbi!�~��� �Fί=�#�>�����<�EB`�d�P�	fm��@��vZ�<��k��R��^�ޚ�b�V+�%���u�t���S+~�xч�^Э�8n{��ğ2��Nd[=���H�KR.��ŒE�7Na�:�H�Y�
 `Si�<y�5G`%��u�p@X7jr �O�|��$G���;y��")��G\/��Ė��<��+g���(��1��1eE�������9%!��{�ʨ�YXBk�1�~iq�v'Ñ�O�P��Mc&��R1oj��߱��)妪���ȟ\!���_��2��� ���!c����pHO��bߊU��g��[ӴgXyQ��Py��%@����:_Z�-|�N��7���B�&�^E�B�/��
Ҿ��1�o�T���9}�D�.E�{	0z�����Knǋ��.�����6@2��89�j�%����R)A�ς��o�"A}���Y+��_<�p5�~�k�/�_��]�n�������}v.8�lJ�V/�����
������pD�$�B�x9"�7_\mI[�I�IM�p�\�`�,}��\�?*����:L5]�z��1~�:�)��B�L��lD�/l0��񷈐����*8��g�'��,҄��p�x�ě.��Ḳ�}�o��e��9��/��\>���5���6�7eЊs�i�x���ƛ �z���-�]�;��w#C�e���)&L��o5��(s@y��H��>��I��*/���b>A^��q���R����j������x�	��I�$��qyQ��L5���N5��
�1�w���1.E:���Fʤ��"s[(����#9��}K�b����O�	�`�Y�N�����Y�k��7!��d���4ۑ:���(�sՓ��&���
5?�{��Y*������ȩ ,�dgn�|��,�U~
�p7�3�2�浱���[�\�L"�7��
@Λ-D�J��D�3T<J�;Ļ�| ���Xf�����.�PP�x�x�'7ׄ�6"0x�9�.'d�s#���:42 ��LX�u����D��Ԅ�PЫc(������ȶH�\��аv�����d�����!IM�}�/�
���H8GK.ā���rY�*�&!h�0 B1%�,�p�6��V'S�V2��j6nr!Î�O�0?y꡹�B�|�\��W=�����MK�pM�fB���+��h;�p��������χ3|mg� K�o��=c"��J�;v�S�q�iԠ"��D3��X�S��e���/B!Z�l�X���K��hs{n�J�Jk9 �{$(Y$�ӍH:S#�X�0a�~O�V$ob�#xCK������U| ��k���Y�Dy��/:�P���%#?�[�:���n���,.h�#0$��RW�R��^�����S�3�cd+�~ʩ��h"�A�^H"���J��C{<�\7���{͍P���y�v'd�G�@_�����d�
�e��3_���V�Ab,(���K�;�=vh�z��QQ<��5���劎��a�נ�ۑ��$��E݌ēv��#�}X!h���5�	D�3��C6ȝ��"ظ�b��؊ӕ��c6�V��=-$^`Vr�?��P�#� �N⦽%����8wj]�X�l��T�̧u�%���^q��bv�կ'�a�Gf$^8��3�AI�}�r�lؤQ��W������j}n�p
����Nخ��a�A�e��K����>dKk��	�Y׻��M���� Ǥ�sm�^xq�3�]W�ߛ*$���Lk��?�]ЌT�*��:h�6�_�H�n2t�5�_�#���K27�.��f@VF�֊���%V Z�n��#Es��gwt�6D�������K�O�����\���GB��b'��W��G����~P�].�����r�>�np���%�~�1ȏm_���:tT8Xz��F���K����?IE1x��PI�`w�_��;��I#2����}rJ"��������T/���w�E�z]ް����&�5�3aƷ��1S}.��r�Jx[[&3K�G���n�Kgը��M�p�Ln,��zh��?�a^Or�}��ai��x��P�}I^�������������f��w�">,%}.ߊ����{���{MHt0��tV8je����U2E���-����7.�����v��@�;\;�c�+�g��iP���E�O�����L�u����d�9$�a'�t�;��3h1$��۞�X.�ߒIw'<>A{'?��P��_q��ڹ/~>�C����@���� � ��z4YKD����о$y��G#5�Q�292�~�

.��X�>���h��#�h#�Z�J�tY����4ִ���2�����|�d�\�[�ܷkuQ����t!AQ�z�a���^}����J�*$!W=r2�����&�L�'�Pʴ:�t���b��;f�2��F�a���g�7N���;��kh���c@��q�4�٢jq��^
7�]5�aX�x��_}M	?M~�;/��il�Lf��V�,��g��T\��a���(��a���S3KqaǷf���G[�N��
Ѫ �q�҂��ʦ	��[��]��P�X�;>�� >Nݫrm��>�S�Y�-q�/�q�Y�vL�k�R��h�ۋd�6y��ȕ�����!����mN�� �~?s}͋Ab-�)�����4hq_�[#:�9)IB�廳��Z�M�s���B-3��:m��.y[�e5��� "<���q��@N�Y�a}�勒�vpPU��uHѯ����=ọS�!S��J��~���{��?�jZ˶�)i�9��9���	ͨ2�BL�����s���U$v���i����$����]�_���o��)��n2U���r��($Yi�2�!�߃��N�.s�9�LcJ����HH6��`A���DC���o("~J)5��J�FT�Z��R)πrA�\�p^+mj'�z����������9��˭�y��$f@��s��悀��0��{�n�h{�ڊ(�����x�����0��B�<M��X��sy�#S�`�[�U��%a�� ���R�"��R-Y�Wx:����h�C3ĻeN
X�O�<u����{�/EG=����<�0�Ȩ��-hlã��j	`G`eY�.n�/�����T�`�GY�<��g6|_��'��(:Ĭ6�MT'Y���+�ǥLa��l�`�mm�O�+v�k�k����T��޶�`���k�z����S���^vJ�)�Qd�,f��$���`�8��@�}V��),�=�*?|�[�T�"v�w!�cu���e�P�!�A˻Ƹ���������s��)Lݔc���� V4�VS� �޶9����AU%��~`�b~��@{H��X*�4�ox$�W ����Ĺx��o��\���[�a%<�\�(�i��s:���d�af�IoNV��fI�D8����wVX��G2��Efh�����<��Z�#'��׻FŎ�m��Q�;X�;��6�>�ʶ�\+����T/z�nm�@%⤲�:Ϋ&��ٱ�t�O�bE���]?�d�;�Ew�w�i��[F���򚟎sG�w]�[Y�s��pYn�9Βh ��[�F��ѭRlp��5�7������ݢ�p��Ý���.���1�Q2	7��\aȥ���|���3����	�~�g�*��ʋT=O"P@ԬO�uW�ڱ�bøZm#�t~�r��^���[x�:`�QC-i�N��Щ4��}���W��F�ܳ��ړ�#����w�#�����K���aFW��Qq*�:v���EէH	̷��9ʘ����Q�V�ؚdk�,�O ������3�	;�l� �i�P�P2~�W�R�S}O���̷��*.�PXɫ1N���ۃ|�`�W�xل*�7�W����_N����!kk�Rү���l�R�����|�9.�EM�]���
�ɹ�F �^����^K���e��աH��)���.D�ɐ�S���K�.���P�A����i���E�J1���83�$O��`�n���#�P^y�cs��-�
_��5���5�$rX/��T�s��+�Ѝuf?�h����RR� �X*~ϝ�>P��>@V�����ˠ-�{���fR���J!�TP]���ٓ���a"��јg5�	u��7��9��YI"Mo�?a}����%lPV:� �@ae��pgj5��0���_Z$���UKq A��p�����e%�}��˂��������=�t����\�I�V(�4����>��]U
 ��0	}.;��4/�(�~��)� ���z&yF�ł8V�ާ�C�g>DPK@�x�v���À�}8f�cW���<�HO�qβ�(���Jt���u�z׋9z�6��oTsg猺OkI�-���/H��4��x1�mʍzys�)�6S���j]��s�a�%	(���}�>9Ҟ��&��4g�o�t�m�)S�A@ �4!�,ً����d#U����r���|�Ҹ������r�
�t�n�
. ȩf����ACƱ���.�A��F��a�U���{3I�_*0���q�,��v}�(�遉nB-�[��C��$��