��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>��`HX����5a8Sjf�&���>b��z�P�͕�[���O���,����9��SF�ĪZ{��A�jb�$�5!��^���4�G�hJq=`��@E��G�В�Al�E�Q�
E���'E����8�j.�V�*�.�Ҋ[�6K�Z��5�Ιjγ*�P7ۮf�������������n��J\�Lt�4�R|�{�PE0|+8���=4���ۨ�˪6�Z���� �Яb�Z�i~�Kl�T|u��ʤ�3f!��H�:U/̑�����Q��iUX���_{��i8�<�֣�[���j��i3���5v��4��R�����g?/�pR�$�9�Ug$��Ȼsw�$�7�X��d>���D�Vm{��}�K�� ^7U�:�Ac��$o̾�T2������d����]����4��o�{u7������M{yU���"lM��ET���-�'.T$�,���հ��K�?wpPb:�V���3zƮ~���%jֿLO�s��Iښ�a�ß@�bcY���ڰ����X�ǽ�P�pFj��d��`�FϦ$����Q�3��o0�T�eV1����R�%�J%EKzm���ʭ�j��
B1���%39�re�%%NT�g��-y�ˣ�r�L��"۫(�!W�ݧ�J��1So}9Z9�_��Й��TLXU��N��U�)i7��$��f��n%@}J1E�R�.z�8�
<%Z�46����`T���z���'��b��S_�-�T\m���'�0��f�'�[wTd�E'�#��Y�Q���2��"�I�Aw7?�ܿ�zRU�����,�����~jp��_D�
��@��x����|7��	����v�v�	z��c#D����C������|b����%ٝ�**cms� �{��H=��d6�@�i)�RJv)�y�udF@���'�윇סk�k����_�� |썟Ԯ�v#W�oxF�a��9�N�,���ŗ�:f]�<$��,�,$��`a_�I&�IP`Pj]��;�m��X�(�>`}Qr�(�j�d˓�(��v�W���7����&��n�Ȳ�A|Шw\I��$ں�7��t��']������W�n�J��3�z��������C�3��`IK�K�Ε�n�y:Q���/#�.ڬdA�\���tbC�L�B���������^��cm�d:�'P�*�>�&;��C����0���2�e��2;s��=a�P ���B���ҽ�R�=,��B=I�1-��_;;�H���'3Q�&YRXH�֢ʫ2&f^�,��!M}��tr�\&�7ъ��G��~#��c
I� a��k��l����ep�W���Q0�P�+5
��vw��[ uKo���T�Ԣ@B�;iMAn� �s�1� ��p'tOu�m�3p'2iE#l�d>7���I�ܦ:7��U��7�`�J�@h?��X���;/>����T���w��f�u{Trm=���¼��?�PF6C"m�"H�`ŇԊ���(5�}]�������a�d�*��*ܿ��pgMm��eE�m����;���Owd��P@c��Y�X�ef�b1�ՅHN"�1ܮ�����k�m���OӾ6\pӰ���<O���+�����bS�>\�+��a�;���f��z:�GI������j��:T]��Sc���ϠZ1u%e�6K$̀7A���QEI���<5����c"K��PLSW��#�� ��F*�q��^�(��~����Jj
����v��W� ěYc}:M͚����~r�>�)�.��of�~e9�qN�t"��`�'��i��	e��f���P	z��Gi�(`]�T�ρ�e��~�=�f�*QT�&L����õ	6��/�ޤR;�n��!Ksp�k�o�1�w�B�.l>Q(�w��I�Q�Ua�\A�XiE<���v�q��Ϧ��š���y�C�����mD{�p�V���������邼+�9�Z�;��Q�l*��L3~�d�K� �to��Q����)�1����\N�Mj��栝CNS�ͣ�lex�w��1ʰ�~�@��1�T2�@�N�
�:����$[�?�dUʱ��_Z9�m|R���P��vBҙ	-Í�������l�3թ�*��(��/�8�Qfo!!d�(�[��mZES��3y�b��Ⴗ{��<�qVC��o	�����ס���hV@�pS��r���)9��vo��n����[�M���DI�@�y�������W��d����� �7�8��:�8�.M�7�*RX頻�7���._+�m�+���8�c���Q�	߯�%rfTMO���z��~_���#�BȠQ:%���|���m�R�L�+e	��>W�Y�r~��[��r4.]�N�v�_�D���eE��}R�,���O��~�4�	n7�B����R��&��diV���W4��#'�#�����캓����2���5h��%����Ӿ�U���_��l��5$b�g`d�ٴR�0L?��Un�mh�V���+�=��8ōߥ���J�s�:���1���~(�+E��1�x�&�6��-�e���,�T0Ȇ���1�QK�m�
�&��{�X��\"���B�@�LWr�H��+�n�R�i�l�㵣"-l���%l!����)0~�+��У�~g������S15�y:.e��T��C�Z��;^�3n�<��Oa�u�f$F>\s��xa}���V~�
��x{�^\����<��~�`��ݔ�����sRe�Rێ��u�`Hi>j݌�f�b���Vhթl�lޥ�Fq���n�Zr��;�,��>ڢf|$��ep�e�ИL�D$��׽��=�-��H����\l�叭S���ٞ��O�,ې��K߳�̒�蝑%9���˰�"B�|5��ޖ����o[�����'� ��ZC֒�%��6v}��%�}?�s\��Xn���M�H����.C�	+M5��]G0����I�d��s�_�^�
j���X�ӑ�h�Ⱦu�ԋ�|��c�� ]ț���BD 
�z.	x�xQ���"O��Ei��@��b��쇤�	���D����G`�����컥x������^��!��e^3YW�`��0['$�S��l������)��C�|.5+K�'$��\�*��f,E8�4�5��&� m����)^�,���t�#���<���|�ĤuK_q�ZW��I(�~�
�8|�r";�Uf�E�����C:@t/\BKa�i����t_���.���1<g���C�`��@wT�4
۲���]�%P�t��v�]^M��D���)s�gl��Q����r�o�h�%lx��{���m$�ȿ��@��)�!��`���;�!1�<�^h2`{	, ��X��@ `�X�G�0��H{��f��!8S'a0�?޼��kx4����<��歍FELx������\\�1T'�֫
h����k��r1\�L��*�]:�-z^O��Ӡ��ۀ�����%�$�{���?�W�v��5���`l��;�Y���z��Lb4�N�3?*!F�#�~g��G��x��h���`����~L���3��Wu���IX@%�Q�;�D��<Ž4g�d!�V��<�L"�|F��k�5 ,�yv��8��O��1���k�_nVx6���H����U<:J]Z�Zr��ak�8߹�W#Xk�1�B�u��8t[�E��>q}�C�pAps����ƒ��k&o/���)×��b��@�U�3?�=W$f8i���HM�k��z��o��3j��X�rs	����Y)[%�H�@Ϡ�S0o�T��#�DX'���A���!�lC�P����8~".�U&�ea�[6�8�#�{��~�`��Q���Y"v�?%�3괛o��r�g���SB����zO�s�c���X-�L1�B2?P��	���>��v��2USЯ/��<9X�+���1��X
+Ԁ���+^៦���>�V Wb$��ǝ�2\�q�uX��A����r_'����@���}]� ��_dE~��0�v*ʌ[��X�	��s�	'q7 W������d�?T� /�|:�m����c�稈O������T�(�:V����(��ڪ��0���̷�������Nw�����6Iu�h�:��+�ͪ7J1��)�'2�24o���Ί�È��.��i��ٷ>����%b�r�X���+�����܌4���܊�V�e�(C�צb�W�$�#lK�,[��@���X�ɔg�E��J G�-߱]>���N��E�;�8��d��?J@�5����I j�X����t�u�����~D��I$�i��M�p��������V�W�̊2���y�2�6+���Ҏ�v�O��9����qe[G�y!3�ٓ��/�V=o9��\[�xN���k�s�	����s:k0`�������}j�>��A�^�ys�a��	Ӄ��ⴇ�a�ŅDTؒA��ltլl�6���7> ����:/��g4h�Ox�`�:�P�ܑD�r}�Θ��<M��UPv6�4�; �A�B.��I�q�l�^��Z�c�|���װ�y��&�	�
�(�,�a;���?�?�C�͙��B%�ױ��i N3�$�F΢��d�; �f�Rw��u�l�Ʃ���(��J���oHzG8��z�v���8Z�����yW��G�@�g��o6��?���C�A^}~)��h�N�����;�P�(��MTĩ|�XX���{FJ/>�\A�p(�<�q�5�O|��LJ��dFt��QNO��ぃW��E��4�E���;��t��G:S�2�j�Y3����ڐ[��b��͖]��Du�OǅIRuj�u)������R���V���=��G{�����fz��rn5+��л1���d�B��gV��9A�#�8�Q�7���(�=��1����%z�vf�23���e93��	�1��R �W<��f� �׵uLr�W1������,&u��(aZ�/9x0W����zd� �j���/J+T��e�Wf�D%L뗹�B��g�0����Q���3�|��Vvp
�&�8�W�^���挔���,��m/2"�z�*��kEn�Q��!�c���p�:l�>����6V�����B�T!k�U�L~��\����r*�a����V�T�ߌ��>a%6��P5��>5�D`�}N��Jp{o�X��P���|�i��zg��	��\)mf�I�������MT <\7j�і�T�5&.�fMn-d`g(����m.��+%���F�j\��'ZX���iA	5�H��`T�M��(]:Aɤ�d�<Y���Cq�e.��Uꄤ� @= �C��1����T���س+���Ms�@����[@�}�ͽ��hpB͑E���S_�gH�"�	[ �Իװca7�������Uf!)�1��S����ّy0'}����8F��sɠ�Y�
��bK���>�ڳ�?��>�X��ێ�����d�8p�2�/�x�����[b�.����N�/rVNE1��nP�q��6�_AkQ$H���}��l�+RfB���o�7 ��A5�Ÿ!��L~\æA,{5Jпf���<��s~ol��r�<9�+k#���al�f�cF����Q?U+��?~+��\��j�w��͊��ƃAl74�޷p�8���5��fz�Y�
u=Κ0崅����tI��+���9�"�{ �^�4������^j�4��){i�.Z����tHD��U�� ���P��㈣�aN�Kf#��  �}s&�~������8[qͲw~]�Rh.����3=ab	���p���0�90~5�}��L���_�� H=�R��NJ��ez�j^S0�}�����[�]��"���`�\�`�?�K��Μ��'$K�X�<��F����}R-��d���b�^��x��Q�?=C������v�rE���>�3�����u���Q�t\�:5��*�٧��k�.�>C�fh�D��pњ`B<d�ԶEݕ����2�.��)�u∌��)�J��yԈ���]Q��9�TJL�����ڋ�n&���F���5¤�a�>C���u
Z�޶�P��v�1����\������z�֍�����F=;O)Љg/e��ؽ�cؠ�h�Lp�>Tŭ�+A�{paM;���n�V�x�`KA2�y� �mC��	\��|e:�{�T`+��c��������%	��{Db�NH1�b_����/yUx�(5��(&C`V�ڔ�%�F�ܛoikMb��x'�	Fv/�wR�"��MY��{[-����k��.W�����5:-Q����S��ͮ�di�$����=�/k���<��R�?ј��ཐ�����Y[�b��y�(�7��� �o