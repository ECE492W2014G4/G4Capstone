��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�"��F9s�`&���a�oq���F�g�O�]�<ݲ����eCL��D���{�5��8̝DFI��Zp\m|Q��
�}�6C���UnF:<�jΈ�2�����<����sf�k��,jڙ�����2��X��Ss�HL��	�������+g?���N�Ż�����|�v7�{M��VNB
��Rs�゙�Ld\��X�'��R :�J���^�����kMkx�Q���3!P}�e���Z�Y?.�U{�RP	�)��lI{tI(S
7ZF�W+h��QCCj�X�ӻ��wcG�_. �S�':@A�5z�zLV��}������Uw�)��eW��9M��d�c���5E�j�e�|���F0�A?��W��|��A�Rȁ 1.�O"��v�j��%��b�T��f���h������I� �$�h��2Cm�1o8y��jt�k�絪��e�9�C��|�RKe�AJ�i��^��ш]��N���n�Y���(ȱ���vB�.}��3�����n�wR��Ӆ���4�)�/��D_~����b��F6��e95H�A�ۧ�V����'�,��8��>�[�y];���0�h]�TV��M�%�,�=!�][��	�C8�CT��ډ��;_�����Y��Y!W�����4y�y�Ҋv�&���]l���6]e�I=ͅ���o�x��3,oO�0�i/p��+?�W���J���m}�4SX����"�f�ոN7��l�po�&7훰�W��C *�t`�� �n˸C�)3����.��=m[�j�D���$j)x��q({��r�8��,6����|�*�tl�����!麞*C�2���Z17��=a����X F�q���_S����Y�G�	����Z���a|x���L�����1*+Ǌ��]S�S��3)�`s�}�S�3�������e���y�|���C\�ꛎ��G?��[��m�%>`y��D~�o�q�Nm��ْ+�Ys���G	���1ZR�)��U�ihh��`b�nC!���B
����k�AREX)���h$�I��N(��A��-�sk�H��W���C�%H�TI�lac�P-�eOR�����P����l�*/%�M|�����Hu�l�����x�d��w���bA�?���v˱ұ��w�i�m.��'�*��}�0B� TP���Sk��+T�r��5I��,�"�zd��SX<L�"{��>v
��m}���h����
�� ��Ӑ"��ul70�U��h���g�Z�ɗ��%N=�9��*�s�(]�b�b��x=�ִH�T7��Z��^F�B�]B�̓��3ĔB�4����	_�[���r{}w8<���:pc�aZ\���b9ȡ"'�iK	/��;j�f��X��@���Gզ���U7T%MK��};�t��Ăk���?�41ۯ�u����V�ܵ+���(U
�oK�?ަ�T��N	�����F��KޑM�i�
�+D���� ��]�����h�h1'��%�n���������{P���^�nQ�֤xa-�����ҋ�{�#�y��<��Q4j�X=݉2S�I���d���M#��y�Eƅ���e�-̽J�Ѯ�WA�Rm��u�)D9�A�h�<�C�W�tGb8���`�%������xqG�]�>D�.ɭ���8�֥J� �7��%9���?Tt����l9q0�U����'�ߍ�N9`݄��W�M�[W�%�p�v�Oy0������׳�o��wH�����X_I7CU���9�o��֡�7qx�FVn��g�m���ȭ;m�E���莇��V�"^<�ɞo�*��Jc�߯FD,8�Bc�=�sr"�@�F��5��G�9�<�g��i��<-��z�I�ntuO�ڎc��h�[	��h�W{�Qm*�qr���*S�k��*y��~��"ȋbp���fR	��>NY�r���f�k������7��p13��-jA㣞X�%G)	F�ٚ���S�g_�mS����e,򫾃���牞��p�?n�[�^�d�� +��>�ϧn�@[���M�[���՝'��\���m�~�έppdv���M{H�)��K�<
�6�ɩ<@�����W�xș�>���z�Ȥ���v���B^�#�r��I_j/*��ۦ��ij�	])WXp��:����*�A񐡜^�quߵ�.��[�b3�����Q/��r�ڔ�u~l
[J�1��VW��¥�λ J�ՌuJ��C(i$r��t��H�G��˂e� z����Y����Eq��'�f W��v�CC�W�6G�HOg��z?dZ�c0�u���z4zy��W���
����B�tgVK@�7�H+<�'�(���s�`4����~u�o��2W�]����W/�(-��5B��Cm$ϥX[��܃��%�K"6��Ȑ#��m����w�Zi��ѯC�㩀E�<WS�1�i�����[K����L���r
L�N��=���3&?B�N��[�0�h+��t=�=�_^���?:h80���Mw����B{b�����R]�<矶���9d9�����XP�p>R�$���9��
J�B�p�#����0쓔4���!�
�/�����!���b�FP�{b�X̣XI؂��~�!�T��/��.ҥ{Ѻ�Nգ^�X穪땪�&Qi�Ɩ@}���	���'+�����w�!�,�UH�ᬙ��4
�g�Mͭ�Q��YKYI!��T�#� ��
�\�r�j���,���4��Y@�&�vt���f+>���{�P��l\��}��7'D��ʚf��J����_�Ƥ_d�˩�>q��p�}gyEz1*Io�l�b�ɑ	B">soKF�|�TV��X�?G՞&.�&ۘ�HD(oA�O���M�ڃ�}1�)u���`#3[9G��{��:8��_;cY�"�V���æ$g�4s)Iͪ)mӻ�t%�c�Ra�Pэ�f@�/�U:`{��;|��XN�V���#�\��ԅ��-��sЯ�
�9�x�����#��y�ӟCY^��������B��h�GCGpD������x��Y�::�P$�ɳc���� �zq��5:H[i���׫�tR��f�Ue�o09�-uS��˿��z9��t�}�n{���� ���	X�=m�=���
)iP�J���T��[�Of��	(�e?,.)�s!SG�3��A�=�w���
fS�lE�щ��y���[W�pGu�V�2r=�G��-�Oş�=_⼒yΉK��ƈ#7%_d��*`��`����+�V�3��:�fk���f���:#��1?F�ڱ�W)o��v����S�ΐ>4;��[Yg�S�&�5[d�g*oH,̡�Zkt���s��+��.�_���O��ܪ�#��ȼ)�a�#��x�l�=�.�s���[l����<��զ���I2_2r����Dވ�*��q;"3��ac;7���,��½Y��R�>��Lk�q< ��I��P(��J<I�$��a�%����K��fMc����ꐿ����D|��ve	zwh/E��Z��� ;�[*��p���D�K����dI�q�hd�|	=,>?�]g�dU5� �[qZ,�hxQל��X���h���"ϴ�>�ɲ-�Z<�oaܺ�	���-\�6�3�y6�_0�c7lw~�;���5�!'Qxؠ]^Й��(ó��]�4�ʱǢ�7�8z�1�N;��0_�J��r���N�!-,�Q�����Z���j�P=/��(��:�0��`7������^p������Y�s�	�X�ħU����6KG�$��y
� �F�?#�PfHE���K�N}���MZ���� j#��E�s �|�E�����j�oØ�t��tf�����/��*.��V��}\:�|}MLXh��(�Lį�Ew��z�W���m]~[�uL�b�K�bx�z��ֶYff+w�d���a11?S��Y�
�ɡ7�:k���S�.w_�9����J��7_�����}�9:�'�����=T<_mH�2���Cf]���}�-ysۑ�jӂ��S8����E��3_�SƇ8��$±ͥ���b$N�ISHH'���|���`�E��з/\��|r���Y��hy��S�~~!f�ڬ�|��㈊e��׳j�y6Y�а��v@�"Y�-��s����B���&6�\q��@���ý��D|� qj.}v�ԡ���Y�r���G"�z�"�h�����,xG�*��6�����[1F7���t�/ɽ̘������ek����%{��&�K�� ė�Cv�I]F�e����G�v�Z��J�ϻ���j0u܊�4(�_g���w�@�{_��=!�d1J�$�9aU[Q��v�3�Hn��ۧ��@+g�����l�,-����%k�`@b�J鯒�B8m<z�d��v�Q��}����ɧ�HƎ�@�5z�Wq�7��u0�h�?�a��'��.���S#}٣n�J�p����=�Au2.����^c[�`oqǩ�*�w�;��ӟ�{�É+�j�F�$TY	*]��i��jDvb�@Ƴ,`���S˂y*�K��
�!�MX�Iet������|�|Phz��Ni ���?��ʞ�k�p�G-?�E V�*�Ӓ��>�U�e^!�=m% G��l�h`%,�4uCǦ��q->2p/#{��o��*�↗���^JQ��b�H�����}tQt)�
pO�"�b����}>��7x	]v�1�7�*ސ1��Q������K~���DhC�G�5��}�m�	D�e(Q��1Cb�(�"��_��b�K�.��A>�p��ߏ�.�L�b���k�PGżd�q�+�ï�?��o�>J��i���qX�)l��M\j�e.	x�?��j�e����Gc�=߭�N��#(K��FZ��Y�ROXX(e�5��5}��'��b�e�뮖g�h��XVmU�ٕ�\��Z� �+�YyyD�
o�L��9Xw³���/J� �U�d�W�|W�qN��ѳ�2�~8��>4��w�^��w�Z�&_EӸ�|㸝�?�=��z���Ȗ�u���f��G����0x�����Yψ��U�����n�vxg0�Ȫ�B������4u��V�1�^!@��$�Y��bX!h,��6�P�To{���!�&��Fg�@+;m�S���Հ��<��]S|�,?гXbK�'խ�������윍Yx�� �'�q2lv@w�Ӓ��bGV`i2��i�!���h��3�y֛�!��W������QC�� �mܺڿ��CIus��� �l��2��P�%��$�̟���ɍy.Zl�&���y�,�/o�N���H�}�[Nf�m�h�j��B�lq?��TfpB��W ���f*�KpEͼ�Z�i�D-�g��F�̄�:��� ���-��}��z�c��o�ٱ?��1���'�=���������5Oa��5�;C0;�t�K��P�j�\$b�xq�F�����;�cKֽb�I0�����L{�N0�r�	l��a7�Ə���bL�V����{\��<F-2�/����G�ﶍ��0O�r���	�f��(��Z�wp6�n��35���Ө_[6r��"uT�iq��W��Zճ���Ϩ*���W�� �WǏ�8پa�ΞPwsu����:Ⱥ���Y,桀'�=���-ƨ؈\{�M���\�^��"J�"�x�W��i���ꁔ�8�O{UL�'��=Ě1\Π�E���x1mD�(�[�K�Z��1�����j�-r��<�޸\�Na�"��71��?���6q���(�y��?!��>�'t�`�v�!7<��#ɮ�?]�2t�V�õ\�Ɋ���jnG~��,)�dI�^�"���3�f��n�����0��)W��8<ߺ��2�`6�:ʢW8+w�ۆ��S������ޞ�r��<�Mp*�^�� �=`ȶAc���.[ ���nN�'g�c�F��kn[X����У���4�Sz&5K�R�^eU��X�?ߋ�yS�B��d�C��0��z�,�{'�{�_ڥ�d-����TΈ{��Π�9�b�(z�(}4n7�n�l�G3J�r���#EwF�$��@kG͓TL��!���Y����d��h���9����Eԯ�ߙ�͋�IUu����5<�2����\2?��Ѱ�`�����_q�ԓ1z�Ϡ��ګ���_������f�R�:��Qzo�S�'<�hv�7�I�@����~�n�|�.j�&�<1R��s��#w ��y{�+���h�@ٲeOXn46L�g���ZU@���N� ��%דs�[G~&:R��fJ\��/r���}��5��vT�j=��X�2���$P}9^ZڣY�˝��ǂnF&E��~�aq��[ � av��UvY�~'|�e�,ջ%���ݧw%Ф(<!�rc�4g�/��t��r"1�1���b+	�|��%6�_@niX�lr�P5���Q��>D6|r�^_��ӑ8�R�"��n��w�ᔏW]i~��ެ"��g�u�y��s�ÂGO[�h:��ŝ	��ǒ�]oZN����9+ZiNcT�E���݊Ŏ�}�߸Z���N�ҏO?>̶�b�	�b�;����b*��4w4�X�Cd/j���
ь5)I�?��z�)>g����VVQ��[d�i献 1��2����&?'��:dwx�LXh����9�ڭ�־��ףa@�M\�Q|�Lw%�[�ײ��J�2�� �#h&����!� ��V4�t�dn����l�DM(ݿ?T�R���o$�a���GI���EhF�+�ؤ�%�ጀ�A���;)B,:�� @�1�ogq,!��=j�K��]�wo݆D3u!�(��,{��{o GV�!�,6k8�d�*�$���
�G|�}o}�D�y��שּׁ����ޯ�����zU��en+kkUC�[/�}��=�O/U���x'�N������ц�޹\���##$���m`�/��t᳠hEQ�UHW0�������

�r�O�}቟�v��-,#�:�wD��4���{����n����IjP�F�l<��S��/���
���⡪�ުE��/ƈ%7t�`J/&E��cη���j�v�j��;� 2��K��bA<���>?���*�ɯ4����>Z��S̆I��)Gw��zfD�U����vB�ݸ�q#�n��E����lj�B���4n(� �\�=�ݥ��NgIv=%�>�eh�W���N_-�z��D��ל8`ܳ�u;����4�'-��U��Kk��tҨ�2�L���sj�̄;A��/��;�����[�aO%u=Z�⬻�u�Ę�'��<e�a���{`�|�&���TE/�>� �8 ó���hK�Z�..<�6 y�/�����W�NSXuo>��-����a��H�v��㹝\�Xۃ}b�cd Y�	�\��4���[)���W3?�<�!	���1��T	��F�G�!�'Z¨���bUyW���W�Q��$GF�Q��A�'�=_�;�r��,L�wN����2s���$ߝ�I�Zzl�Z��X3yI������_k�Ҁ��S��k�ޫJt�0���RR^��%A���DME��"oc˴qr��K���#������_~�mN>�:�GC���)��(%��A�`�����n"]Hf"< ]�~�S���-0]��#4��ӳ��-��A�Yh��6��S�{|j �%�Z���o��X��׊'�8��#EtG�1e��g7E6�aR�d+b�o��l5vH&�Yw��v/�h��5����T�^·��!����xh��LXB9ś���{̩qfR����E4^�%Άy��Z�w��%M��Gf�w�i;]�Ҽ��f7 S�-f5�hs��%���槄��p7��{z���.�(�Ӣ�U����I�|Bk�h�����;������K7[ߤ��+RB�����)�]��&�0�pB�����%�~ ��Ó��!)YyV��`�FpJ7|h�}5}�4B#�8E6��iы~e��e�v6=KMI�	U��6���9;��C�)�|�H�xX�UH��wm�,a�����L�w�e6�QB���F�H�1�g�|	N�S_Q4�7�8i�8�[�/dB)�L������h��Y�e#y�*imF�s��,;��Y���G�#B��Z|�_�.�Z���� &�L�5�y0�}�9/�'!c �[9]��h��>LQ>&;`�-�~~�������'k)ܬڀ��q�ϐzu!Ì���qJ�I9�n��b�����, V�C��󑖢�O���g2���j'�xzg�����bp"P�T$߂�r�Ш?��v��O�U�u�!���}�yKamJ��K��E��`D��ū�psI밧#F�Y�Z������,�r����޵g|��UlS[���>���<J	�:=e�"��&<�[��)e�8���`�]��xq����|�rN-)��4��xT(�4
�&'�kj$ y�����Y�$�g<����2��3%�n����9ϰRY*SX�Qo�2ѹ��c􎓊�9��@ya�qc�̡5	�c�a��aǕ��*��3�OV���{���+�yP�}[�"lx�7Fy0�me�p�9#K�A�%mhCA�a����u�ny��S%�>�7��3�X�0���t����{p\�������H�Փ������搰^�(�[�M0_������A���&��Q����x��׌!���&�6���Sg��bR���6����`�ָ��Z����:�ڒ�C�S����T�t��zN���D������x�N/H:�:�q�2�L��|�y�p��c0�����
�g��������ހ��i;�,��\4K ��W�;����5�JZ�c�[�魷|l@��M�fL�-�!O�`��T _]��������Su�9�n�<�r���`Ϩ[ɂ�D���p��?����y�D���=l,I��:gAҤܻ��U�a��tP�����A��я������l ���p���<��#
~�z`��5�u����æ�D�҄�D����Y�B���'���	@�l��|������Xd�|��t�B�~c�₨�9�5���F����I:c�P�b�P&��-@�\T�h��/g��c�{+����M�BoW��p;�����"�a��32���������&�2�Z4�WXT�>P^w��R�Ehd���KM	�.���c�����c�u�x��,˶�g��0�2�)�2"�E-���>"x$B`�J����6ǡ����|��"�矟A�ͷ�hÌ ���
����![�Cwi�S��AQ�V�ҩF/@LW[j���CM�Y��|#��@��`���ڵq��^^M4۪�ܜ�P�R���F�է�|Nɝ!����"�ۦ�t}=�ɉ����$v��/Ԃ%��xP���ѳ�0J4i������s��ʵ#��?TŲ�"g����ʾ������%W:���n���]����d���)�aL8�RM�gm��es�O��	��qj-���6��QD�Y��2��C�T����\/�6���������{I�ɔAt�vZm{,���P���"
Z2LJ,d�|����[<��
E�i��#;	���c�ʕ��+ե�I�-%�;�_�R�M+�h����`#�V{�D�O�S������j723dSu�" ���4n�(o�@	���m����(#у��Vozx�^N,J�w.�66�k����>NF�MT*tCv�ř�ӡ7d���N��O��F������M��'W����25�K2p��j½���o�>F钙�����T��WWx��O�������Y��ƈT�AQ!�Mk*������&���ǵk<V�K���sY�~e�<�)�Ց� �nYi�f�f�׾N9�j81i�ZS^Z��	�+���Zn�	L��,�J?�e�"��ڕ]m�݊D��Vua�c,'ʧ:��қ��@�ӭ��S�S5��&v�A�u������#<$Q�U�,����=Z�����������!rxGj��[�'f�M�	iq�7! 5\�f=�)[���d�����7���OG�ȣW����(���7Jg��[�$\%^D�dZm2�zR=c�k��*S5�o��#B�c{���'�A��ED#K�g�Ctז�K�]`����)�cUf�������،�2{O�.-VwUz!v�19Ǌ������	T�/�Wn�������=r��A�_�@�հ����E+3o�4��|+Fsk���%����`q��1x��9@z�=W��U:���gy~%��[s ���]F&|��sRx��/��sN��/�d�hzJIxt垀ҍ��1��X����٧�6�t��)��\�b��/�?�p��a��M.a�N�Ű��n����C�AaƟ������@�1�cw*��1[7���ZѨ��k�A�*[aj��?P�z�VQK.���cM�{�3�]!-�*d �m㍭%�5>�o�'�v�Ċ����Cm��n����䯗V:�Ȓ]P|���-H�ܜ&��Q����L�LZ��� ��8	 ���HP�V���\�V�}�G���5�j�X�&�/9^\o���t����~�x|=B&�a(R���p~���g��z����+��|+Z��*^�<F�L�eU�"T`�V����F�r��}Z���ʽ�W��*0�*�B�{ ����b�V�v�Lz=e�	^��h{.�W}w̧�WM	� xj~ʗ�j����0��	/��a��`��a��Uެ���I�4=�I�d^��u���ʶY�l��@I,=����k�����#���Fkc�J����/�$�8��yI���_��+��q�d����F�v�(��~t:�N?�j�����'�0�57`������M'D΍� _{���}Dq�c�>�� �䱄����~���J�f9�7�'孭J�X?,謝m�"��B�j�?����9)��A�U�ǅ�6{�w�{c�t��}�<@ű��V�E�0��h��T�b7��e�A��!ςG�z�'mV����D�;5���2;u�&�� �*�����[��l��?=�I�-���(��PBg$&vL�۵�"w��YO���D��͵�VL���%u�@��Ee��W�~�����A���C�ʵ�a���@!x���ИH�6���E�dt>N�������p<����#��%@,8{�|K�efF�g�Ӷ�x��٣���a��&���CZc�:�G�<�O��a�%©ƚ�:dz�%��n\4#�߼?��^0O�u��a��E�{��"�jq��Z���;o�K����k�RNh.q��eqx���n��������G�xf���$�#:���]�В0G���(�d(sl�=p���?������������ܫ���t
��7�,�:��Q��ı��w��D�������P�Dn0_��:y���p�'@�1���o{�vGLBN��. �p�xb��%��߇��u�D+up~�/��;ׁ$��Ɋ�yc!�H�C�
�m}W���/���zd
/�`#�'qi�c~\�01��<>!0'*Z��
�qt�~$�j�;�Ȫ���_Vl�����;�Y�4//s��	�3|���_6���HL�;�ħA���Ç�ّe�(��o��� �-�*�~�����On�v���U3��=�:��Ϭz����N���A9�5[�����\2�m۳����%>F�]�O8}���F��m�Gw^���mr}��>���y�������H �n�}j B���3e���|�-C�4?��]�eg�L m^.-c �!vdP�T����U��v�J]��Os�nm�+��2����mtخ��-���gpl���+�j���Ɔ׈^�sb{%lR:9,9���Di�-�X�%+���͙��{r~�0_G����:7��ܻ�'|+ �x��"
j�s�{�݁}<5�g�!�A[A/�r�O��STcqP1P�!d�K���H�؅�n�ZZnD�%�]Pw���Y��CX��������hF�,Z`u�
���#�����D��z0�dF�.��&n�3����]x*6m���:�����!��g&Z���p[�� v�q��?��������(Y��Ԃ+�WA�I�a�����O�C|���`ձ��������{G
)�f�d��)�&k�T3A/��O FD�_j?fl����QX�͝7vR�/7����@)���s�V�˞��XRғ�݃���*���n=bP<Ʈ��X�˜�7 9n�a���Hu2�>�+���@R҈�[?%>��5&'�0����vP�G�ݖ�{�X��g�++ ��A�Z�"ɠ����+���A��ҡ5� �8ɿʁ�\�BZ�Q�v v������ߵ��/�4P��{�>͸�}W�T8h��t�Y��r��5�i�J��_�Ę��[��Лؖ�0�8S�`;�ע\5 i��8&K�i:q�n}��#�jS����?�K/��:	S#-Z!37�bj�n*�C��)���5����c�ja���{�9�ԡU�����zv�阪j��?�%�$��9՜�4?�6���a�i:C�K&U�x�Fs'P��<K�ʘ�"���=�f#�QEd�S�-�k�YR��s��e^� =g�j�{�aL�n���P���@�=���Ƕ0�І>�Z/���	g�/J\)���k9�w;�Fr�	_G,��Vgu�]�u"�Y�M��)��Ng�@s��&�6|�S���A����D!�C�q{
�铘�T�u�	���so5�b?��I�:�y�RӨ>76H�T�\P"OSZ���h`�p��.�K��w���]K��}�A�`���x.7�<�d-θ�|�F�1f�%T���q��W�yx�	'�؎���?�+̬=��P��2C�D	�(c��TQ�����!b�Q�ؒC����q�hy�u¿�*������d�����Ts�;D����/��i+S��G�>�PH�@M��݌l�d�P#�)Fڔ��f��q�D�����΢�R5|oF gR�o�r�(f��
�6��G��N�h�N��d��n�I����\���f]�b�Q����~X�-(V��z|:"���s�h���qvZ��+�WN�͊���g���Le��i�	�{撨|Fn�~�Z���D�'���x��!��L�� �dn	�"c!eL��q�i��m��<�oi5W���HU�q_Eq3�BSYtm�XA(q)�K���Ś#;7���}�#�&�(��ԝ�M��81���{���p�#qk�僝S��s�ãNf&��泲��� BP�!���Z43�c��x��F<���rM�n�$��z�B��}�ħ{ ��ֵ�Je=�h�����~�>;��z��3�Y����Kde�>��:��A�%�.����r��CjK�0m�>U�{MʤB�nF���_�n��3�ZBiL��+�"�!�C2|Fw���Ϥ8���יO67d��JV��]�M��l̃��t��i��6��)��aܕ1�rP<*T�ci튙��A)�:�	��߯ae��T��wѤ�9ֹJ *T��떄���	*�V�S�� ϣ�ÇP	[��j����$G��l�)�[��?/�\�(��m4��e�8��(k���� �=K�I��u�F���.O�UJ\��jo��	H�i��i��$�9C��w��b�e#�E\˜����Z�X�p �M�kۈp�T[G��I��c�f;dS�Db��c�&�k�jm�A�#�����ũCumu粳h�-w�ƠEҶM�?��D�z� �-�2��,?p�p�s��P�Pwɦo���{��ی�ff�a�Z70��5SJ����t��|%�GS��&�����������B3as�/0]2��y���N�w��>��q��D
3h*6�f5�F�Xuc._���_��#I�w��5>����eO���%�gY�)�!�t�����Q�GW7��.҉�� ��a��)�0::"�)�����#�g�K��*��-����4?�~/7(¨#��"��n�� �%�v6̻�������B4�+�(��>X��q ݘ���_��z-�4��np���ZFW֚q��\f�R�4J;3�*��ⰴ?x��i�G1��� U{�Xz��&���1{v�����n��R�3Wq���5]3��XT��:�z�����2�!�jx�v�w�B��u7=��ļڌ�V�#���X���j Rn~�E�r,/�H �tCL�[��F���������o8~ �]\F@���f���X�"�gQ�_o���R	��Eiu��Z�y����"��?����BD�,�Kd�N��cϬ�C��8l�l>�"u#q�ŏ3Is�^C���O��̐bs�+�j�k�{S+R,���Ƕܳ�
o���Nk1݋="���\��r���8��=y�PP3���\�B�!�[$�51G^���Bmf�+Cϒ>��|EK������Np��b�[�c4�s�@"n�W��SD$���u�[�ٝ&9�T�/[Q�\���k�uQ7�.�l��b��E��T[ݼd����$3�]xj���z�`�� ��.1�L���2m��q��4Z�������F���Q��H�Y?�o��7�쥜ë�d�ъ�-|zw"sL�ph�b�@d(�nt���3ps셆�g�����^����Vq��O=H��(�)o�]�LB�#�0���xU����1��y�%�Y�5H�H��C�9�f4݋Y*P��p I��F)D�.ja�����g�'jɉ�Ød҈����n���t`2X����qΐ&A��I @d
�0)�)��|ʢ����_�vXl	!�^�r�+��7͛�$�M�_+��p8Ϛ�0�-�êiy��:��@Gs{����I5�J8�����uÇ4�e+�R����Y�߽�z��3�tm��.�]ea��G�(�C�hFǼ��!J�>�0�BȢ=|�,��L�q��������`�Е���D)�kz�����i�Ws������}+�ec�SRezL"�x�-�Y�x�Y���K
j��ux�>�G/���|�8���՛�ԁ'�"@0�(�f��������i�C��^�z��&���3��D}�$[F��N_�Q6�g�Hi���2izmq*Ź�����H�сF%��N��u�<��Y�S�S|�L��ZB<o���92�v��?����!�/��s!���w�Iw3��*���Ze�~�я���2���4�Ēg�8�*Q����j{S���7>U�}�˶4��bUU���6 �f%���Y�FA>�
��P��-��Zz�l�4��F��ˎO/xLڢ�I�t�������%�*\�X!�翆^_Z���\C�M�M�|)zͦ�h�/�ˎ�,r�x�rm��#���n��"4��N���:z��8S�JU[��C�����W A܎'I�3��
���pٺtI@����. ��S�iE�i� ���B��q js�n+��� �����+���_\ �x�_j�G���O�kbs�.Z~li�c�x�C��D`��c�#z_ӌ�86n��?����@��_X��l��>ڀ����7WN�����tx<g-H��f��a�j����\ �a%�N�&v[�1M�<r
u K���rcA}f��:��&�'���'�}��aA����1IJ9՟�fս��\ g���p
<F�҃ԝ�Rj���*B5��Y�[,3�Dn8t�2L%�k�_��~����ޙj���!d�kŊ6.�|~^���Z��D�CŚEЇ�ң8c��:�}1N븣(��SeE�P��?��HeI�sl��L�G����s`��0~�&�J��g�"��eGafW0�^���'�f��zo�8+/���xca�ۻ�et�*�I]74�xz>,M�����d��������1k�2�p�(4I�n.�/F̦��,&�:�0�K���UB�Fԭ_R ����3�y#�>��޴_s��ɔ�AE�V��ԉ7��=X-!r����>@w�>mQa
Z/Vg5����^,��~ٹ���d�R�D�b򪉻J���/�V�[�����,�]���)�pU���O3�]ۡJN���+�^�'�_���k�=HK�<�o<?��ۥ����ɯI_ul��WF�Ȝ�b\�E<�m�Ƽ�l��N�>���;M�\%�"��Ȥ�Ԍ���3��
�4�0�Q��&\�]F��1�?�m�5%BzDM�NW�u���C�����D��w����K��'� ��L ��EJ�����P��p��q��>��\�I���0�~m0�F�8�N�|*�\Q�ІG�����$�Ѥ��@AJr������̶�*vS�9짤͗��M_o���Y��Uu���;�򑗃~��2H�w�J�89_�Xc7���ZTK�˻��]���B��_��^c���D+��5d1�c3͏�s|i����ݘb5�&#���1u�XH�)�.��%�#��f��X��v�:((��>ӂC�w���{Z����戡n�.BFCO}*������@c�!�v)�����<�~~q�7�%�N�;|̓�ڱ(�&�{ҪS����Ww�,:��?�㉿��	�C������`$�ӕ��<b�&��{E`�Bg�)"�g�z�R<�+��Qo���+K8r�bF�\����
�&ޥ�E� Ҁa��l _���>���9�1�}�GZ���lW�*�j�y��j�+��1�%�)3U@��Tq�$�Ё��1�hʯ'�D�v`o_M�O���������|�$�5��X#<s�c��v���!��?z7�(g�[OQ�9����֪LW
�m�/N�S�����������b��l�h��qU����YKu��`X��6Y"��w$b�d�\��1�1����4-�(\y��Reh�Xy(&5W[CN �Iz�pѶ�Un�
���tط���7�x���s��ϓ�S|�#�P�U~��Zf�'뾱� O!-��,]h�����ɥ����+�.��#�;^5��לN>���}ۡ��A�L!�щw)>C�g����#*J��Ё񨰢���k��fcqʀN��!ۺ�.���d�u�q}�H�1�0�+0'��{@۩�)Z�B6V�,�ǈ=�N~ndh;a�.1���}���8�z��NR�~g�/p!(�r ӯ -�۫���"���W���,&-+�s<<@��2�袖���xŇ���v\P����bװ@�i�l��1�F?6C�3wX���3��Md�_y�u�2b%�J�%�	�v����Ǐ
�M�Q�(%�e��Q/pL��|������"M��X�DX�ګ�V�p���k�m����qV�o{��ğ�2���'�m a�	�_)a
�/X�l�W��_Eڛ�R�r�8͗�M���p#r��_�Zw�q�_����Y��6up]aH,2��.D2LLќ,-딱)�s��Te���؜�?!��|
����]^!�/r O��| ��B��JD{��%Y�f�njA����T-L�����RC�� W�� @�U��T�����v7K<���G$�&p}y���sٔ��_���i\1������vJ�p�
L�=7g=��{c�L��K�O�"�����èq�+�����V={xs�q�
x!=iq��	�ۦN�«"�]�. h�i}3�z%f�?��R<�U_�U��/�['�����w�.�QX�-�?؜u�SHU=M�����q.�:���-7zg=K$*N�vdlG�Ou�"1D$�[p��0F���u�3,"a}29���5�Ҽt����E�84��*�����ϋMȶJ3e���pҳ�y+�[l�w��K�!�Q�CPH�Qw��+q_0����^@m\}y5�	�O��03���Cb����c�O���X�ٽx��bTo���&��>O����p?*W��r����g�r}�̳H�X�u�J��Gu�_�����-���eRX��,J�,^�H��q}M�:�}�eB8H�/�G�%���MՂ�햦�+�B�+�6�>Ol����OA;�F�e�ZÖ�MW��M!.�ng�G0 %֏�4>R�,�3����\U�d��������i��Tc�;5l�Z������Sss��kISyo��R*@>^n-����]�۹,@��y�٭,�
� ����Z��4\�1\f����2A�֐�Ƹޒ��UI��VԀ��u�Nnk�mF�b"r�l����d���	�_��|��r��YD�I��M�8�1Ep.����g���;���py��9��#o���x�[���P	x��	��7�(lS||�]U�#d�
�S~s�1[�0��J�Ah��{��2��:�D�S���Ꜫ[�󬍷K�m�NX��_���ޡlK�r��񸣰H��\%bn4���~���r���}���)H��#���Pfie�aDƳe[\IH���x�9`��0e=���Uұ=��'�.��� ��Ԭ�X���<*R��qy��I��1$ΟRx8�(�XM �4��q}Y���n���p�O���b��+限;������	�֖����&0�a.�N;!����~��Qo�n�T�	�К�o����A�N�Vg���D����frk �sH�	zU�zX�T9�Iw�Q�� uu�'Y�JsmjN�pl�� �ZIk�|��V em
@������X�I����8��&� p�BߡiX��v��r��9�y�����ف$�e+JJ��\���=�;�靁V@�;�R�'ӡvhA�U�K, ���2�	�Z�p}��������2);�L}�\���}�+*{�Ժ��$�_.yU�D5��5b�ܺD��R�TY�̀���̩���.jroX���P�X�>��+�$���Ǫb��� �`�$�喔2%���6=�2�!��3� G�>��V
��ȍ����_P�K�Sq��i�8����̎Qn�A�xK���PH��C�A u�3x"LRȖ��� i�׋���p fd��+��73,f�mw�ۻ;�֘�FH#���a��ŵ�6��[�k�UL^Q��ܾ��������.+��Z����V�;�����J�щ���e^�긇����u���߹4}��b*������)j��>�G��OX��g8��TK=:Aʍ��ZZ�^��;�i"��)�n��u�v���=w~�	8�"���0��J5� ��uP=+�f]���Mj�Yd-����&T�"�wE6L])��aS��f�/���PXw�Y����؂`�-��ˌ���vk���D*huǳ�����GEI4��IhZhEy�kX(�:J�Z�q�}͓�e��&ַF�T�Z�j%�v�ҧ�����v>�6��4���qRc��K1����h�?�����8�9SQ:h�c�����.(�;�u|x���Q|j��#�4Ւ�h������^�^��J�D��/j+�*���S�(��R���kRd5]�&��5UM�8�Yѵ����u��3(zO�$�ކ2������k
p��h�6�@f��d) $h��q��������� �����U�� 9�7�$H<]%���$g�E�7Q4b��A�|o���5���\h�Hjt�0��jZ�.�@o�P��ȳ���`E�����G��,ӥ�n�e�h��<D)�h����l�^<~�P\/[}wB�Ҝ|��l��J��C��0�
q�O�َƂ�}c��C�@�����&ŵ���>vFB�I##`"l��w�����m���[�tP^r�$[O!�j�+)�OF���Rv������aE"[�Io���n�C��v���z��E�f� MP�������e^�眸r*s�����w�l��v�k�󜞥e�c�����p8�>��I�5f��f8�?�������6��2ȥ^��������C>�$�=��6��|��N�L���B���YdzLhV~�Ԫ�#�C� ���[ �gE�o���"CZ���l�ںH�B��Wv�j�����۰�.��:U��A��1p��1�r�b�V>Cf�C��2ゝ��/a򅲞�����X��&�{�nf�ߏ��f(��⌬D>�u��]�mn9�ʡ
��eVu�D5��?m,�>
���aX)���r�(7���	Kk,��<�_N��vsr�9�q��X� �{Q��N<@z��LFYA���ׯu���I�t� J@R���mvMP��#���0<2~g���Ͷ#����ݯ���"V�'��B2�X1����F�,��4R`���J�98z	�̫b{;F`�d�/����9̶�[�1������h�jҾ�z>���W�Cnl�=���=}�mB� ��k���mB��R�V�I��f攟�*@&5�iI��^͕v�c?�-I"�$7� �(N�`H2B.:Q�d�Ž4,���Џ���Hh��7/5˨%�@þ�������u{�O����|��*�F"��MzSe2��15Z�H�ԀQ*_�TF���. RӴ����~�M�ʜҰ2��|c�(7�:4���n��=�1���;}^���2�|�C�]�"#"�L�;��\�'�C� ,���f�ģU��:��uD4�0�c��|P|t�A^w�0���6�-�#��K�39,X�'(��ir��m�7ᷩ�u ��ܳh���?�@��E,��5L�8	�.d��P�}U��½��Їj�0Z����ծ������s����.��FvuӠ�0�e 1q~z�]�'�B� {A�ر�k�mip_����-��z��M��e�%D)XY{zOl�0���sEř���Q�ȅ��������A*X�0��L�~�⿁P�!H**eY����}{�!�l��I��&���N�d~`$UK?�Ϡ �˶�>�ʂ�Y;��rH�/f7�u,b�z��]���r�7Z�	�x��&�aEzU�Y�5rl@����R�W#���df�!�$	���RW��[��$��eb5�|���1�W�T���-�đTw~�r���4�K���d��#���{�#���1r^�Ӿ��-jB)�f��G�fO���Mͼa��r5ߥ:�J��d�&d_�x�Yt�G��:g۪:����t<�R:� _�}�]_��{@"�8���bcȬ	*�5������n�g�s��F��ٵ����4���	F~��ڢ<6�=���~mx�6�~c���ޛ��}Γ8K��btB&�x�sJۼ�H34�y�&X��L0!�b�����<�xV�p5b�p?�I��{��5���T&۱�4�B�P��Qjd��{3�*��ȣc��~�=�����f�2��9m�.ƞ&�hG}�Q��!���.��mFJy<x���on���ˈ��q�l�Gb�����p��)xIIWW@�.��J���A����v�Q?
�u䡡)|`����}���QY2R]R�<����9 �u�X
����-8Ƿ�סG��p��U�JR�O��q�on�'V��k�nǡ��*�8P��;{!o����SNi���jl�~�_Ç��Z���
�zW�Y�D�"������k���m�qO�ʬuq��QC�����t��T��
{��MZ�T��	�&�7H���?���K����O��>Y�DNЦD������Ϳ*^+���*�_���)-����T�x����.A~ˀs�F��<t͊��,͉ȏt�#c�Q��.ڕ�
�"� Ft����h�:j�R����$��x��21��A�C!	18;Ih?���c�#�S�廥�CU���t��JS����^��1wn	��oT|���������x�
����D��`���dj�6��?�6>�.m�J�!RJD
$����O�Mu�Vfl�Rxk������>z蘠�-<2�`����{Fc�%]��pAcu�*�(j.�ipӯ|:o=����D�xMx�e+�M�U�N&k��ڽw�ᙽj(�-��k߳��c�e������_*C��(Ȓ�d�nF��c�kS��[|�@nS��ш=B���D��� ��(���v58�x�H\�1�ݎ��m�5T��;l���c=|�9r�	�1�@e���b�����4c�L<C��,Je���� ԉ��E�M� �5^Tu*�*�G?�vO�������Ÿ4N��A��CU?TaiD������w��v����u��.H�{��Xl`�.��k���3�ҷB�V���@�#Ve�	8�}��.\��vp�i�!~�s�Zj>8�4\���n��LI+۸�*��P��	R����D��g�������N5C��J�V����S�*���ڐ����7x0�,���j����A��J��y��Կ���8�Kt��	�x��ψм�ZKztN��h<[����{�,EK�Y_-[��8����l~����`���=��v���npD\���U�����K��ȼ&o�EO��5I�2A�V��w�P�N������Nx�^_��p6Ó�i��2x;e܏6��.�~L�=k�#/ry��6��8x�P� �Ը1PΝ��z�\͉����u��!�$X�ӿU<6�L�d�t�4�T�]^ _ɋ!W��ݣ�-ŻE֠�0��5�~��p�Ͳ������P&��>B��O���L
�B���* ��l"Ux�����1���S$�ma���nL��T�ng⺘U�i�B6�dC�=&R-�炈����E��w�����A�B��)�X��>�x�����M6�n�p�
͵�|�ۦp��d�e�Hh�6�w׍��7&�ЃSX��L},R��zx��k���U���´�h�/Pn�iJ��X�Z+��c�n�K��(F���㾗�Uc�s	!�S�"`y��r�|����ݼ�9���i��#�|.R�sЋv� ��l�5u��dO"D�,c� ���GL�t)}N��?����0���p6�E��4p���}�-�+�U(�y���´������'�6�s�i�{@�u�� X���i �N�2i�چn�2�g�f�:<�ɂn:�����?��#��×G�Eq�mN�bgD���ӠSIdq頉��@�XV�E�"�C12�I�S�k�5}�W���SC�a�%4�zi���Nk:K�t�Pv!*e�$�O����w��}�`B�!%�G�j>FE[����Hx���vcIO)�4 (f���m����d}�U�}@=�i3��UNv�����W���{��&�)=��RG��~ Wx�����o�rC��� {XEe�>�ٛ{�(��tt��ɮ�X$/^� Yꗯ5[5���i��k$��_�P�D��w��k?+%��F�}�ֹ�x����ALʀ!�)��ܾ��k��C	��7AI�̆��Sh	3d2B9rO�.a �M�Xۂ�G[�C^�2��8W^��~��ݠ���Uf��?6�+��2	��������
�/�����2��(����?��\�S0�x���mEҐΛ�йX��@�fDhQ#�&�s�E�_����u�P%lh�mHi&v��yƜ��$s[��)���Q�9o;{��<�����_'�|K,J�2�/=��%�PkOy�1�5����ڝ�M�<�qo>���BsW���7�h5-MO_���f���5�r#h����~�*�/
6x	��{�su�ٮ�����s�l3�Ҷ�'C��4J�C���A��!vT|�$�ǁ�W�rɁ���]25ƍ��Z�X��Pڦ�^Ns�gS�_�%)�~�w�
�1S�O�\j�)�8dx/��9�!V�Pl�
�ܽv����+��J9A|O>})ȴ0���*��i�(8����M-����s��:0r��C�ƽ��>:W�$�W΀e�����ȑ���R���GP*Y!����#���a��`�ƅ�'����x��6���_�|�;������(���j��
�g��Nc����g�`�`M��Q����=�V�����?�mr+̪��!��(��g�2�Ź�N�aL�,���_i�!���������*�g��6���H�%���K�g���]x�|����Z�\6��CP����qY7��U

����S瓢Y,�4�+���m����2���w`���E�� ��o?��(O~�p�ofaA>�f츉8���P�N�S`f ����$��.���
��m�xZ�m�z��O=��m<��4��<�{m��=|��s$D��P���X�u����k�/F�z��譅�?|�<�n<�R�~�%�]�|Y�2A�H�����1X��k��>L��.���jE�M_�b>�<��t�ً�g�\9u+�!>�"#a��"�O 0��U�x������<��`��w�x����^N܌�w�`�V�����җX��p����`ys�&X��)'(ox�~w����F|�#������-�Y��Dξ�o?�kG��d�\H�@:\#x�V����K�n�U�?7Q���`ͧ��kPI0YZ��O]��i���W����4F�DQ? <�:�͵2�l}O�0�鷏r� DNn�H�c3Lu�\o[�WV��9�Q(H�dTg���y��:A&��2\��9����V����ӖU��?�`�#��e4�W.2䎙���(a% �h2{�G)'�*j���.t7I�95���k�2�z�T��0"��n�̻�����6��;˟9���}TC^r���￝����?E:л���$���D��ȁ/!0/+��13
�Δg4�*����n����ԿۅY��l$kp/�f2��+�qpQ�?�p����ʚ8GF �x::�+ޟ��(�W8.����,o]�I,���W���j̄��q�T������:_E�8�!7۪���Nĝ�|Q/��.�+Pj��[Ɔttˡ��-�sw#i����}/�Β��;vD�Մ���;��x��@ˁ�g]�~�p��G]q/=ݡ៟���X��,>���(��[z\Qۀgr�Z�w*��vH�1�'r�-�����^VJ�b�0��~�Q�rݎ��г(dD�{��?��[4�,3��X��5���ͺ����� Uwm���!N,m�w��*P�]�p9���e�:����B�1�Z������?#�n�9���D��a[�)F��9����Ũ�hm�0ȉ�� ��b'XQ� eL+A��ϺF<
�Е��D���%K� �V�h�F�~�7�Ɍ���)��{��1xIL��[����l��f���$$ఫ�v^�����Z��X�|H�YG�;M�w��\[��K�,����.y��[��SR��>���EZ����9|;]�ۛY�nc��*�����r�ô�5�}ও �K,��6�\���_q�4�Vf�uH;*5�Et{k��v��]�n�o��
��:��J��!��p���(��TId�y12}l�T�*�#�h��Yjm���	�u-̗��%TF���A;	�6]�0���x��7�u��xaEn��%���?o�s9�t��Y�)��9�y�}+�뻨N�1'�;���f�ݠ(� xk�7�s�`+9J�%IќMpə�`���Bq�cr^�f0���ߗ>)�k2�Ԃե�#�[���i�	3&6.g:���A��7;�ϰu6L�2|�� 8-o���;��׺x���]���T��[�����nZ��3?�~!u�@	�z�|��و\ĴaF�vT���u��	y^�EJ4
�J|4ǫ�0��!�l�@CZ�����3�Y5f�Ǯ?C}�+�l�^4T��;M�T��
ir�.L��LM,uva*��Θ��������5썚0�U�H�.�aw�6�+u����sY@�(���S��4�fQh���Cy"�[�uB:&�n�bu�|��$t��H�Cf��ѯ)M��ڦ�
���ϟH`�<���?��"�EQ��?���z���u��ve�'����lh��N?�;��1��p=Ǯ?�dY�G}�� �/n�-04�[�6����u����-bt�]�*��a�!DT���t�5r���<ƨ!�'D�1��J�¯� �P��!�="Zr#�@�^bL���q����p�{HyG�3�/n�3�Ox
lYy�@^l��lr��¸r��(z{\��KUJ�Y�� ޓ���79�db�v�����M��}�V�[/�k}�������q�{�p����e�j(�T������EkqI�>M��<���
V6�_�\�O���:$��G�/�V�sU收�8k�<K<��G�^� a���xj�AOf#J�wF2���*��j��#��IW^}���`\�,�.ۗ}H����
4Ձ�,��e�4u�^�%�ǩ�m��Xl�����C^�p;1U$�!A-�?unԎ���� ����	���r���'d��m\�C'"bN��$���^~W�ZQ{���x ��ڟe��{*(^ô�3WSK����\�T[����e�0�,1�è�)�Zj�@�`�~k0 BxC�d�����4k_1����q9� ����6(�J¯�i���MN��Xr�%��r,����J!�/���!�j��]�
� ���Ŀ�t�f���HZ�0���\L6�ǐ*�V� �1J��)�V�>��sX?S����n(�����ɦ����wJ����p�q�|tc#���B�-�>�W8/$�+�������\5F��^�N�M�Z��-��wK����d�������I%��Z|���iO-�c�G�݄e���#>d)�����,�Y�:���=�O�C����^��:1Y6r1�'�8q��vt#����/!J��j���FL�K9����k-���5JI-�����r0�V��}F������h��՚��Xyt]\z���GK"fn��4��`�O��rfz�p��Y:�h���|֟5���0Ԓ�����(�,���H�����w���L�a�I|��w��)|��>$0H�ꙣa��H���N6,����<z_O����0i��pZӹ��EE"����Z���i8oRP�e���?ʗ�(wC�_Q�}:�����:j(gI1ʯ-4��R`ʿ8r��m�}�v���ǹ>hf�,	"OR}������~���FX$�<t��>@U��'b!F`z�����IW�
ҡw�ޟ匣��7��j�¡5�<p?p��6�d�R��<ɤ���I�R� ��0�3��.5�Z�gs|t�ة�];���� �Iu�G�Vr�AA���s%����Y�>:���Df�&�Df�����ݲ���)���@�tE��Q��W�D~OAE��W�YE��i�����g�kQ0y{K2���;pO&_g�	9D�����C�P0~�D���<xn����*|�oطD�®��ht}�P2�����3�o�w +�2�$����ʲ�`VF�*>�7t˷�3ir�3릛CZ7&��~�T�_`�(�&��jAγ�_ÂRTw��2�}� )��I��iL4(���!�Q��W�J��R��v��M�S�D6f0��⇆�o9��5�ᘅ�djT��g��%�[+v83��IZ#��Ud�p�U*$��|�����Ơɣk��u�*�!�5c��+�����m��[�:C�HF�˞�u�˱�7υ��{<s�2��͉����P?J���C5Hwι��$�z�`Ku�����u|���ZBnAJ_���tK���I�?$6�]��j0uI��2o�+X5~�!<)�yāokaXE\�-��������|�NUx Z8u%я�K��C��m�=}�y���o�q�` ��R�,� L:�}��:4��i�`������*֑�|'o%�>�$���G�I���'�D������c[A�8�ۇ|	�Z+��Q�	ep;������ES����AY4��������<%�.T^5D�ޠ��}��9���g�Nx���?\��ʂj����9pĕ�uT����W���K�#j�O�/c�[���v��d�݈��Zr�R]
T�����ǁ-M��P�� �c>� 2K���8Z���OG�}kV� �ο̢�#�UX ��ϊ����yi���[6d�Uϖ�(�����«,m��][���u��ڷb�F J$j�v��  �vW)��j���_v��>JzD7
vg:�L7nh�Ü���TY���ٳ��߳Z�xv�\>R\�Q,�p���`�RV�F�M��)^�G(��[�x��o�ئ���sQ�j��a�Tz�8}X�4�����|MF��{���,V%h{F��p���0�7�	�3sH+p2J��J�v٫����J�������N.�'�:]X�r���Xs��|��M����&���਴��=br�Sh閘���'�o;����\6f �*���8K��{��އ¼GӐ��QAV���Z�W̸�kx}Z�'��[g��;7����k^����mo��K1�V�:�@N��U�j%R�F��L.oGe���;ΊC��<����\V���k��5������dݐ�	Ӕ4;�'{�s�r{
�L���>��0#�
� �p*{��#;�N���朵���a2l[�_l?{.��7��?���>�f����ܸ���O\0�m?��6��_���͎n�sE-� ^�엱o\�KU��(�6�8��Gk�D���ͳP�&�t�s.�UA�_�[�3��	|���؈��F$LqG80ӆj���J��}/��q"�j���ty>+�O�W�Qx�%��Dx0�
+�Sg! �;>�������׬݅jlR�gjP��ɇRH}u�`{&��p0��,����� X�i̡�-��v��j���5;�'B�r}�xG�ݐ@�Ŀ:ҍ�ظ��H76�7F׉��s�1�ş�	3��f�+���W0�AN82$�#GEa��z��y��$o�ͤ�����2U���0TC{ H�i�����d�N�������������M�ϖ��g�@V�m�y����M��M��³�")B�n�v�l��F�L��� �_i\�=�4�U��&3T�<v	d�,V�k�0?]�^ET>���R�/��mQ��1�߅�H��f���t�*E��<�g8*�r�?��q�r��>��� �c@�\��x��=\�dO?�l5b2In#���V�X�e+����LȾ��в���
`�B�!6�:>2�=�Q�;�UԃOE��׉�ra�('+<�&�yGr�,�N��E�	*�l�<�yV$�R���K�K��g���?&#̄?P(��Umz����b%�j�^��	T���S薊���L�ߣ����P���w�=��	���-���x��M�&[�>k��#)Ծ-�G�3$�b��-\Ug����'�Z����N`�eoǚ5�y��%]�)��Ͻoy[6(0x�����5�^" ���PIy��'=�p�L1��?>��[�mj����
�+��OH�Cͮ���bŕ&�.��t��0��ԹuE�s^S �����z�<��!{x ��Rs���`V�*��1��?|�`6���\�f�On����.Z�#��~�C�+L J�!#J���Y:c�/���b
԰�m3�&	(K�B!6)�VHCR�K����_�_��K<�����������X��!g��sܕ9�IohLa�;���S;'���c�r���tD7�,_Q��M�_�M�}�cV����"��R�d��1�+a���pOŦ;ѐ�UT�$���d����
�c`l'��T#�0��d��'%���0�I���B�5_�#?0��7L���lmh���ĳ!�]Gk2uVB9}���@��I��:)���0W\���ҏ\�K���&�ɺ���# yk��%�)�W�?����{k4y����a�
����l4�z��M/��,��91��r����T�\���΀�|D�4���m94���T'В�]�B�v���Jĕe��NZ/����@�'�N ��#�n�@K����G��凉�����`w@_��y-�{J�>�:!�È��8_�@�lAeN�k�%Ə�9��E��| �[�ռ+2X�k%u�����ł��6]�	�S{L��s55͖�+�ouS�>�x�}�KЗ'.\&܆�Ӥ@ʃT�oZVb`�T�m���4�e@�ό��gʟf J@�4}]{�C�`�HB�?�i��0��rkb��5đ @Q�YS�4c���H6~���X@uj>�<���2�TJ�-�_!0�����+����[ w�2���8\�z��ėM�����D{�:���;Qa�l�� ���ˍ�:����~p]*A_u����\O�"#���⷇m(uÆEh�ZY���������v���!d�Ԭ����T|ջ��5�?ԞBn��z�5 (���u]~&�o�����RD�K�)� �D�+B$>9q�~pe�Q+A��^��3��t
cz`|�z̧bD�r�L�)���TX��dG/@2x݉�[%�$5_�*qB��RA��#��~�ZjES�>&r���3�6ކiZ��v�F�;��&� +|��4���1r@[��c� 3��1��C8vlhsڕ�Š~���6ܬ���Y��%�ݘ�$�E���&68	_��`>)Э���l��w�Zx�������P�n1��(��E�"���	V�-��m�e�g�}}�^/ 	��$�&�x!t����uK�n��Y�jb����q)�����x�)<�y�,e��L,��|�.�.Q�ZECӎ�_�{4g�fO)W��A�N2|F!b?�t�HLp�s�^���wB������=g�ĪS\�3���+���['��}�:Íym(�~+v8z����v�o�.햼�S_��;��߲�p�(��J���Q��q���l�=����=T-Y���u��5-��5����9�~��P*�@T� "P��h�P�Bzu���Q>GM+E�ݸ�:늑�����d�kq>��*Ycz=��(L# ��/�6{�;Ð�����T�6���,{�U�$Ņ|s��E��3�%I��d��Y���Ԗ�����m�J�L'�����8��	��������ܥ� ���6T��];Pۢ���2(�5�)/�_O&WjH�{o"Qr������ݠ�m`r/�s�����;������=B�����S�������fr`�4�Rr��c�[TUAh���;���׈�n%����A�����Hl<���C}_����봥A�u�?J��I-��8(�X�^�nX�q*3���&�K����w=y)<P���k�6nh�}�p��>��ӡxSy�u�e{dx%"ޟR�рş�d��_VpֈSj����r�lަ���%mS�A1堝���
�]���
�?��ſ/�T'֚F�X�1���o���+�U���~��{V$�sX���A�- ƌl;�S��c�����7W<%z�e�c�R<����5�c���5�ɛ`I�h�ܑ�|7�+م��:/��]�٠4�/��f��7S��[����۟ g�ӈ�!)����q5�'H�ħ��<y9���Ea�a�|=1/!	���3�<U���QML:$�POZ��T���歧,*;Xhj������!�P��P%�Z�37-i�����E���*(�{�4�����k��0��?���C���ɡ���O��U*jX�����N�=o�}#�G���x�K�R]a���F3N���0��o�0OZ銐�N˨Q����,����>͞�@��]����zk�ג�ϧ ?�p���Z�
�R�:}�q.1���j=�����g/�u��1���k��e�1�T1ee��°F�E
[k?�bP��H����n��CT7E�6ca�=^aajFޗ$�7K��θ���j��˦&z�c=������<(e潰@�/Q]��S�=��頓e�"
!�s��R=w�4Q& ;{����\���F�2Ds���0���T�%fJ�gC@I����Bѹ�m� (���{jѷ�8'�k�Kb�@��"�!l�Ԉ껻5��Kz�`�N�О�(͹���Ϻ�!d�k�p(�P�7\�$e4dꍀ�b�~�Bw)��vD�!y`�&.��u�����r$*���l�Aʥ�z�����+&�$<O�V�*3��h�T634�d������E�%�"�Y#�ּ,|p:c�'8�p�.^:й{Fj��i��*K^�s�l����H��H�E��8m �]��B�if�[��^��c֟�G�}�0F�V�dH�"z�Mz����/�p�A�Z��\e��y�1R�+��(���ҫ�U�o��-�&���_U�X�s�6ڭWo��,}�ￌ��"	[�����B�5�?�H�\���C�?6�f�" �@�u3��6a�1A�i[�dB']Y��O��Lٺ"�`�m_�а�u���^�_�-��e۴̮����AR�����1E"�09CRbf��R�ǃ����= 0w�K��U��-��Ș�e�cLn��ݡ��v�C�N�!�\���dl�9@���2J�tB�h���]G��������=!�����n�;҈`���kv��j�[�% �X"Zz�`�������������~��Uh�]jG�n9t�#�N:v���(nEs�a�Gw�康�3��S�T����jG����sU�0�|7�w�ozWCS� ��Zߘ�CO~}�t�
W{���;�	ÎU��8Gzi�k��}�d���N�x����u��l�w�ud���^ixgE�}Fe�%� b�d��<UU��gdI�	�jD�l����\�	ȼ�C���q~�[���TT�@��C�R�Uyԧ�H��x(vF:�;�����]VL] ��[����
A�Z!OY`����+a�l���4��]�����@��=޲�t{ỪO��͖�ZS��� �ax�f2:�nꠦ�bM ߤ��%�r����)�t/8���&M�AG� �L<�l�GL���u?^����&R`
g��4��|�/LO�aJ�U=dɌ�����lK�Ka��l~�!g�P�2�qG����<��kuխ����:=79��6�$�V�6�"w�rڠ�� '��������X� _�IU�,2�hć;F&L��RT<����{���F���R�m��<Y�u�L��QEFW䤅������d��.�UrV��P��@K��bz��0d��T+�7s`�zd"B.j�*󤬗�u
����ȋ��k���#��ܷ$BU�%����ѫ)�F�pg�E"R��+I���N�g���(���Cp�(b*�p|����@GKz���]o�Y��ձcE�¥]�uQ��5�s2dH�qQ��P{����?�"�||�h��Xt�Y�R3�EIǖ�ai��$��{�M��0������(o�������n��M-�i�c����'��h��I��i'�ã�S���i�qܳn�D��!B",�}��E^'�U��@�X�[-����xu,h��+�&\*�%��1��A����d� &��E�/xz�z�N�o~#�yv�DӇ#:p�e{C��}�M�мlNf%�?�<��7��4i�KV�l��� �T�#9�\�{-�߶�"Z��q�l:q���$)e��1�-�[�z5m&�ĺ&^��怃L��p�{L�hxQ��(����M9Z�����b��	Na��+�l���	+$�� ��i+~y�/�e��r���~�;V�)FTE
1�/�C��l*N��%���x�|��/E֯"�P���H�V���W�e�.�'o�NAv���C�ŗ���R��C��M~kn����e��-T��jV�t���{3�1�Yj�PsB��^�W�?u���ūx�c[��g��j���i�� �1�����r���W��o�1�Ȋ�'@6@���;��3��aWE�����5� �4�Z"UX�|�| t�O��Z�����2��;̊<�p0I�r��Y�m�]�\�c��>�8���QF�
�.T\����&s�J;7�S����]O3=��E�E)�c��	��b��|ni��>��$m��L��J!�`� !%;��7|a�J����,����7)�$����q�� OSZN\��Yl�`�D\����ZU1�P2�O�N��y�5�ImWI8�p��������%��o���S������{�Q�{�8?:@P�"�MuB�W��B���HyKc�������mH|�:�C�y�F^XT �cej�Z&;�����)�8��8n/y�H~���s�g�n�������$�8���/]Ip�(�*��t`/��Z_� ]�?!m��{�|�I��W_>���1*<t��Z`=�gU�2ಸ���9�*:,�߉s+���\On�V�5����v�oZ�o�8�Y��	�x�RZ\���F1���݅uo�#��=,��t����ÀlD:;smd"�GC6���YG'�����i)��g8Hf7rq��JZU�x][�CYP��q�v�t�A�-��څ��Z�5B�Ψ�v'����a�~-�hYG1�Lp�O΢�h��
_�`R�\*�k���� mX8x��؄u��TӣעU�l��]Ѳ�0�ȷ꼵D�	�v�P��lͶ^���NŁ�r�4=< sY@[��БW�xO��e��oF�s���i��צ���I��u>���"�a�����j]2E7+��pT=K��)���b������U� ���l��e��tY��5�s�o�T�-���O���E�SB�TB��x��7Q��W�������WL��wj.�9���=�T�-M�W�Z�m k��Ⱦr�����S
D
�yBg/�Hŭ��"Vh�>9��}�*�o�I8M�ݱO�H|���$���EtjߍbI�j�YW��L�k��N7�P��>�r��Ԓ��Г[��-�'y��[���%�Td"���Vu*�3ف6�"U����w��S?����&<�P��M8)�ޏŒ�T���0q>�483�j'i������%8��{��ۏ̵���R�`뢋G&�Gm���٪܇Q�	��ͦK���ֵ�E�y��%�s_�+�{y�:�?o�3s�܁޻[ ���ڣ��Ë�XN������D�JN��D��!h�͵�{���G.s�*)��ٚhYIG�(/Р�O�ߌ�g�f�@����������N �`Ş8T|�����H�?��б�mp�����ȥ�V�tX&I�ݸ��P�>�J�3B��|�R!�2m�,��*|ø�'��nX���Սy�1���	7o��J�*G�ol�6G��]dV�t���7���^��O�Udl�aqw�7icgk�������f�~Ɖ,ХHP|㐑*����wv3SO P��[��ǯ�M* r�pt���@���H��a��Ef}I8�*�_��N{MW˴���5�0�ͩi��ŴE�������:�ͥ���ނ۪����+����a�êF�N�3�L����/_�a�-�r�[2���}�'M����\j�g2&�������:)�Dw�ˌ�'6g[>�#���.��dU�J�3�)���~�lw3�xg�)�V��ȅQӱS�S��|0�M���aBO<��s�W'��%��]���sco}�n�3�Y���9\��F���,Q_w�h��:ٮ�-�	J���`������$"lBڻL��v���pL)?bɢ���3?9 �^Yyn}'�h E5Apb���q���^}��y"����Lc(K���{@"�݌��M7z����q#�����m�xcnb��	�]t.�=!�r��A�Z����!��#G:��Deҵ?!9ƌ�%��k���s�9�a}�:�����'��r�zu�r�3�/��ֱ�3d��D������K����NWѭ�{�
�$�l�!D�̙�x�V܌٨5�����퉩�޸ ���@ʍMzPNn-�k��qp��q�Jq�����sg����;ip�,+�ڜ�sf��s�2>����w�͹��vZѦg�A�,RG����Gښ[��Tr���"v�~tŞxhQEf�������"���g|��eE�}�Ǆ�ŗK��nq�?T<@����&2���R�t��?�R�mI����=���K{:���-Dcm����v���m��J��:,<���_��5��]Rga�،>6 �ꃙE��7����^	nV����w?2����	�G�?�`�Q�֥��~�A���E;3�=��:U��Y?h�������ڧ�)?#3�}�gY��M��ڹ�S�M�X�lпo;�[��GsOn/�k����@��CUK�j����9@��(ѭK�B�]�O��n�QN�(�Bu0���-U??G҉ �Lx�)6�����b#��}�1h]��RO	�@o[8Q�g�B��\$�T7�u�W�c=������L�6�"�0�B��j�����g,]}n�6FJ̧|=|�x�	$Z��uM�{0��&�Q�L��d��+y�\ʸ��s���Qx�U�A��IVC��e��B1>"	Q2�Y��q>��P�>���xC1��P���h��nӲ"�ϐ+���%\�#���q����BO�Q�-��&���;�ٯ*�`��ѫ������\�`�4���7��Q�q֬��i�@��7�m�hM��1U�5D�3#��� ?7"��ek�/��(�+FT	�p��E�sZ����+�	0,|�Ւɚ�9`�`��an}{!ڂ�iK7oĵ:.R@-��G���[f��IE�2�/$C�<�=
:H���Yr/g�+R�=Il��N���^ʌb��<K�c�օ�
d��9X�?��~f�$��D��7%}m��=Jd�

%��џ�]�9�k�c�U���+z&lR])��# �Xh�f��z�
/��U���7c5���F4��U�o� σ�pu����wD\^[W�`aG;WM�Nؑ�z9yF�ԏۋ:�� e��3OB�n�	����~���,m��]��"�m�p����N�XJ��V�8N�Ry��u��W�J�I�TՄ�i��P����5��,�٩냂]��;�SW��QB�Z�y�ۧ;�KB7
�	6���	s��ts�!$qn�
������������6S�ގ|��ߢ� ���{�����?ty�{�*'DB�}����J�� �E���i�7>�'+ ryJtZ���\�>��0� M��b�s9JJ�6�4����A�k����ti��W�i���)�X00�`�a�`UW\ul��3��x%���k�S6��5�Cv-S����_L�ۯ���8d܉���gE�3��δ&�v9]���#
�H4ek��]��}z>ǂѪ��ahsO��\�8g�C��Y0J���#R�&a���%(9�!�����M7����A��n�q_�s���휒�Xַ��`����t�53�JoZ`h.,A9K{��2�(F��Or�cTHAo�m`Y}f¶4�I��?��d�������ڤ�Q0tT�kVHQ���Ċ��t)����\�)���]�����
�[�8�����
�=��6��yG���E��p����0˺5���J�N� c����A�]���YS+8'7�|-�ӎ�e�8.��-E��.���B���(�8mo�'����-i�!d��_4^V�B?�-��{�c>�%E�K�L�8y���\���דP�{--�W̽Ԩ^9��THS�>I�%��;��>�o�o��� ueJ҈��!��!<���
9y�1`l��3��D6��c1ي�&h�ԥ�H�V�Ìߕ��I�h���v*���J3�w�����,�yk��/+R����F�6�H�e�W~|��s�ǷH�}�o����8��%Εm��q�-!%��j��y]fL5s	�@��]	!��F&�'�ls �I���B����=�b�.{p]�\�*%b�5����o%(�Z�kx�8sE���[��-�?��> �I��Ca���e��Ͳu��l������ȹ��쌼����P!JRCo\�,l����V�u�LTm;t�VNAZ�I�49='��~s�3�,pj���z��"Q����(	J��tnNP���Y�9f�o�wW�·m���!��4)���ƽܣ����A�1;���_$�ROx>��X���K���Ā����m>mV�غ�#?s\��ѹ���Q���˺ѰjW��~b��?��|��ԛ8x�p��x���P*&�����8{ wXO�`� ���c���e��4C?��4#����%��~��MM%���Q�"�/t|c�@T��s�^�1�Ì�,mc`%�~�C��F�@BPvV�-t��T�e�L#�D��MR�<(rR(�;��r�t'����{+w���U����Ԕ8���t�.\~�n���u���f�a���D�U;�6�[2R7��1�t{�������<$u�kF]��):�τ��b���,�
cT�3�߰�J;-.�����S�c������h&Kk�A�vq[�.��(�@d-�!�i�c��HK��������[^���R��F^�6��o%�w{P�s�0�Kx��7S�]_H@7����ΣΨ��A3�ţ�th8HR��O}0�#	0�\����[@�B������4:=�ՃY��?��>n/�	�A� 7P��m]7G�g�o�� E��Q�T�!�E�dO~B&1�p>�O��%�[Y)�B�:�*�Ҙ��.���g��SM؊��1��I�VcV����ȿ�h��P�����hSY4Gw����nh������#�D"��y�^�ܶ��T��L���j_ih��s߀�h��ԁǣ|�'�����6 0J���ƚ�9��T|���b�ɣ"�M���N�������۾����YNr�q��ԗ�v��Е���l�y��6e�� ̵:��×�P�12�@���(B�",|�tM���}�����C��`�]�vr!�F��p�����3��X��[�J�>I����uW�J�*>@���X�]��M������؍x7���� �*�ƜZӭ�^�J.Mo�
R�0���ɡl�Q���Mv �^�x-D4��өf�@�k�!��z�a�
~�Fl]�V)7�G\"��}� $�lPXS�;����a�Fvi_�N&I���+�����_z#�KN���zTTȹL���M��Ȗ�Aq:tJA;���$��G�v��u�[��)ޅy�-5��l�����p�.� ����9u �g=B�\1|��)�����.� ���4~�i�4���#�4;���N��UG9����mYU5C
�H1i�j��Y��~���0B�	�y��V�{�x���J"�'j����V�F���٦2�&���%�����5��G����v��� \2�v��\[�m#1���2�a���i���@�f#�bǚ��^V�U��,��Sd��Q�! I�ɜrJ��ѹ�����İ�6e:�i�]���:5o~�}z��{+1̨!���?�><h�3�a�Y��q�}�⃽��T^>2Pg�8~���(�]��3a���en{)%����T�٬�_	-"���P�s��,O�M�]_Fk-�v�ߧ��B��q�{8������:(�����p����F���oSN���!����l:��,���1mAeK�1FU�qs��O��J��A���]Yuq�n�F�6aG|��`d^l�L@��Ћ���S���p�;��s�p%�Illl�#�����$���
�>U�l*S�I�~���$10��̴3f�
����O()hb��Sa�N��e9L0��;H`��ƉTY����N�B�d��j�f��B�$j�p�>�7d���ON���K��g���i��x<�g�嵎%3�0�SqŌ\G�i�Ye�%QQ����6@(�MƪXc����<�C�f�Z���H�U�*�=t@��3�.j����L����Jd�O�H���F�*t���:-I�쉇��6�N�#�$Y�
s瞘�{�4b�ബ���
AFv��j@�T��;���x�/�J1R�"X&�?�m�~.JC�P��
�Y>�k�Wo�Ώ9��f����^1��C̆��R=F�r������v;��]�P:fV��3w)Aˌ	7 ��rOPw��7����b�,���U	k�)%���	����NHb%Z�f��l~���uT�Eko���&�,��>�����.�X�_��e�Y:!��jī�,7ek�������Zr��A��8Z��
�ŉJ䩐���z�M��J�������l�u�R�_��6��^�١�ІĭU8��c����1��R���p�Q!��D.�V�(����'�!��$�L@j�3�x�fx�-)�Qr�(Ԃ���c�O��S8��$���lgl*���Yw��=�z�`�(ROtçU�@��W��ծ.
��LS��C��e�'��31W�Kn��Af@�@r��3?�[㖫��^�2��g]�kf| ��0��\�LO.�ʨ�aSl�]2��(��bJ|=�յ��&I�x�a����J�)baj��s*~�~��mKC�f�͸�[�d[�3W�&��cɎ3ϳ�5�?��*��t"�b�|�ۥ�J���:�0e�S���3	��s�bv�����k�gD<6��N��#@����b5�i!�M	9a!R�?��u���tkգw�ڢPê:һG�\?�|(��L$�v����ց�*ʻ��3�v��ژ�p�c�9�R�џX���J�`��j��D.sh�%]s��� ��2a��ǐG�R_�صi �B�Q;�͖�>3ƭɄ#�������p�wO+6w������L����i-I�٥r��_�ӡ,��Z$9H
M���;����da�J�M�0992H����RPnm'q��?��S�l����X�b���)�Iu��_����s���¿��'I0�3~*��Z�~�Մ��.�ty��<Ulp�k��Ў��gO9s��K(��D�a����6���n)�C}����_�F�Q�3��ɩ��A鶐b���B.��Z�-���Q����ub�R|�@�Sє;@i{SM[�/����{j�n��멬c�ww�V� �lLwq3�9�M������6;����"G��a<m�T5˽�l���0�߱���I��y"��3�@�1Y)� �6�"�-���"ꈿТ�<��4^��j,�hV�z��ן�W[�v���aZ��@'=��~�K�t8§�~"[�K:&�m/�2���e܏W!�+*��L���<9�9��jۮ��Y��C�i6r��1���T�-�KJ�tՉ8Z��� b[�o@ҭ:��� /��KS]
YXQ. B0�]��x�F�����<�Q�H�<"4���M�:�:�KP���TrVSa]�Ӣ�bB�'1��1��՞�p��#��w!�J�fU�ST��X���/&��t]Q!�[�)��E�x,��y�=�ʨ-�����ɪ?��: �9d;�\a!�8��x�S�_Y��qm9G"����\��{�P�OP��˂��`7�8X�9�/.�P�Xj3 &� ���[JP�֑���լ�� C��f�j�@�~�4��-���C.r���30�g�rD�24��r�W�e/-�ہ���hU|��,#����{b���(c��8��r�s�uC���L)P������1sw�|L�5�;����R�`_�g�=\�	�b���)��L_��EJ����f��[��#���X��^�O(rH�N��(Wt�o��CohGF����<�)_�En��`��7_�e�I�Z}]M=���8PM�A�SɈ,o��LnK�*��4���,H���nd�M���Eq�z��y;����+Y����T~cQ$��.�yJ�C�D%�CC��[�\�p)Q����2��]vآ�	h΋ݕ/��[ned�r3Ί�yV-������6�1�щ蒭�|���	�_����E'�,�:�"`�����u��RB�Ո+@��6�� V:�mS%���h(�@JZ x��o�HSI#՗�dvd���/%��pĖ���(8x��q�j�M���o�Q�/���v/e/D�4��&Ϛ�R�	�'�#��Hv��
}� �q�&�ر= `�a��OR_a��x����9�j Kŷ`����[�]��n�u���"�W�4d�����٢� t�eAEk_Ϫ]퉄�
)�Ƒ	�b��*Z�"�	.��Ơ��r+��%���˽`���M��ϛ)�s{>s�IU�0��Ѵ	:�nzT�/}����1,5
�_�t[����ٓG!�Z���m��Ì
-�3���T�C{3�3� �K��ԟ�k;���g�)��t�����Q���r���J�g��	��G��G��&߭ҏ8��6�S/��7a��#�&�>�(��A����S-�s>�-����f�|l�ƴR�W����m�@!׿�=����7�tň  ^�c�RE����������	�NM�(�V,����u�,�)�v�	��i�i�s|e��3��K&�#���^!f� ة7o��ҋ��K����~�_�J�w�ʜ ��m� �}l�Ap�~Cl�ÔS�~�t��򒗞v?�RB:�/�UTb �Č�e��ziu�h��ޯ�\G��W���|��V�ިV>��כ�p�z�h_A���߰v�H{Ox��X�~(c4	��ܭJ����Q�Bc�����0�i(#m��� ���ꏕ-d�e���R��NU2��Wf�N�ފ������^*͆����o���?�׮Ĝ�duU�ǙzPg�ZY�F	��'�Ȁ�Ȼ��5�����n��`ݭ{b�f���a����	oϡ�f&j����*�_1�w�-d/u~Y�W�Z�4���N��@���9r���Μ��p�Zl�w=��Wy�@�[jx|�޷7Z�Ձ�@��7�Q�LL��Ƹq��F9��yRC7�c׽�:;�;10�긂Jf�n�%�j������a�f?�q-�&+{_����G�h�QA�9u��d�P/� ؖ˕߮�����_��VF
�aq�ÀA�+���ߕp�8+E�z�K+�n�B�s�+�~D�R���e�	��]fX(e��Fvr	$�.�_��Y������*q2+���ՋCq�T�5��A�KT#%�j�zE��)V;���Y�L���/��><Gå��y���X��6Lx\�`t� [�f���o�~H��������#�7G[J�T�^�٤n���p!n.)4��#5&��g7�@�&,MZ6������a����`F#ِ���YH�
��#sS7f,�g�.D#�ҏ�O0�>��^N^ڪ���7s7�	�� X!�W�O��$��%�b�",D��yMJl�]�,klU|u�nP����{�ND��_�J��~ur�	��5�0�(Ō�;V.�j�r�^��)P&��\��o�!��~���.�{��c�w��L����Q8�b��,�s�H�C��e(D�0�'hP!yq�p��`����^d�ھ����W_�QD���	Dv��ж,Ɓ�����-&�{��C��&m�mLruyۥ�h�|�ϣ�\�������T�R�z),?7W#��c��.� �SX#sC����~A\{���q��hE�{����bj�o=��H��D�т���*(��}����T+�1Q��T��?�?��_��F����b��mé;\CZCZ�xN�[ H���\��;�����$����ݶn�X���׏d� ����oMJ����C��sG���r%*�)/i��m?�϶7�Yd��x񁘿}��� ��� �r	:N�)��m����罆��0I�g��G����Xp򖫘�>蝫��u�@AQt� �� Vx[�� ,���ը^�bԆ�ɋ�7 5�1Hu���ݖ���
�N2��9��������\tB�R,���ؼI<hL�U_�f޾�| ����V���\����ԕm.���.wtZ�� ��5a��C�23&<��e��dL�N��5=b�D�xb������s5���TQ�yAC��ȡ���8��k}(g���=Q��)y�����XJ�z�ˢ�����^�!RS���B>h�P�p���_D3��:�%V�mLx'�����c�%G�pY�>�-@4ʷK��5���p�FÈn=�S����P������5������C�[P�ۓ�t���e�����A�D˅n�'\%h�2]�˧[��&3C��A��������X ѡƩra)5���\ׅ�w/������碻oRH�����,�v��A/]y��zS�={s��p^3�˹� ܏��Jr��
*B�٪�z�Oc��� �����1܍�K,}`b�D�Vۉm� 9U�X�A�m�ҁ�W�#c��n���CN u��]t��-<FQ��B�ϻx/����I�v�_]�
	+;�֍$�>_o��x˒���1�] ;��rp�^F����+�:=K��_��L��+�.���5�j#!��
Ʈ����X<	���r���{��Y�v[�s�d���jnf�)ύ��A�a�G;�pT��10��}�[6�������Đ�= F���v�k�bs�Fz٭/K��F� ����F�� ���M��,gvc��8(�V���H&K���m���2\]4����Ov��qd��F�ڕ	�]��H�eY�wErȓ�Χ��LNrl�^����0~3�j�߱��D
5�	�<V�<��V�J�EWV�5�*�E�)>yE܈�!��M�d_���î9IsN�6����o�����@zE��8;�U�'�|�j�k��f0�$�D%�2�d<r_1�8m�!agɰ,�F�b��������}��9s��k���;�[S4:etj`O�Bw��)2i��4o��T��&=��Zq[��?cK�X�
8A(�u�N��U� {�*�S<b�J-��#{��ᱞ�Y{�
�a*l/I�z���Ub�tx���Bi�8��F?�����ia�Z�����|�d�j�ҹTXa�H�l��?�"�u2O��
�K�(^?*e��. s(�:g?�M����N��٨s�t@�����[�h��fp
��e���Y.�VS�h�]�mҤ�g0��kŶ�@��)���Eu�����b0l�v�����-i{v��iBl�DN��b~��2�|GPJ-[*���Y�a3����1FW�*���!
�a�r'���e�Zf+��	��zĵ�y��1����2��]���/*�D�aY���u"
���j��gw5�if�@��*O��3cI`#�oQ�QvA� m�������kY����IT��ř�E���FF����R�+C�BI�b]8�Z�?K!��Sۓ;1'��|����W�AX��n��9�A�a�B<� ��C�t�e��(���v)��K��v���T_y�(R��d���ձ>��IF�.�^����4���&V�ނ��l��t6Zd��nk�&+�0R�.�2���un"Ыm�K��9��~�X��J�|n�ڂ�Eu��|T�	x��:�߅BѠ�g��M}Q�O��َnB&�>�f�;3�`�Z��n��W���
�tO�`����I?�yg�iQMs%h����(-�
9��s�Be�͞;,	�Bgl�+��^�_5�������y�@E�N�u�<QL��=��v�us�)4�F�"�A,���Ϡ��ݍ�Db�R�����|�}�#׼SO�#��v97r;��T3	��i�)�i�י^�=uHA��{�QR�gkxc�8���Ӣ9�Y��������O��Ͼ�����3bh��?�&��0v�Ź`�7�V�Q;����Ⱦ+���ǳ�eT�?Ѽ�y�I��`I$�2d�՜]H��0R�1J�lt�fҢQ5-�y�t�	�g���qW��}��	����XL�:���ʳm�
:�mΠŚoҟ��UH
�0��ٖ��,��jx`�ʀ���0�eT�kz���n{��_�F9F�
Q�iv�gt�1}��5�o�E��"��L��'D�0:F�3�
�g�r/���=}�);�b���\z�� �gc���1�B��W��l��`۔ A�@d!�b��v"��\�X�(l���]��M7?`+ 3 ��Y�q��*A�� �	�&��oZ�lx��G��=����#���f��%��|k(d܀��d}
���B��1����mս�L����:,÷(��莿�5o�V�;��M��q���;����"o}�r_�J�P &�1��)��c:iI��$c�1
`B^]�b��gFSaT�,\nQ�T�>H��m�L� WY�\�A��!�z#&$p�}������̛�p�m������\6��H�f��ւ
� �F�/���J>T�vS(���S�q��D?��_����[�U�
'�|)$�BP��)v*7h��4��|���W������14���Lu��M��j�C�{�g�Q-��:I8���e�f�Hݽ���h��'R���s�/��4	�9>(�Ɩ#�uCU�YZ>֢ʹEn���g%�X���2Ǽ�������K�T�M���F ˭)HE�&=:���l܁3&�/1�U��ĵ$8��uV�ɥhqE��>g2h^%���Uv<�	Hq���Wޥ�����xga#)��a��}�#PVF�ȥ�����z�m����˘k��;����{;��!& �#�3`������z��f�{KP�x���nw����E߯�J�,����=�z.�t�$,��N/ݪM�Eͻ���ouP�|f��T� e�MJv��@v,�A�
�דt=��r BrU�V+3�Q�n�!�����c�A5�:u��P/}9�b��/܄�j;������d>K��\�����ob1�)m����9��^�ԡl
 I����`L��-�v�K�(��CB��(�kR��ʐ͊M^eWnإؒ �6qE��'�;o- po ���[���O\a�Pݠ9~��SO#f(���a�I<-o��Ԣ�k�����R)D���#p���YTK��{w�ؗ�V��m�����R�	w�cctE���������ˣ�ۃ�_6��r��k��o���P�Ľ�I���|��=݇�����I~@�~0��n�P��b�!�p9\sU�&28��;��^�G_* �L@߈|N��d&��"R��W_�l<���ruev���������h�R���zeM�a�6���DMu�&5���d�Y08眠8D�G�[�6iM�f�!��P����0�m�s�՞[����Ia��P}�86Y�tt/
}���� ��.So�jq�8Zo��X�/n:�+��j���TC�`X��.��j����N�4��'���S��Y�-y��E�wT�5�3�l
8�vu�k~��U��ֹv�z��ΐ&NɇHJ��1�Eu��`��i�(/��D�zʤx���-�O��䝧U�������`�� ���w9舾ޜQ����{�o�����/��Py�V�cvM")����w��*Srřa�3|"LH�4[��l�:��}�!o��t�RQ"ESfD(�܌	^�2��jQ� vعvl^��V�M�Ҥ_��Nv�5bAx2�(5�>l{�H\�M1�����ҞZ;~����<�>�%֩��nxb�7����#�m�{s�0�#��s�6ѫ�8ڨ��uW8�LI c�kI9H~u/��(;|�=/����\�b>X��?��P.wp���3�ї���Ԓ��C�Ĝl�u|P���q"/��^%JQ[�=���wlw!��7d,FvVk_��#*�0e�;�e���
���k�y��Gf�M��%�g�{��Zg����!�q>���w���1���n�GT�ܷ��(��`M����s	sL[İ���(�Γ~e#.�N򉀍R��H�&�y���(��ɄE{0���Fi'�f�|�ܡ����0,���W���	�'��L1]�O��H�A.�L�c�˄�0��'��6Ņ��N�8�)�Sr�BGD�� Mo��2�/�� ��5�x+��)��n���W�	i�s�4_{�$K�+Z/���a��m�xId�����������������߾��2+�}����z���zW2�P�����F�FT��e��Ǻdo5��#L�#�ËL�`���a�Bk�hw�,��n�d��H��������JDY�!J��$	�ڡ����n��0�ch��sH��^���3va`�`4%�1�� �S��?��5�ː�7�fw��C�v��f��.�"fcK��y�ƥ��I����<ɒV�iv ��`�(�	�N����'Z4te�V1씕��V�v�D�D,g� x�h�w�0q<�	W�\��JĨaj�C�"��*���4��F�R��A[E3�a��ڿs���u�,$ݔ88����[�㤃�pۨ���mW�>'��@x�E�{�s%��˻3�������x�h	Ϋ6�5�~�E�F����&��(�lⲟ�*Z&Kl�W��P㵇�0;D�|����-��ǧ�T,J��܊�iP�c�*ū��������3xǜC�m���Q������ 6ѓ�kB�+����R�*ħ���,h�����������|�m��-ib���0f��i�>�8�,1�4��?�QQ���pf�8p:�D]-<X-mK?��jj�F㣃��ds��SN,�+�����;���$zd-?�'�#c �����H���<�1��1t���լ9��V5��a�X��.�kS��^!CR���M���2���� 7���[��Ӛfa��i���Ս05"�&P"��e6���n)�b��YSo�5Y"�Uޟ4��t9%��$����O�� i��h��{�O�[d��\rp����.c|ALnڱ�7'����Wv϶|��Qb�pln�ELD˪�t�����4��L�Z���t�F�Ě�����]�V��
[n�T����#YjQ�J��X�lO�Ab.^�qD��t�� �!S���l&B��1t�R����� �ɀz���A��"�aQ�z={:ըRƮTqy�{�Z��T}���:j���
�=�h�,��0t��C������h�!��y5�ksr$���{9�쓘�������
ax�G1Z�]���dyO�e�9�����O;T&z.�L'|h-mq���m�yq��2�Y&��G�����~b��4�LK(~j/,�άHQU���@��Iĸ�' �]{��P��*����qtf;�����hz�V����s���Ė�dp+�'6�i<#���'aq+��z�n.�S
�R̭:��Yf*h�	x���:U];��/rY�į�&ճ�C5`EL���������MV(HV#�k�ȭ�7�=���I��� �)��D�������PfH]�e��RD�m���4U��+�2���	��jY�&��h?ꢦ�!p渫����sg��{uݒ�/�r㮭<���:��O��R�r
�(�� ;8�~�z����� B9���R�Uo�H	�FB����?����T�4��Ė�|���LۥB|OD��,p��5�Q��6���lL�6��Y~����\ZF%.��l�k�yO�ʘ{N/�X�t��5y F��/ă��zL!�J��r��Z��Oո �ib��NJSk�ݺ�X���e��/У{�8U�3ra���Z��~fc�&|��� �z��;�Y@�Zo���nQݬ5�:�k��˸�ԯ�����hL|�U�%G�a�wqߟ��;��X�'fY��ӳ�u�����VVQ�*"���b�s�+wy>�*�{�=O�w�3.O���ZtYv�;:x:�
��-j?�߃�G�n��k�'��"�RxԂ�)\��~��;e���Q�H=H�W|�9���$���-E��*� 1Y��-nHG$��i�iA�����;������ ��>��!��b@O�?�h˅a��&��NI����qdX�=3���z�"@V�/~�=�FЪ��*
�94��\�"�=�����)��BE"���&A��&��1N١y�L�t"k?����>��"�>�(#7���v�#'�y��9��b-�a;2x�[�G�I ����ﱸ�%V�m0����H�#�D*�?�LH�1��b���������	~}���Ы��
�@�C�kc�>�₇�e��W�6��bێ�����?.@�����q8I�.7�6�'b�D]���]@{4�V�/�C �\5[����lZ�?�C�>wG�i��ð,��b@�;���rKs��;���G�p�,p7R�t�?CY:��@�kY
aDH��1���Q,d��\����P-j ʆ��p�U�P*��7����k�%ף����o]\^:�,YI�,@�[��� �>��Sü����sV�j�6v����p�0��Ud

�Y)й��X�g�w}PzWB]!��ҁ���4���`�dP�.՛n��Ps��D�ee� 7����5��n&��У��� g��}�u����A�B��@�N�	7�b"$[L�=h��m�	9o	ib�u].�heȢӪ�}}�=�$���;Gdx�k��g	h.�9p7l�'��=�����C��Lʭ;�i^mE�T�@A��IQb�-��le��=plzߑ�p(NNC$��:�%p;������lC4h�F�9�̌~�a!��1F{\��T��޲ĭf1���X���4�[�>� #�ab�����^�& (��@�?�#z�g�$.{\�x�v����D�."�C���
�p�(Ch2�q�#��9{<=Q����v�wx�+�7JK.�k�g�l����|�Hsf@�ͨ-�;4j>ʝ�o3�djN��+J4{33!��d@A�1��Gf�FW���o�o&��N�Β�Wq.�1IM�ʓ��|�QeR�`!{���.j1����?��z1j���,�Aן��}����]��-�?��(��$Y-���?�������@�/�k,]��Zg$�$�������L�Ϳ���,	\��%`�B�O��d:Q��`:�՞����V*��t.O��p�$odT�RH'4�!�5��hX��Xެ�
�M�\���yE�D��LǫjՋY��QØ>E��w��1�����V��W���6���l�˖u_��O� �I��j$� u���å��%q�hl�=d)T�杣ܠm���(��#.��Y+@6��h*��j��[��BE[�b)��������5{�H�E쯍�rJJ|@�*��o����--�X��A�ywqŅ�l����@1c�q G�2/0"�5���Py8��ᇗ�U�%��8��A'�Y7^��40M�{U��~���kv�S��<�?��M̠��0�l<��n���^p��;�6��Wͻ������t��%�����<A�_� (�L�gy
˲��G�A�=�n�+���+)�JD��<�z����T�dەE5"��r�ؤ��<?`�͸�n#���?��ӵ�O�N2�wI���=v����㽽�I�e)TPO5���`�gu������8���ͅ;��P���JS(�%������t��VȰ�R�ś��.i���A�W	����t�`9���ZZ��2#�o@T����,J�͢��
mD���P5������/�0�UM�5�=N�%�����+����z����^����MZ���y���⧈йH%dJT�DZL���%AO�r��lٛ��2���O/�����҃H��/��rM1�R�BP��t��zl
U�c�04U4ȴ��f�NXd���{U�")���td��}�־W^Cm�yx=�m��\�%G|z�n�	.����8T0Ĵ���5�H	L�KOw_��o��_f�����Z]��ǵG�M��� }<.�*��y3/V�dP/��-�I�r���U����	�z�Ǟ2Ϗh% �|"����Ʊ:2\+a+v@�]pu���c����Ѽ���9��n��퍃�)�x�����*c��g��+N~h\H��8o|�����[{X�b�����";�Á������˒I���$�k��N��'�S�:�PΟ���A�c�7%�p�U��[��8oY�\�eX�N9�N��(�Z	b�� 8�7�pwo�k�p�0��I�!j����Ts�� 0�ӄ��ɒUQ��>kF�X����9� :�h�^�o����^j�'�AeF�F��6���3�ß/�-~i ]L���)�9鲢F��Dz���.�&���f$PcUi˪�ZX�a(vP ?q���&�����RV(X��5�Rx�Y���a�v��yȝ��#�>²�C�7?`��4�G����U���,��6t�ȱ�"��vr��XOM�NA��AO�G����2;��D�߬�4؈)zC�z�������
a��LT���d`�}�*�Ð~=b� �N�ݯ������9���z/���U���]��B���|�{cX����)n��6����(<�͖�m(/���*m�|��%��*J�>	�ڏ��J�h��j����9�1�vض�d7j�UVC�P�m�7]w�r���xR�o�$�z���ȖxNM�������Kn�Agrve����|*;�-ѬM(�����,�PS��2�<�t����yͽ���)/*�+�ϕ��&���V���x�TIF���[��:�b���P11��!�O̓w�Z���{r,�������GV��X���FO�<�����CE
*��@E����	����3��;��?�9G��xĻ^a\�V)����9�W���U��w�>�#����;���b7���@�ZM��4�=� ��'�%"M�:���Ӎ_��p�m*�}��+�&"�FZ��m��:{���)vR14{���X.[���m�"�+��YT�zKj�R��z�@��do?n��l�c�� �^6�+�Z����g#�]�j�x��֒�J�n�MM���[�C83RH`��G&2~�VT�[���2��5}����@������z�!.�Cu�]���K��K��Y�r]�r�tg���3_�`��\!�%�$)�'s�bm��>�|ue�_�e�H�!���Z���A���m�?g}@��Is���9���>j���'T���b�SپgQ����W�C���M���xΎ]�m��S�Y���]�����f�����G\�Z���ǜ�2��h^�TWݢ�tp7	�C��&9�4'B����X͗@]MnVb���j[L�Z�ʟ���gC*��;4��ǏC/Z<���`e��� Vw����c�$�#�Qp�U՚�p����RY�"U�;3�����C��u�m0��S4Y>,���|�i�h�I	o�
y��5�<�1|nGT&e��'Xxb�]��-������u�V�`W�s�Ɗ�4]u[1��I���,w��_�(nz��xa�?�(�S['+z��]��>�V.g�lb�̛�2W̜4�جU�Pیk ��L��-v%-p���.���ັ|6�<��1<��c��۝Sg�A|YW��^���b���i�zC�.3	Y����O"X��� ΋B��Lw�R�W�ގ��lq}�A
�h,��otƐ�/���)y;��JI	
E�ӥ6V��'�L.�g>?;��^n��y#��n�p�EB���(����,�H/JJH�6�P2�1�jr���z��hU �d��+y�5]r�� �ҕ�p+��Zd�!��s!�4]��'Q���@h�=^;D
k�`�����gF�f!z�x�|޻є8�>M+� /�78�n��Q˼]��b���:ejg��k����Q���T�8f��ͨ��6�AF�~���#	��?	0�K�9���z�����w:��F�2��= b��ȁ!�x��1�;�����*lr+�'�0Ɔ�CK�b9&#j'�qi�F��oQ'�B=d�r{�ŏ�P*5Tc�.�d�#���Y+��4�`���7X-��)immq���¥J���5��b)%c�O����'!�2e5$�����_�Z,��ߒ�/�@"3;�]nm��:�zft���}�6���bhQڄ ��%{��-9;�2/�~R�����j������7�����H
йYO'Iߊ�_��s��u38��}ƟT�r%KO"V�������P�`Ghd�?Ƨ��a��4CAj�K#�f�ٝMn�b爍��h=�3��)V��9�B�2���8��)�a�(�;�B����26�3���"���$������8��V���j]0Y+����DN �O��]fI�X���j^��6B%zVJ���p�+�?%�bhz����7�� �P8M#ګ�N�^$9i��l�$�WX���{ˑ�r����A���~r�_�/tN��U̞��p["fM�j�\A(A�1]�8���:��3��-w}*(��3ţ<Gt��v���ܰ���U^6��/e�;0
�.�Kᙾ���݊��rL�\SP!
�K呗�p���~S�B	k��0���"�N�[o�eLK��qΔ�4��uX"�)�1t^j_����x�L�����BэEI�F�����Bjb�ʸ�F��������&( ��,�߫(hkM��o�Ş�l@�t?&M��OFE�N}s>�s-�o�dF�<�����p�U�,�1��P�xĥ�'�BA��t��A!��l[�h��u9�k1 y4���͝��~y��5jy�:��o4�sJ'F�l����&�̉�b츻��d^��IW�fL�*-�����8R�`0>��?�97�`о�%<kt�J�6r��8���B��?���+P��EW��|LP�j��:����<W���9U��ϫ:���;�֑��T�����`���r��~���L jyi@զ���XK�=Z�R�Sˁ>���D�ΈG����p�kKS8��6�0j�d�V��ͦ�A�U�޼0�+��u���I[���5h��!u�Ջ���}�Ix�QT��`��n>���9�q�ϕ�L��_�x��cw&�s{EF��R
���1x`p��P��|��ä�'��o��Quⓢ\� �p�FT>`��{���Qf핅K[?���;�my|��T�I�3�/S^��!I�� ���sjL��|v:[sf��:nu��!tc��}���$�#X�E��0u�)�F82�n.H�j�IҲ~j|��j���œ �]�\�Q*sY�*M�Ѵ��㈹>�گ�]�����nS������kw�V�\p�!,f����&��dÖ�3L8�L/�f��}�9�Xߊ�ߢ6'߂O�̐2(�+�����9`��;�ihh���PȻ�7�k�~ě���p|�?�����E|��;k�I';V�l3�~�Ǯ;|l��oo�`�ؼ`��.���/�W|ye��2t#ۭF�흡S~�/���G[�����r˃Sٵō�[HPel�Dh����7��Ж�W��>���Qbx��D���Ԏ-h*�<KP�b�[��5��im�ӯJ�Do[ǊD@�~� ,`{�M��ZG�'y\P^
&Ԗ�J��3H�dx�=�Ҧe���g���NV�j�uHNe�cZ�?���)�z�!�y,mV���UM���~I-5�z7�OٌX@�(e���
4��BS�-#���<�xn ���i��z�_s*��C�L�KT/V�@;!�]�y�i|�������4��J������[�c���qU��R�v��ƶ)��[�%�֌2�(l��)��1
��k�Z��Kd��e1f��K|G���&���_J� Q�|y݉�@ξ��8@c��|������+�2Қ��
4_�\W��!)'�]'�fқ��
�Kg��_�&_�j�z��(��B7h���%.������5Ţ����&ce9]�*�!R�+��d:4���|�I���t-��CU��ج��I�g�������$ᡞ/�jz�-���q�0���
�K距�Z:�`&d��*0?Z��v$4r#�P�ݰi��Z���1�l���Ft�0��끚h���L��� ;���e�������R�c��-Αy#C���+i�Mo��An�uu�ZLCu�F��M��ɨ>:�͂1��Ng�+|q�%�>y��Ɨ��q(��O�t�K�Zնꨜ��Q��)o�b�U���6YX����<�%�SH��*��U��0eI#Q�����2^P������!���a��w����D�JZ�NM�ŚYp�͉���<U6��Sbw�e�f���,�� ����j�~�I���vtD0ii/b�̯��P��w;����F�������ޡ�<�ۣ����5��=N�h�`~��a��}��*���W<!�{���WR�Vۮ�dτ��2�T�������~:��[��$	�a���J��z�ˁ��rC��ƵE�(�c:`ik�HeL��*��-��K�w1"Yxc_���F�rDH?�V�?{de�bbY��x2��a7�0����ɻ��x"����QT{�E�z5�e��~��`�eAV�{�8tA�š��9n�S�c�e�zǣ��N�ο�~a�q'�=� ���z�>�L�зʸk2f���Ӽ$��=�tvF~C��Y�^d�K��+� 폅P��-�1Pݣv=p����S)c7����\Xj���;y��
���Z��|�ųQ�7�����z��H ���uE�h�%3��Doa�o�Etj�����R�&���8�����3*�|4J��Zds�uOD�t��ݧ=�U%l~���0V���!��.FgjV���nߒ/���ֻ��n�q�f��KWG_~u���
���LsU��YuQ9��~�����ɔ1��z϶y���'�/w��i��L:1zboL��^iw�Q�f�8��o_X�6�^"���+�Za����z�UP��g�#M����d�ED䝳f�"�/�0��-���v�#�+�٬���.���≔�"��.�l��b@) �c�ٳ���՛C�����!:Eeqr
�*c�k���,�pCoX��������扁�V�S��iD��r��d����[���7��)���!���ߍD�5������ɂ���#-�a7�����;�'�cH�m��ޤ�@x�-���7��P��L,v��"%��U�V�C��+y��%�����B5`K]0��j�~�@%Wy�DN&���/���o�V��>䊶շ@��#-���!A���o�{�/cM��E6=A���<�hs�&�[~�!���3���/]�8��M��5G��ŉ���p�9��l�E��?0��E�=2�E#ې׆yL�{�ѹ���b�^~���x�2?3��P�ڳz���H��%�#V������sAN�0��
�����ҎѠ��B8[�C��q����Qu���Ms/���+ۗl$�۔ڬ�wRk��n��="���C3	��2M���&���9-�um�<H�V4�G�R
�75���#*_޻���ra��ov~S+��Ղ�X�r���6�u�%$�� �o��i��	D7�b6U�?n�z9p���O��?hP2�T����4�	�꠫o����6�b�%X;y �+�86�z9A3濃m7e&_4�h�ͻ#�����-J�~���HR�H�6x˚��D��n�9���V9��&Z7��.���Y�mj��fMkwZJ;�:P���=���B�ƮG7REK8�k����2jS�):
d���m}ë����Y\$D�}��������n�� ����GR�2��M˔C�zawn���3��8���:kX���=�6v�qm{>ûu�`�i-R���K�za k��2҄͌�a�Ś�"?)v{h�o'��if��3��_�)�$�}!@��%�ĆzK$�*�4��),��7��S�r(V�>e�zΈ�jO2!�*��uv@��Ò9xZnb0Y��rG}#���R1��D����h+���P�!d�5fa������y`oͭ����O�f�0OeS_�C,�.~��K����w�&���Ԛ�M>YCu�aoݜ`Z�����R�@��r���J=��e��Op��4�MV����=(�줛�������#��]��͡ �w6N�s�}k��P�Q�P�e�����tcH�F2W�O٥�;��6U�0���,�n�o���(<Rۊ��K9��sG���6j���8����#�l�"P�1s�B$|g������Ϩ��n6=j�u��x���A6�r�q;L��U�֛�?��Q�2�s!>d�nŷR�i-��=W1�4
�Y���:�E�#J���H�g,��3�m>�??֨Z����[��~N�>�vߐ3�^���J�el�7�nX�n�׋�Ͼv��$���|���� �fgRk��i���<n?P���B��)[�ם�PeW��HCU{>� �414��{�y�?��9켧�ԉ�@[�a����YA&�ߕS�jm��B��6d���x��Pr����{-�!���Np��~��B��$�F�E�lW�J���_���쏕>��"U�6�w���8 p@�z���|�G��ߴ�e�w�&��i%�!�4-�ܾ��1���o��
6Y��D����F���yN0��2�5������T�
NH[�=5sx� �g���NK$,�;����XN��$��,R�"~I��)R��Ar��C����AE�%z��A5���/O�V��ԨH^^Cl5^�K}l�k�khXr }.��j�F'O:��2z
�R�}9�j G�bf�2��׌*ip��0#9OcBF�MX��r"f���4�G��O��ɘA���`(� h�}�����4{CAx>F�Z�]F{9F���i��me�g�`)��`�i���|K!���T�8�rq�C����jo�X���"}h����)`܅C>\~�e{-=�VϠ�h�GLaE�Y�̈́��@��\L��@�	����P�.��=g&��+��^�ގ�`�ݙ��W�w-�E����d*���ª�"�J�����(=�w�j��aJW/� �3�!M
.-�-9�qx-�H�!��M.3�rGk=۔�(�n��認M�f��'���pJ�����)U4����J�1��L�544��v+��X-Or��Z�7��@�١��ů)r{*
�ݕ��\F�v������@ټ0���͇ML��Si)m,L�]��y�G�5�O%��n``�H����Mpv΅8�S�$џ�$/������"y�Plf˂|q��V��T�ԟlL����H���ص$�P4�7�Z�(����}e�����M��ml'_���\!�4�ߵp?�_+�������ġ�PY���+ð��\7�iI�CMR���bG䷹Y<���ѕ��Ʊ
8��.L�C|��J٥+��?���)
.�L��ʫP�=҉��+g��OU��%����,ߘ���6�3*v�(ko$�V�Y� _�L�MҔ��E/.�X���O!6���-|��QĽ�	��u~[L��W��-��Tn����/$78l��������!�/�s�+�������S���ޤO}��{s��(�\��4CY���(}	�i��IA�&�������'�H'�p5Z�;��D�(�<�dm�n�Љ����Aỵ��u3�K��u �qjT
?8�(9�߲-�p*4'Quh>$�
�׭����l�N�����u�)�6z�ϲ�mܢ�{���H�\p6}�ݢ�����Q%^��ݟH��v{���wxH���?;�?�4AT��c{��&���)����_�7mc>�Ќ���k#���=��:��9�^����A��z�/��Mg�Hc�Q��d
ts8Du�����bI[A��HDY�k��YT o��ь��*^��s��ԥ��lSPX�j�q��"!��І��Z��]�	Zpd��T�P g@w�Kԛ�B�PϹ��e��z�^Õx��v���������\(���\�X�����4��.�� �J��+83U`��q�T_�Lo���DZU櫯���L�U��i�gVȟ0~�U���4DaKc��'0�ۮn.J�O��r/�$��X�Ȋ&�+<��?=/�uj���(�O�7Z3�����8~ DH!�󖔉��)g8��	(@3V�֢�ȇ=q�NC�g���%_k z�5�����﹡����+����7G�6eh��d -���IB�p�O��M�(��t��/@K����7FKb9ibhS��:���1R$&V{��
T(?̮,��9{�G94E6�z�Z{�4����-P�D�>��?���r�vD���js�#X[���c]$x\��;��*��Na.�m0��yMnC��0�T48������R~b=�r,���x�>��M�
 �j`GR��O �7�9;�����'fm���h�j���<��U����������g/\��R�*���	;{�KفV���Q�M!ø��Л�UE��T�R��6��)]�!BßU��E�8�����~w�0D�X�Ar�������A�L�*�YpMezVP6X�|r�[q�%����k&�T�(��z�͓RE��w`F��̅���t�ߌ���n�4��*��g*�ZO�w�@l�/e,��E���n�KE���8}Pܚ��>����ܨ��<о0����s���aNw�(�#�c�Q&�v ��)����*tRu����S��!Iy����z�Ԓ�H�z@���L�@W�zi�ׁiZ�,J�7QKBUr�ͅ���d}���� .�N,	��k�r;��i�	A�P��'��=b@�EZ����ܠ������ӫh�i�шH��6IM1��>H/�6eɐ����\�Y�ݍ��ɋ������jG�Q!�&�K��;!�N�>6�'�V<��Pt-���"��Iw̳��>5%t��+b��<�@5�"^C�h�>�'g������\D���IM���|
&ec/,�:aH�#��H��sY�خ�=�7��@����Cr��|`���m;��L�i�<���S��1����P��RA��63�.X�o�����v��H]'�c���&_����ZĻ����:��h4�3��8?�Q��u��R�����k��?�r2��G�K��/ Y(���V�	[�\N8��R�%�T*�0���V�x3���I��~U��ؿ,�9����œR�9v� ���(�]��#�1Gm�k}���h�S_H
��6:ĤX��0)-ߒ��͆�����H~������;U�����3�y����"�d�;uň�E�8��ws�͇)_�G�I�j�d���M��Sv��E]?��%jK��������ۍ�EfHŨ��X�0�G�x�D94(�'�r|�OrvAy�[Wۀ��"y�h���+{c�'����uyWh�S�%��5��)��V�~�$���~��k��̃̄(�3�˞5�(5+_|ѭJ��K�E.�_�Ujp����B��"����`g���XX�o��@���P��o���}�$H���\�[����*�����_צi}NS�5|H��G�-����ݎ�۹��71���Ȅ$q�b��&�� O�ų������Bd��kWBF�\�����t��Q�jX�#��AE�	���,G`�.S{��/'��eB����E��{LK�h���4�]����b �Ny���ΡZ� ����O�"MU��a<��>DaJ��2���&M���g(��Ya��I��{�]d�d��ݺ�O���<־��c+�G5V�ۧ����w=��G*�z�x�dC�5������		������Y4	�F"���~��Dʙ	p'b�����1��^�ߏ�n�?$��-� )�]���a��$!���#���a���*�����&�@���+^-Ca�7����9Y:���3#��V�����wݽI�O�/��U����t��r��Db���=o�xi���J��UO�S�#S�LQ�Iu����5}=�,��qn�HB���;��?#��6{_������x� ���A~����7�7,������C�<E5�� ɹ4��S�3�i�^�1��R�MlA�/��P��7��fs)�"�?����O(��M�N�|�c�j�u�����Vt���h��E��An%�7\K�E��S�	�J���_lk),�l
�<���������9gѷ���xH�[a`'���&�E���4���L�����2��ž�*���Fc�8.Ue)�<�`������-iE+�P_:Z����0ĽyӲ*_^x�ţF��ҍ$�n�+g��G%�-Y��;5L��_j!s3��x���z�%������^ۄ�Tr��K���o�k`�	��@Nv�I��E�>z�3�9�D՘�m�R�I�B�;Wp�a�w����)�c6�ɧ���(h� ,~����3e�%�uP���%[�^�d'.�w) ��[�oLW�֠�}��8�
T���Iqx�{��mŴ�-b��1����8�V����]�V�:�5�a��Mpu���jc�0L�?��E��De�Q�N�����x�2��3*<�;��5s'edC��
\4�)C��mFf7xl]ʯelp�?˒mW��i��B����k��*���Up=�V�3w���!s9��.-?�$���}�ل94��/Ř�;�0��v	� ��?[�����O&,�'�b���"���2��N3y��Yӣ�PL]����: �O�}r�SS��>a������|g~�u�s��LQ���l�3QJ9�KN�׊t�Va�޵r�"ľoլ`�M@;�7+�p�Fp�^~"���iyO�FW�7�?�!���諮"l��w�=I��_km��?�H{����y9�}���o�Χ��	�E�����ɽ��tX���R ��u���$"���_Hd�%�����mq�&�/Y�I�X�+{�I_L�/xh�yC��	q������Xu`b�B��A�7��5�cLA�b4<L`���$�����Sd�9Y����n�<���$�#``9�D��ڸ5��|��K`��R�vW(7ܪ9ْ��?�:�@km�_s<O���v�����ǻ��e���7�_a��\ک}Wf����~:Q��?��.�Q�W���Ѥ�,��|4�����'����P�o�Z�O�������}O,%+v���՛q�G�148[]�q��P�\ؒ
h�b��t��w�eж��E����4�{� iǱ��<���y���\�3h���ܯ��r��GD}���[2��2�i�,y�x���8^B����Qt�yV�j�yt��o��L5!7kޭ�)��m1�����{!ڐ7���}��� ���W�����O�%��б,$G�,G�]ܯ��BKD�o��{�u�w#,�&c�t�"L��6^dy\�r��ل冇1։�<��Of��e��܀����z�B�W/�@#��v;���*��c��3����2��t����N���T���S�~�N�\F��%&�qxK��.�
]5,[�m�S�9g0v���r/�<S��k'�< ��`[�ܽ�o�0wFZ�⫰TMdmJ}����`��XX��/E8����NY�[En�%D�)f�N�ͫ���˟�B(+�>�ޫ���O�b@B\�&z�S���#�����љ�s���IM��j[��'{�p`|�Q���n⣯����[A����9�r����c��q��O�Н��?����������-0ۚ���L�zZx�|Py��vli�1�ۿ\��N�yU�J8��������rٔٳ��bR3Nf��P�o�ߐeWv��Y_TG�ĖY{����H�v)w�!��J7A�II1��(Z��*�w���:L�}OQ�v����R�4�(T�T��z��tM�{�$y���tD/Gk�Q(�/�*��4�P�v|v�y<����HP*�����w�>���1��Ɉ|N�й<�>y���u?�@ELI�́x�;��Яp(�Ν^%�z�%�ZSI
�x9�5� �Ys�g^ٕ�7�l�ix���a�1C4��q�E_>��)��~��*10n�jU�k
IKi{�7^�W`w1�������`�hs�8�kb`Dy�[<��N�E�kѳ������c��]��M����e��)f�n![�,7��>Wvҍ�)�&5Ox����N`KH��	��6�/DirUj��v^�t��D7�����2'�&��$�ZC�N�ʈr+4Dr�g����)��K��{i/E�����eO������K�S��x]d�7��a')1)lą� ̵���@-�6�����eX˨�����N^�����v����Gc��$�v��s�H�眹b��q��@��{��҅'���RM_�����wL%c\xo5$��[���a�@�ܠ傸���l��@P�E�T62��V�)� Q��-�O~1�_ekBD�Mo�u	�*��(���b� �S-Y2Ze��A�
A�W�w�}:
?��mcD**��	�"�XX?l�E2���8$!B#tS!��u��K�������ڙ����*^(�^S�o?��>�l"ݳ�.��W/�y-���1ȸI��6���J@�6�`��BɝZ��*��%�Et�Ctu�.O����2# Fh�p���+_���8 �7��04��4�v�U�_(m����9~aQ�`��#W�̒wo��z��m�v�db����1� �GZ�M����W���tci��}�$L�Y��������������j��TR�Z�]�L���ֺY��N��h5�䥟^��iU_��9�~rm�u,����J�M.���y����/k��+��N�t7��T��O���x{CF�Ay|��ZUmA��*EU��e�3�&r�5�?�w�g2�p~�h�����qn}�|�\��G���9���m�'�����[��_ǎ���t����ʩ$�:�{�T����v�4�~T�*�j�Z:(E-f�ަC���d��U<�7��}q�C�ֽ��r�R��4bJ��_�nr�Z���d�O�7b��WK�u�S��''~Fm;b��[-����Og�f��S$t9,a66��,� X��#�WOR���ۦ�߃�d�G�i�?��(Ѯ��� 6���f^]n�rg|��5�!:V�A�8p�~�񅐰Y��%�o˒��ώ�� �$�%�%���A̾�h���W�VvR�y��}��媐R.}��e�<<?�dvT
�;��һ�A p����\�,@!4R"���aL!i��K_�2�[y�8�F¾�����?p`�x����̹H�/�T9'�֜���~9�" ����R��.�����ne��r�y�T@���eU{�����4%g���]��Ŵ5���ǝ��ʛa�#�vw_Z�+u���geF�j�;��W�]��������iV�[!us}XM�$�qE,�|{Q��q\�b�LA��Ex�&�V�cUĶj�(8׫W��qφ���W�~�o�tw�%��i�\�;Q�XA�B�!Y T�H�4޽7|{<e�f��U៟zJ�jS�x��3]���}�5l��sNgnԱ"��ɧ�$lP?�N��U�5=d��-�s5�1�>�����u��b_�c$��|�B�`LW���#o��qsW�Ԉ1����}Sĕ��C���&�]�)�@%z3xS�&�<�Ѿ�6���=��Ԩe2h	�7�+im\�~�=�:u�?e��s�t-�C%�[�#����h�7KMD�.4����[������W~�j�u�;�	�@���7�|E�4�e�0>���Sro��S�Ѓ嘋����|N�aB|�{�X-�������~Y25����Q�#��"{���B������
=.���{ӑ;;n���HdN�f����	3�yb̻W2
�q��Q��I~-$�MLK@�4�k�5����Vֵ�(��k�����B�`�\T�G|��s�,\Q��\U��V����P��CI�z	\�����{�u��{��m|�(o|��h��[e��Ad�J]�}jQ��~3�����D&ߖ�	Q��p��ox�?�A">��Cr��	��;�5LqS�i�&O9�I��A��'�A7&n��-�7X�V�AV��g'���U_��U\SHC䈭���u�-�Ϳ�4'�&��>Z���kwp;��E���p)�k�p�St7����o�C�~uf�+�4�z�QL�w.|����V�	��.��Yv��_�$'=*�0�R!�װ�HR�=
Q2R��媀8�Rr�l��`ufs���M!c�>i<n��h6Ewk�i6I���1�l8@#P'����U���ٚ��+�ۭO�������b:_�*�Nf6�� �8�/���]��z�N'zh�ލ�8'$Ym�ۧ�S|���	N� ha�Dc���y��ne�8#$��X�0����X���`�Bc̞ EWc�����q�ؼU�i�}�|?�X�P�O_��8�eK[�liF���,�>lK���p��ŮL!ҙ��Y�"�������2�%��˄���hg�]4
>l��P������u���Y+&�@�#���fPL��S���-����)US|�����7@����¬ª%@�o��a��?�e����D��"��`�5�ߔƸ"w�=vi�&(�=���cd����:$�#�^c�K���|X�xQU�+��@��dJ: �Aq�1±qxa���.FL�'��c�-?Ȫ8`~^ꖏt�����N���mzp�	���E��;d��u$WCD��������c�	�Hց���2������e8
�R�f41�˪o���C�zy��Q��}�����ה�͒M}��R�.��GN��(�F�Д�^u��|����VZ� ��˹�:,k|Ө�O0��5����+����D��v���������y�=r�1/����d �?;�:D
�p��^�JjS&�Dه&�;��3�5�T��t�~���?�@,�4��Gg�O���T9�6%>|�
\A��E��c&����d�c;�=$�����h� !	�n��^J�������Tǋ���.�d?���̉'�v���_>R�kU�T�wl���R��B=��?B9�|rG�`:9�B�O۶�L�el�e���:&r[�|�
ŅC�����,y2FJ',�ݰf2�XB,r���%�¸�K�5@������^mP^P#ǻy��o�5=*�˙�%Ϥ��A��>��dnim'���}b'4�h�%�
��1찇LSyBs�u�Ū�{����*�(����"#ݦ*,�t��;�� ��I7�
�W&�]�A�|s�x��3\1��Ꚏ�����Z#����7u�ygB3v*K�Ǯ�{�P}c[$��q2"عue��$E$Yf8�&��:��5bu�}N`P�?�@�����A��bS�%b<�	���N+��
�����
8�9@̊)'�_EE��:�	���G���Vz�%�(ڒ\l����@��	he,-?���ö�`���T.#|T�E+�(����@���b�3|Q�l���%D�RrX7{��]OA�#�MA:\Vɿ+�߾~e�Kw�{��:_4U��n9�����-<��p߄H(�T�#��D�=���O���:�;US�0t-;���bًD�k���F��Jp(��R.����8��U4R�KF��9�m�H�.���D�v�_�Fk��R�ĩD�6���f��u�7n׳�xO�_;	?��y�?v=$��ic�������c E�*��w����
����2j�^�Z0���Wvs �[�l,�]��6^.�ˋ����<J�Xb���[G�6��YT�݆�/��� a�<hjQ��L�5;�#nv�5�y*��f���e���:�����le��f�H���&#d�P��keoϩ�ߒ��$EԔp���>K��@g۫w_]7C?��<r<�˕�7F��܉e���@��9Ko�=��JP���-�OM�bx����ɦXS�pc"F�+!�Ҝ�	f�j�Bv&�uv=l�|��O}�y[݌����$
�;17�D�E5�m�؟h�)�!�ڋי�k�.?x�P@�bO��T8̋���9���-{!�RXv����2${���l��&��ĚX<DN���27���,�v�d����Z�#=���ɀ��s]�����k�
��8^Jsx����1|lv��% ��\�|�����&�w���e:F��S�2�$��.o���H�/���}��e-��6"-UZO4U�#K1�QN�ʬ@�
���iH_l+�ՠ�LW�e����5j0̎[�<��":��b�;8�/���-[/_W�����7�!vů��s�?�A~7�yP�\�xua���	��d���UW,~0<aG7���98��
�܏6��Ǧ�01-�3��hܘC��'cL��?��8g��k��;�N�na�u���@��E.|`A��5^EMtw��������ad���a<lC��$C����A=�����������M���h��IMz�ޢ�Q��Iϔ�A6�6�AbD�;Ym8���0�R����Ε��N����ZQ�yl���M`��ԤxrQr�_�a(�N�Y�=� k�9������1�iO@� j]���b�aP�Dh�<[ҡy�\.�T�'��K�$�/���+M�R�m��)��V/[�~�{�@iN+������^̴�_��c� �\�8�2ve�?��"8tq�@���WCz�0Fz�9�W���"�y��;�35��{��I�����S�j`O�n#��6�V������c3��W��R���t�V�j������@�:���i.B9zTm�JT�̀�}@�!�[,`�JWe�,�a�վI{��� ����6�^͚XJd�mC�UOhI�1:����!�Ek&��j��)[��X.�$|?�M�0���s��eU.�_f�J{�̋}JHX�6ɍ�������n��\
�oӑ��F���m��79��r��º%^�v��w�ާ}��{�X�P|bm���͎��|ݶί [0�ᴢ*m�'�q��J�o�Y�.��WT�u��"� F��t5���Ɵ\^>ǻ�3��E��~�,&\	���wl����m�b'�ЀA���YŜH�c��;j���!���my�+œ6�2޻V<P<��+U:	��@<�Έ�m�f������/|%����;�R��{:b54�ԕO)`��!:�k�R8:B�[۟j�1�V/*�M�l��L����T�F �o�F����5�����ޙ0�ز��7�n�<u��Vl�D�)ȶ�n?u�mP0�ef�bj,Ay{��'䇑�Z�+�"���Mj�Y��H�0m5iݮ�&�y�(�%f�Z���Ho����|;1[2���O��K���e&�98~�̺�C��9��P
�����Jv!])���pu��mb_�� FU|�����U`�bNu�Xi�D@ӄ�X��?.����)7��VFq�/��/Ć�N�f�w�I1�G�$
��kGc$D�ʁ-�=�U+N�_e(t�y��o��~���ʜ�8��n��AO=\�ء�w�Xh����s�&����Q)��1y@�����?�3�.��8��3��	 uN� �[p����ѥ��R��?VeE��O��vnm�5A�nڄ��ﰍqQ��^�8��?/�n���C���~�/r�)�C3��Eo$'ύ����o΃��Ͷ)�x�SP
��E���q�s�����1���}9���ѝ�m��ם�ȧ�"���I`b"ǧ��{�`8t�b;^7r�/����}LM`薘�������F�AfƖLOS�,p�o�|_`W�:㼺���Z��a�ۻ`�!1L_��!p�??87A�DC<d�4� �o�_.ʬ�ҿ���\��ߡlc�NJިu�s���[���?���X����uT�]N���7�g�%��A{�~���p̈́a�c�搃�CzL�SG�o��U�.j��I�c'�&��H���f���Dw��;S�.� Vs�P�
�7�L���nm-�?F�)T��p7�]]j!;#���?�1�DQ|��F֍�a�Y�ӕ�.�$=��M��;�-�8P)�g�Voq���{�?+��a}U��.�וh]��1@!�)C���3)���ֻXе��Me�s.�c�����1G1�yH���J�vS���\).�SG����P}x'�"�|��4�m�2�z+����L3���$��uvD d�洰Y����ۮɚ	3���\�.�g`���>����Ό]����rO7�HGriG�i��hD�J�� ȽOK������
��*�I�r�����{�%V��W��']�o�[~	��Gp�0��9���>�5~���8���gR�V�
��a�U���E�E);Uǜ�����r<��Bw�%S���Yt�b-.��2x�L�J������ƒZ��1�Y$:�����XRӻ�Q��;�R:r����|Ů�����ʶ��ǫ�7��8ں�v��Ou���w���Bv*v-��+��7� ��p�
&>��oR1��$u]�).M��A�f���V�!�H�!Y��'�V���μ������O�J1�����$�NƷQ=q�S�q3C�I�Vӝ��n�� ���p<K�U��ga��D#��ic�Ro2S''O&���
�/�t����2%E���`c�#�x#Ş��zo�<�"q�q��{G$^x�E��kq���L����TyYo	֞����d��p������js7Gd�����Ib�l���-|h�ӵ�-�e9/9��Q��E fc"b"�B"�R�7e�����P��	A���v@
�Y(# �2E!ݐ����n��䖳#[�U����&� �t'p��#�Y��ey�z�����y����X�L{�A�;;)&ّ�T��a���:��Ct�?��@��
��s��js{�5�D����:����U"\Mx	�n���?j�1�9)A�ݦ�HbM��R���K�~�  \c6;^��,]��uV�d�І<��o:�y�欠�4�@T}X�����k���=g�c��~�{�[����^�驹����!��5 �.h	;c2d�ْ���yh��i1�<���b|Cu�E�*؆
�e��X�ٔ�>m�V"�y�����T���Cv�L�e��I��2V���$�)iO�+�M�:��w�3.�挮?��h�宊t6V=��-�^.t�?���O�wE�V��=�HDsгf����T�f�/`ᇞ��u5��v��[���O� �'���s��/IAҫ��X)༡ٽ�\2���k��VV����N���E���9)�uN��C��պ����r�$�qDS���r�m�P>��Ͱ�O�{Ȕc��] �=���̳���7�ث[B��O��"؈�} �&e,c�?w���"\����߱��W���C;��]��\?Su�Z���D�w����@�D{�"�$���k�/s;H�[EA�4�>7A~���V�/	�9��%����Y�n�l���s�ߑ����OOW:�?�.���Z1�u4���"e�c�Wk����H:�/|l�j6ܟ?�QQ�N{50�/��44�SGozD�|��uq���fޖs$�ѽY]��s۔���>%��ЫV�6�l�%�N''����~%&���S�0e�+%`%t"B|�p�������]�}��NU;*>+�0��\9��Ҙ���._�Z֭�I뻖�cE~� �3�lȕq�Jk��p���#��s%�ݙ�u��X�dN�����E�� �-��������q�:�����R_d$� �\��|#�ؔ1�c�+]���[- �����OaO-@'������g�~��nZ�����GS~��sC"�	Սy0�3�%v%PmG�Qv������(��A�	���wLm�[$��9��Z�o�Еl��� ���׻��i�l�m]vL\;��z8>�+c�5O����xy���k�� �}q1{���1z}�A���`	�� ���4�����0q�.�^1Y����}���y,�	!���]X�� DU�J���1�p�R�n3���Ų#�pG�pWH��evZt�#+j���N����
:$���670f�7��(+Uu�'<��v=۳���v^�Ԃ�=mS8�� ���g��j�9#Z�] �7���F�g_�"���_
P��z�c$S8��R�1S�5MW�ǡ�G�Q�..(t��o�YU�u9_��w�b�`��ݺr��Z��Џ�c_Sv���S�h��	 \k���xtIi$�C��V��'K���i�g��cH��1���Fm���՚��j���8���Z����Ɋe��:e��{��ih��̢7V����@H�"���� /���`�#�2����LY٬�?~h=�w��Q�o�QXڒ<W�߫����-e�R����{��7y,���|^�F���MG�XD]~�� A��á{�#$"bޠ�}CJ����� �8�{�����`u������5-%��K��g�
���4
���M�2��W�f48�1�����}w��&%\�
v�aF�#W:5�
S���/y?y՘�a܏`�b+>fHKӕ(���TOm� O �������c-���a`V�0�z����+�3�����זz���v�T�6ʆVvѲ&_��0���Q1d	�.!�]����� }}��{�1/� �`>w���������/�q@�;���.���i�ȿzQޯq��0��wG����k������M�h�PvI��=M��H��Eqi�� h��%Bg8Ͻ�X����6�k�)���h�g^�n�˒s�S��������U�"'������#�0��A
���q2��/NH?�~�Wҥ�S��Iƨ��ѢA����c:|(�G����(�3Ҝ5�$�Ҵ�@�f:t��/���m��1��u�̨�e+Ţ,$�c�#?�Y~�;�*��'C���1��cf�L,5[��u���.�I��*h��_���m��@�|���m�q�s����flMi��a�H Ԯr
��$
����Br�����R���}C]VF��90ų��eC�R�@r���ɀ���^�eEV�@症�T�����8$�Ҭ��B�������T����@-���/��=>2܌M�#��1����tH��R.�)#�R�����r��m�,�lD���_��7➌��C���%2*�:g󡭁C�˕��=c`v��XӃ��[o��f��s;4Z��Yvl�^��gz3��i�%t|E�kV��3�x�I$���^�D-uhi���b>�ʷ�<H1"�z<E�t������.v���9��{��v��h(���c�\�������钕S������P�g�[C�	�ċԬ3zi�����3����D���h�Ì/cR�I���}�q��� .I�ek^Hy�ĲF1s��Q����@���CMZ�ˏA�Z~�&)����.,����E�$]
�u}k�8Ħ5�~W�����ݘ��`wDX�l7�Vx�I��1��.�ǆ��_ޑ�꒠_���8Nøb��;HM\�n�Lz}��=wc�'m�*��iBV��|r6.��6�!2����ټ��1�aW R�=�^�������&<"7�F�R�BqjZ��m ]�����&�_E�d�e��!��ȃ�z��(Yk�A\T�V]U�Q�[p1�A�^6Em��&�Ԯ��D�a���	���^%�L�L�,�\��:eF���,��63���&.��ɵ��:Y�jL��[�}��v�ڦV��������v�-"x6a����0�W"��
�
]��r�kA��	�t�v҄ޠK�i<�����6 �#(�h�3d���>P�w�ʤЗčHt=�!����]�1/�냛�*�o3�S���޾E��y
d�{�تz��@2��YZk2��G8�_D(��/��QԬ����g\OdmB�x����c�O��ҖdA���/3f0R�ځn��V��y<�f�V*�I��q�p`�`����W������u(�͆yQL,E���<��@������_�"1���&�nP*���(�}�|�`b��@�2�����W~�����u�͏A�*��1�7�'u�n��xG�Ҟ�2"+���E����m�S-��;�˴�eAa�f�o�?vhL�YO�gQ�i#n�ei�tD3
x5j�is�����&7�[���ʗ�w���7����u_���Y�"����j�r� �F��b�z�e����s<�ߛ���/�"S��~	�W�{����I����j�DL0&�XѬ��+U)�3�v�Y�,G��y�5ܼt@}5�l�	����|N1IQ�w������d� ��@�#�/�� x[ʹ�^v��Ì�pŐ'�n�h� �-���U�A�o]�ҸZZL4?�s��N=
�Z��h[���sGe�eZ2�E�h=�5$�`.=�Վ��煑��u~$�a ���De�f:��s#�y5!pHU�O"$M�$6c����R��(^��_=2A0<��!i�nC�E�µؒ�/���������ONr���w< HC܅,����-x7�T�G�����@��_���U^q�vC]^��Og�����Ƌ_�����?�-�+/rq	��oN���zo�|��vp�$ ��ƅ�.V�ƴ,ϫ����$��o�	���Z�r�9�ȱu�Y?,��<3��I�n
���?)	{ĒZ�/@���k����p��W�ţG$c!5��i��'��j�U�&�"�rCAL�c�����k�T�c"I�ېn�!Yo)W!�d�����Vu^9X���ٳ�}��f�q��jT8�)���ih���u�xZ�{�@��k���@-%+L���{x�'�nӆ��뵛N�k1���l�\��LvV)��q�P{�~�Iv���'t=!f��b�a�)&��Ƨɸ̯P*�UMFCαyYN+��U>Jr��M���V����?L;��,���"Q��ʨ��ӭ�=�WVH2�}��ƙ�gՑQY8:{�̋�Z���O�*�t�y�=v7�׶� �U�o�+xv���$�n(�v��,V�<D�����U��]�b8l�
�U&�:��~tb�i�9�N���� k�I�~C"���hj�Up��-��t~���:�Ox�9��Ҏ�,�4I������+V��U��Sd7�oY�H�C��5-H+3��w��M�0�`�v�hZ4C��x���ʺ�y�tи�Rﷅ΍FD=�HR:��M�\b��8����1!s�gF��F<���M+}f�����D� X���w�֒|Eˬ&)���g��a��}�XH�Ђ;�|�p�@ݛ�kz���(�7�OA�a�5� ;���Լ�Y��]0{+jT��C�Ճ��s�0h��mWm+ P�\MW�"���X��t�+�h�f_�Re�+�^w�;iz<,�p��7�)�;w?Y|=/T����)�����nW@��Ϧ �դoлI�2Z,L��p���'���S�W��;�G֕7A�:���?�uǓC
#�ƀ<�W�}h"0��b<��T�)hV2���&��͞�Rk1ud���4f6�az���O�**^�����V���qT���1l�D�����F3��Il�)͈��?�ӎi1'��eq ������%9nҎ1T�l~��E-�A�޶�(�#h��(gD�G_���P�S��Jyp-E�e�[ٱa6���<|K��}<@�_�r˅�,ӿzt�40�|��j����������
�

�7U�����^�Sw_����nT�U��;E*U�
���e#��Z0�D���v��;g�A�L��$��{���g��F�����N��gD�0ⲥs�*ɡ��p��٦LIO��d�)}q�=0��jsGP�Hw�gt}���0��T��t�4:�S>e,�\n��Lz�a�� s��PY+�˴��;�r����D��k�x����ĕ)������ �zpn1�E�e�B^rڍ�@k���ͥ��a���kFEG	�H�G`Y]Q*��k-�Xjh�0po���#aQ=L��fM1I���M*jD��!Z�/6WQ��l��b7&+�p2$8��D�)V�WP��Ӓ��l��`�=yK���|+�}�t�	b��$ˋ{�>����ҧQ�~� )�2�X�K��X�^y�@A��������y֗5cА�n"�'+/�k�i"����d��[��nA^@��V�2%\�޴ �+�2�%X�X`����^�A�гΣ��8n�1{a�@-ҽ)�.ډ7�Q��p��(�a��|�j]�s�>�0�g';���Y6@�5������`S��v�R����䝚
�̒�#�����mV�=��_ڱ>�=Q1��_~.[z9�$y���0�-��l�|!�EX�y@Z�0q�A/�t�7��s���1��B��Fr.cE�s�zVX�{��:Ch�!n�qvGtpv�6G2[�M�Zr��O�Q�����'ՍG�&m�o��F���k�I�"���煚���X���F�E���F3@���Ƕ,��e}5��Ԭ��7�s��5B���	��-�ޘ�c+6`��CNH��Jǔ�$n�?zCDapG��j�[:Nzx|���4�XbP}4�XC�Yp�Z؍�3����٦,�c��ɶ�v>�Y�5j�3�?��T�Urg�d6�#Z2��MR�j⤿�=	�|O9@�[T}^��yw�[p��n�]�A+		f�<���T��ȷ�M�{}�(_�'������ V�\Z�{5#��ˋ7�m&B�' ��<�%eu�+���4hB�HH⚫ul�,/�AM��3�n{�>��B��ևUB�WsHW���A_�k���K�����CҐ�MŻ��f'm9,���>{��D\���pϕםנ�`Ћ�f+W"G�q`im�x6_�U�4���e�mG�<�Ƭ�Tl��`��ɷ,$�Ϥ���ϪQfv�-~S�Q�\Y�)gZ������!Q4曺�@���!�Udy��k9P�s�I>��� ��7u��x;�ow'�oz=c��y��":^X1Y�$�:+Yc��փ��7P@c{9���Q��}p#nc�)�x���A=�<LF6�r�r�g��쏥3��B���>��Y�F�q=��#�jF�6%�������A����8��}E�ɾG	��t)O*�/5Mڂ �M%I��(�%�^��eϸe��ns�5�PI�dU��We[�� ���>n�+��Z�΁tۮ����d�"2j�l�3�6J铒O=�@�Jj����ǈs3��c�'a�5�S�ć��bi��'^4t]�dHP�KN,��kk0^e��|@�U8w໒|M�F�`:*v#C�:����O����'�����/Z��g�~�R���f9�f�+�9���>�H�j�T�a��% ��c�bIr��O	U�>Q�]�E�Vý�+)��� �`���2�C,�������t*�̓��{���K��E��G��ac�ɋZ~��K&�lA��� �����@"���8���T��躀_������e9���[ ׂ���>�ҙ'Q霄��{�\z�F�6
LL�Y�V<�߳١R�Kj����ԭJ���o���vZ����ƫ:�7�@��^���;��O˳5G�y�����4�A���-�3�FbA���,[�I�c^��*2r�!cKu3���{�B���0�0w|���wR,L Ҁze������;�(�w�ЏSg���5�HX�>�
��'���hY�]�|`�NE&<Pq^)�3;�0�_��DX����H8P�0zpQ�J�%iN
����Q��قS{��4���v`G�8"�8��s}��[���T|ۙ�TYL)HB~��Ġ�7�]E6y�H;U�"���+i��=P5�>Z\=�z� �ݘQ�7w]�sD6k��?g��,���ҟk�����k`x�R{uJt�Ϗ��)��7\�r����$H�vf�@z�t\�x�P��������&�lF|��7n����z�B4SüwR!A�����,|�~-����+�b���1�l8 �g����\=������:�b���D��.�t���_��hH�RKl,�V���<q�Qq�JPup��������������oMj"%R��i���7�(F�����ġͿ�z�,�邵B�} ���.,�������F��z]_]ᨐ�^E��ص�� �I��[6�16�F��m�W�
i*�f4�%�vyZ�/�J�1���'��mj{1�0^����c�{$w�m�����3��ǥࢃ ��*���b�������h\�I��\QZ<+��G�i�Z�G�޵���^�3��5	3(vz���(�j)��x�T�_@y�ώ�!/�7=E䱍�8�L���연�tt.�;"��	S�Y��	�PX���{'�q^.t���c���8�#�Q~���'�%�Tr������:*&b�p�<R�a�ĩ%~~�K�)KS�-�:���"HĔ��nGA8T���� `L����_��WnE�8��~�"��m� ��f׼����Т��}��z7���@�i��XTU��ڱ��Fm�M�0�E;gY��$�.?�o�^p%I�Mct���(^�z��d#�V7&-,�"��/�ɸ����^ϱ��J�k6�^}�>3�z! ֬Ӥ���K,i��C���1ac�)SM�7e��w"��Ἂ?��dT��C ���h��F�Z��E� �_'¡��6������,����·"?���~�N߾�������3N�'/K�s?�i` ��]|�o�NZ֋&"�6Ǔ��!n[ik챞A40{�9���F��#܉�;�JPS0�87	<��)�B�iG�j�Üf�(l-�>]��(w������6n�a��Ԫ���h��	��ZY$����2�@Dc�\X%\�)6
3,6��Ƿ�N�5�P:�r4�!Pm��, 6�I�R�\8f�e���b�ҹ��yִ3u�T#�"@~��yg���/y�?��!϶-E/��E�{=c«L'����U}K0����}'�G�{�1��4{%ԏt`I�T�49�m$}|@��p�Hl,ZS+�\'QO��2ơd�s�����w�s'2`�yŽ�c��<��'�հ�K�E�P�(S�fy`@���̴�me�r�RikE,�Gv�
������$�}�V�� �+�U�#����fh��~]�A���-/+Ϟ>x�Ზ����K����UK�@F������h{�����m����"o��!��(��ٸ����ےN�o�@mxx��&�V CD1�n��{�;9�	 �ۙ����\s.�������h=��l����E���$49Fx�B�N��a��������ߧ�wqn��;����7M�sb��ȫ[J�˵��5A<�'��'a�j�#��2��+OЁ�)����Y���5�3�^2 q����8�z]�OӴptَ��Lu�b�䰨�7�"�s&����I$3n$h-�H����������ʷ� ��H�їG'i�oE��7�3x��劎+p�ڬ��St.�d�&� 8e��U�����T�x��<L���Нh.��/S�,�'N�����ߪ�-pe�����s4ՔZ7�^O֍�
�V��>r-P�um�!yMt��-���˰� K�R7���⎈o�|��"� ׳�\#g�i�5������9�<�蛗�D��F�YM�7�\x��W=�b��҆��N��("��𪎰5��Zp��}ʻ�*�E�:����A�Z���d��ɥi[�7J�0�lxu֠�}����<��������I��V��}/^t�9� w�u]����3�UA$����7䓘c�H�b���~v�Ι�m�u~���gc��	�<����:��$u39�-M(��U�����t RP��̱�&�K��$4��pK�d��+G(z���^#�z, e�M����G��fw�4{E�!yt
htɧ3m$�1B( ���*G���Mk�Q!�E�	�*F��'��5�l�.PI��r�u�+h��	(G]r�g1VAQ������!��-m�����szV�R8F�D�Vn��J��C��&m��U�}���*:'��z=%] �mZ0�s�F2K�)�>W��~~/OO��F���5��)q�p������V
$�q��ˑ6�����s�����(!M�����w�jC)������xQ�%��X����§�+�B�����r����Io�&�ъ>�8#�����oP�i/J�f��,�?�m�K�����-B�dcM�Ϟ9R�b�ü֩�*Q�yVDב��-ӯw���_�R��G���Gk0C���c�\È�4)��0�^Ӎ0���<E�/�`h�NP����L�&g/?�?�T*2�������E���W��d�hv��oRӮ���d��4��4�I��E�C�U8�h�����z3$��PcqfR������_��
�\�
�	!+gs]F���C�m���4vW&1�/�#��^d~�j�ta �\Q!���/�:�+]�����������
f:�bG�]}J���V(��p�������)�@*HiE�Σ{��K̅t��`E�\IŌ�s��N\�� IJ�J���c�?�]a�Iι..>�DHي�&��y�!�}l�E0���"�;�8����=�6,*�t/�%��x����瘾����Q��@F�bB���Mf��T<2�R8z�<'
q�K�A�MF�@��1Tj��/��R��6P�OG1
��n��T۞zJ]Z5�ș�:"oV[�U.A?֒�NӷɳQz`���e�<�}^��eR��O�x�YA���0�rt�< T���롌ԕ�Z�ݚ��V@V�fK�=T v��4�!f�5��c� =(�"{�,^�sZĳ��M�myY[�U�B��n���=�?(�D��_�Pf�݄կ�<�)lc� ��ed��ΛB%�#��~Peqc5N�BJ	Y�$G{ pw�j]nv	WFM�9⇩��Ey�R���}��K*$���[ �|�uPf� �~u��H�THhUZw�},SjB w�v�-���������$nf'}�}�����r=�pD*rԛ߰�%�]]��75�X9��2@Ēr[�C�n�T3֒q5?1hM
��TK�G�/�#t�ν�D���(S�G+1[���TG%�F �c@Wܖ�U�"�	ϝ��É'ٍ{�e����E%�>-��-ܘ�U��E�G�ڌt�g���1��_�ٕp6�G�W�o��+�t$�D�R���&��|`'-I����ٟ�l�~tP�F���Ҵ��XoE}7�#!'H�m��H	3j-6�(�I!�fr��?�a-�8z`B� ��S9~X��
l�)#\:��e�bй�(�bA����=��p�I���� �g��(�1�b+�H���D�SB��6|�����d���;�Ԣa�A&�Rf��H<�+G���
(泙���#�|��NK*��[�N <��T��h��Eu#8�ΰ��0�Cθc�s����5f%�f���^c�B����.����L�Җ�ҭ'�����ЅxTTß��.��6��[]+�l�����+j2>�cz���\+:-�@�xs��PFK��T��w8����5Q�3~ė��^��
���CEd��՗���'�>'z�U���X�仅�l���+I�	�Tf7���^M��c���D�#�S��J;�6r��8�^fV"�:���9�y�n��e�� ?Q|Gl�L�0�P�LuSA�O��-;K޼ɵ(���E�G̙�S9-9�������v�V�{�/S���c���AQ7�G���SP䑠�A��Fo!�>"����>��WzgV�"h,����q4�ϥ{���4A��A��/�0Z,���]BNPp±xNJ���ȘU��z{�z0(�f75��Ty�i(e�O�v C8�=$
ZN�SX�qm{��W���7��I�.U���0A�Q���~t�JV�nA0�{(������5A.�;O�/L��M���h<�Z��PyU��F VX��=�^`�P �7Bg}�ռ1%7ʕAg[�Tb�\�P$!���ٜ�4�!��OeZ�c�FԹe qY���VҜ�K.����z���\W8gў�v�7W�4�.���-���PPl�,Q�U<I!���%�r}k�j��b��߉B��Ĺ�7�K��f�(���:�_�S�����8+UH���I�x'��*�-���b�e�)s�	��g'��"{���zz����@��^���;L�'�h]ԉ{,uB�C���$8s�ao�G
?h�WҼ�Jȳ��:&���ف F�s6�[�>����
��ܭ�>�rP�O�kVD�c�k���:�ȟ;�@-(�]T� � oA$w _
i���g7(��G�RN�1Z�Yy^�(�2.�TL�±���O��j�%�ІAĎ���5x������&ų���Pe�й\\ZX�P�&�/�,^��=�p����4g�_�b�J�R�u)cY�*�w4|�h�����ؖFf,�שC��L�)�!��RſD�ޣ]<�o�n�t��������6�ʩ�J��杺���P�Y�j���I�i���zL�����(��2���r[����S$�� �f���Ez�}u��>�'OK
����@����/�ez&@�2	1ڥq�	�	����rp�}	��X�s��`�%*�ӳ|��N����4f_^���l)`U�6��w|��C�xFh����J�yĖ��j��!�l������O��69-#y�v������m�W&���L��F]���+�=�IѰ_�ӔK��$|�2�I��m�����椠�b1��ڙӧ�0�D|L]]��tb٭�~o\\��|?y�1ۀ�%�𕼝P���d�ݦ�$ɹhyb�P�G]�3��a�;��\�/<#��}_�3�O>�%#��ُT�1~rv���KPB�V�j�ꞓ�� >Z��>n�Ok���g.R7��W�m::8�NN>�[��o������c�`��
�U��'�̲�̕�ZRJ�xDڑ�o:���a�7J����-��ϙϣ&l)������K�b��
���<O�s�����[VT���N�$f�Ϻ�M%F|��ǈk��5.�c�H|c�]{�g�?��n�p��m��Z<Q�f�ʶxҹk%�#�P�n#��g�����$m&:�M��n��2�[z~��Ԝ��w����R�v����7Q�^bLw�9� �e���������1�1o�?�D~r�w7l�w*sô�$���-?�~~�~̨�*f�Yk{���У�y�	'�B�����	����s:���CC�y&J����Q�$�U���]p�C'+�gpU���8��P�"u�9�p�h��Xd���Y���v��L��o=����2cYU
��F��2th`�|�.��@M��a�Y����חҶ��[��k�JQdU���m +j�s��ԓ\��5�&�m�/� g�E�ِ;ד��L�&
�%���S=][�Z<l-A�O�V�Xu�U�OGE6��{ْKόѯp�L衦���Oq�����SYD�2#�U�*wi�!*���kN��1,���t�a.@p��Xׅ��V<���T@^����=��ny���m���8�����s5�7D$�C�j����:�:M���W�)�Pzz0�w���*n��G���7֠��^nim��;Td�[���m:�j	3��[,��'��'
�\�<�.�i�A�"u��g(K�Ⱥ�ޫ��qi@�E�6�[b����]�����ig4��LA�M�	l� N#�:hUh@a�P8�%�p�ju��ct��,'�>�p�T�=�����")�/�k����We���x�5�S�Kj(����f.GY:�V��ښWN*�܋���d�K
�FV�^�ͬwE_:}J��;���dd�b�d�\+��G;���lp�vy���׋�z�W��E'!3��=Ϭ��:���{^��=�E*�+�Ц?o�e�5����7�~��ֻ��l��X%X��@��i�~$��������Zg��aW���t&/����;E�q�q�}BI�~~��em��zϭ��ܦȅ`��5ܹJx���1֋"4�s�LjP2�$M"��"GY�L��������Bʈ����Ic�YzhF"� T��bp7�q�i%��W�h����|1E
jP`�7aUi�gU+�������y^�S�U�pwg��c�����������j�X�b��Q��n0]�*�D�j����pFk�P��4-ػ${D�o�Z�$0��ڥp@n�"�ߦ�i�C����j-��s�!��|���������lW��Qm���x���j���v� �}t���⧎������ba]٤'L1�rdw��[�����([_�ݢ��;e��%��W���|0#��g�^�42�cKy�u��,� E������	�1�[ֽV��ǋ]f��bC��7#����LL2��!��ԔWC��@M�pf����1�b�Z��'��`E4H�jG��{}���Q��@ �`ࢾ�"��ݨX0���!!�ӽ�;2�r�$��5:&���;����3#���,D!B��9D��-��"j��1\�����_��E���ii̲�˷��|��r��27���#�F�xGTi�	jz�aU5	j�p����V$ k �H�0�0�ٹC4����O�K�`�����S�1��~R���*x�1��U��Fg�R@��!���3�enFm��E����[�!��z�Z�jf�T�8Bʊ,�;�oe,��mS�� +�S�����g��^k�W�X�^ʤA0(�����
	��:��9��p�ӄ���ys���pO���-�5�+̍G��-~���Tbx����Z�������	2��P�=�é�%��	LR\�x繢1e��������"�$�M��٘
�z}�4#�He(�Ia&Q����ybE4�p�e���ON"�5���6WK��	asĉx�������兇��v�{���!��s��e�җ�K/��D�ŗ<���E��H�w����}�R���g:�/,9�%j��([�P���Y'h�W�5"	�F�h˷x��K�ۘ�
��Um��>4�^�棑̶�u�� orш]S��K+!��q��A/�Rd���Y�&)�mYã�(��"���#��NB�����6\�UF����
PEI)`���m��+�pUx�4��H_#����H=u�w�X���*�Q)�g�T�QT���>�<�Ѳ��kp�:&�|��\���X�Ú~:�a�#�Xfw
�*Ct����z�����<�i�M��Pt���K�J���K����Z'���z#/f�1Q�0� %m��r�+d(�' ��Y�B@��d����6�����[2Z�F�:�����#�(�(I5=��#<��E�BYz��-*�4 ���6?g������|�`a�5�S�_�kL7���M^�nI�10������~�~H��\���L��
^+�u�g5�fA=�N'�ƤdU�B�.Z�[EU�r;r�r�Q��
��\s�7������dA[9WX� ��9l�B�묤�+�V�L[�	�6����m�����|vflj�ZJ}���$� `H���4hGw��K��
80kw����}������w4%]"Ϫ�!sH.��1-�@vD�8_���IW�D��Uep�ʜƧ�?&$<�Q�1PB �*�BpA$Fy�����p�xɺ*A�2kvo5>�皰z~ �y�'-l�p�m�ُw|*�CF�;R�?֢��ѵ�c��Y���l'�r��|����B�ˁ~�i?�������F���@�`�B&rZF�v�@�dy\�}����"8�5�}�κ���0�/`nd@oE#R�Gm��-9�����p]���AH�i[B翘���P����5����u���	*Ht��95j��f3ǭ��znU"?�y����ւ� �<vC,�,:x��t�5��U�9�2��O�$�ܣ�}�c�)?'-��
i���e�ۡ�F���n���hϖ#�v����rv�Y)Ǝ^�AmG�P�����Y{�!vI�鑣&�s.���\��,o��� ̚O���,5��b�
:A\,�m�a�D�����^�*%��b�y� ��x(Q���7}s�Vk��$VDY�#Ǫ3��R��?Y^�}�����0|�nA3�uͳL�7�ytt�>G���ՈS��,uʔPs5uG� �m�t� ��T;��}�k��bz�nto�����
� T�tܘauZ���&I�}�;4�"kݼv�AWh��<��{ɂU�r<�:�Y�N�K\�rR��D�#�f20D��˨��7WO,���Ț���L����x���]�X4�eN��h�Y~fk�+I���� �0nQ|QI��HQ�q�Z�Kk��d
- ��Es�&��W����d��N�zٳl&9�0�Fz�Q!��� �E����5�s��~��^��W�Lrfq��xq��M/�9�ק-N	���QX+���ayW�����^r�l�W�"?��]\�Q�pnjÐ�U��uf|�9���s��Baە��9�$�4���n6(���c[����Z�E�n�܀����]N�O>g�#�=��/�{���%�z�򍇖	\�����0W�M���(���riS!;
�Ѯ3�l��E/zL��怀g�UwFp�IA+&�Lȼ�\��?/��W� �w��M�av_�[IH��a:J���<�WI���Y;�/E���xv�7Ѵշh�g<�s���@!�?Љ�}qG$��Y�&{O
U2v�>�f��9q���ޯiWǩ��>lF�Nu��� )�X�����2�`�`P�<��GFh�4v��UK 9��X%h���~��b���g������Q�-du7#L҇��q�����2E����01�:�S=�P���7��,�1b���{Q�0�'N4�{]�@��/.s�ҫ=�1R�%فs����Kc`��ם-�.�q���ҷ2TO�^��g�v��é����ez��5�|���_��jʮ��`N�\|I!L7�����}�
���?:M7�/�i�ږ�A�)9�_���7�֬Ӻ�O����h^$L��e�*n��o+�T���I}���lI��<Z��e�ȫYo�R���얱����Oo��Џ��zhŎ
���uv�.z.�
��5�E�ޯ���Y�C��։9}} �{�9�f$&�v�=6���٣#����M�{ �������k񤅄W����T}i�)���*�6�5�W����2��hq�7�(�rx�o�"���{������W�b:���5IK����2U4����#�\�G�#��V�"m��X��9�<��6,��Cn�R���s��W�������) T��ص=�ΐ��öK�K�ٖ6W8�Ԁ!�[ j��o��J	Rg�Jz�������}7:�ˌ�t�J	tθ�1�(.d���ro*�d�4��Xq��/���M߶L?�w-�����B��Qo�6���������
���{(&N7�w���+��g���U��~��R��� �Ǻ�=4�Ǭ��kؽ(;��~V�MړzX��Z:8�8��Sv	G�h&Sm���}��͋⤳�N��bM��+�I��J�z\�&����j��K��*졥���yY^�27�����i~�ٲG̮�{x�&z��wV�-���E���Mwc���EE�.��s��·��;P��Pփ���7V�R���M8*��wk���M�Hg�.��ʜ�{F��"�%�n =+Y^	{F�w9�uJWoo,�� U5;��q����8|��ҳ�a"Hq��WPh�ӆ~9���^��'2o�)�V='Uۨr`���L��v�1:�O� �![��:4��x.ӌ��W���N�P:g	}R�.�#�1eź3�t��6)=��F#�4J1����/�}+~V��7���AQJ~$:����i1C�����/X�����H�;��\%EfP�
J�.��t�����NE�a��Ơ��b�r�X���J��]���,]�v�&lh�o|e|��5Uib�/���K:G�F>��z狻��_��� �|ϟ�P��^'S��s�p� �3'�sB�����?�ʺ9[ y�^2�	jUn�0�L��� dy�bG�yJ�i=�R��l-h� JA	�i�� Qsв#�h�ؖh�=Ϗ��rAf�s�0ZM�]����1 A�:�)�҂�E�Ⱦ�?��>�
]\�t ~�e(輪�R���ڊ��������vY)���V�9�%)�+�����+�m�C�#҈�(ɡ8�?H�W��zWy+��sɤ�<�9�	EE6�
P'!�9&j������N�fSMA�����p63����M�]���+��[{j��衚���R�#eF�T%,�|l�����'�(W�6<B��Z�9��/|h���:���q����y�5c[7䂓9��`��d!�-�}��16aB����j���؎�����Eu%#~Piq�!bF\�芋O�C����,8k&;K>>�B\w���ܟ���1�H`����}�Z��|�@K��{�]_dN'�6��&n�	���M/R�C(�}��gA�mu�C���8��y-�_-�2��,���=*^ys���:���)*�Kf�������R�C N�_�{�5E����y���G��J����&]��q�#d{2=Hi]Å��~ueI�2gUZƖǕ���$ C����@�{-ەE5u�t*H#@{���S�W��6�3b��׶�e�0�F�F?��YC�4��{�ӥ˸��G�����@�~܁m��x��z6�}����U(��H@�Fn"��Z^������4L|��f��S���p��\h��fk�O������;ȑ��~?�k+	��S���:��'���;�lm��4hK���]�!���a�)�3h�����#pRJ�D'kz��o�椽����?6��ٸ�o���G�j{�ƈ�.Rᓰ!�zgX�N&Ԁ�u�Ņ�B�׸s�6|CgSS>ˋ���&�M�i!�%�+��w��M�jg�rv=�z=��u�)��j	���Jp�ŉ�2����zI�9"�?��3��
��jB����;��	/c��6\f�n�Xӥ�U�-��^l��#��M���#I��x
�_���T�9�B��<�K����R*�
V�v�K�9op*P*�SL�q�]�"��̧�R0@�_c�)�k�M���c@d~��ȀYkrY���$��<�����~�#��$%�w,���zʢ'X�t�T���Dק�=!b*��oݨ��D�G5!��� ����}c�9-� �tı
໾��,��a;0���D�+���$���0Jv�U_��ݷ�6C��ToP?Z}�B�_
Sϼ��i�������HZK�KA�(���@�$�
^	��8�@d���6o9�_@�:�#�sX�%�s�.�Z������Iԣw�#Q�����,�dq��Q��"�ʵ;$�{ʝ4C;�2u�h�?3�pR��~k�i�访0�f�&�Z�s$V��&�9��E6�ӆ&���L���y5r��Fv�;$��o�zͭ�6�������Wg�[v�����&� ��^����(���WH���@.�&@��Ix��\�7,�#-�Ej֋���5o��ٯ'�R<��P7�W��p�<&�x�8!cQw���a��G�M�P'�td�V����qQ\ �";��['y���?���
����/�e$m_$�K2I(�9�Ǝ�"S�8�M�g"���'�=BR��8�rO�	]c��W]��:y�^�pp� ��3��h��Acemq�Ё�җ?�݆p8�l���NH�Ɵ�|[�xr3v��N�Y�ڛMbPrJ��q&6��XL��8Z��#���zg�4է@�ӣ<�\G\$9I͊�:�,ww5b��,��F��E���?��Ph
��s|���I�58��_��+����A��Y��!+���h0��꼁�ˡ%V~�a�=�+D�Qe-���1V�� (��'�x�{)���8p���@2�6g��ۿ9�/���o�2tN�$�K�&F��;ꠘ�dft��/$cux�.�Q]t���ZlݵuǺ�@܎KD4�+�����8Z:(@5,���:��ㅁ���d���n�Q-��:�{O��ˌD�g�U�j��%���$�Ɲ|c��l�S� �F1N�1i/fKm�?��5۝R%^Yp0e��h{�k��Z��-0�\�`��]ٖd�8��Pۨd�D���<�;�uI'zcA��� ꡖ	��EN!�BN������?l]g��Z%�3�y��x��j�%:,!�qB&��5�d�����K�<�2�=)U�a\�;�46�{�$*��\%1�<�=�K����X~]�p���l	�IKNr���@&9^}��v���هEQ�f�̘���Q@Bv�C�/
0s����\7?h@�K�F���kW��Y�͎�V�ZC���Kә���'�1cR\�S���I�0�i\� �EtYG�\���k�ٶ-׀��P
�+�-��k���~�yt��z������Ye�|Pɨ�>��x�������4��Hq�q��!�#c{��������/�r�69Qꂷ
�"$����D��.���%���'��۝2��e�m`��[��/�D�AK����bkPs/�9�{�C���L�9����C�d����9�2V�n�0j�?D��������N�6�֩UuÛ��0���*U���`^�ޖ\���Ghu"{e<ݛ�1�u�{i��gJ��*]��AI��>���<����-�.x*5Cq��c�1RpT��T2�<mh��ŭ��1�����{���}�{`nϻr5F�"?K�6��%�_Z��s�t�ԛ��ׅ,�}i'�^8�4@-�?���@��t���i�����%�R���Xm����ޞ�$�����/���l�aU�Y+��	�]�7� ��@�j�?>�+���s�¡��J��s��iC�<��h��VU�u�CN�.�p:(1���}�`��T������C���m	�UV�_��:��d��~q��
��%�B��	� ��kDb���}֧�y	�5��X*+��.�!��e�w�-�I��Q��G���<! �ԓ2%��kZ �
����ܞ�!l��4�C+��v���X��39ìv~h	0~4�t���6 �Dc+��e���8�j��� f��s=m$SAH�e��z��ru87mǦ�n�%�$(:j~��K>C�.�j]8�Rb��o-���jՅ�׌�WgUb��]��"��@B��R��授�!ip���W�T�u"�����J�������a����C����I��R� McY�r���uG���_�Z�[���L��N0�I�60~�V�RA�{�P��v"l��H�A6AL �{�<�c��*�D����"ZԹQ�i��D���	����H���n�}��XM��Y� OeS����h0"}���;���cS��,}XH����O	��%d��48���M�M����l�����%ܺ��KM9���5�=����I�����G��eFwP�;�)�q�X
�ͅ3�y�G�E�tD��%�i0�VQ˧\q9��4.������j���vY��!C�	ZS#+R2"D1�Y����5$*?��6�C�Si�Q����Wѣ`\ ��n-;��W'^�.���)�H���}�I�e���*�R�UUD�E�ՠ&4�tNH�#��N[�[+"�^o�zlD�aVn
##8�/��K�6#�y%�O^����a=��HB*n�{ܐ⨗��m8���`��]�L)��Cq���{��`lO�5c�+�\��[&�t\g��%�\�ղo`-1#j.^�k��S2C� 7?�4K6Iѩ{/^�Fa�\��ѡ��0³$=3�m��g�t�x�����~n�"\ǈ�ZC��w��u�Tg�ϔ���h�M���Hf�A`�.R��x�5 ��b�ɀS������fڧc�X���f�/�_����쮯'���{�^O��W"�;�
��~F.C��� �Ic�I�n�t�1�C����W~-PY˞ �`x��ۥUDf!B�D���N�����A�^�@� ��ƨ�#�Ⱦ˹4}�T��:���&I�;r�,���zޱhset~� ��8���x�7�'��^p�܍�i(�ڊ҃���dD&�,�
���-����g@6�i5�Cْ�#������7),ǚ��q���
M��ݑM��=�P��WB~l�����#l;%�_��);�������31s3�i�\L�|%�ܧO޹�R{�5�_�k���|ų��~_���ޣ/"�+��KI`���}�����+q9�@6V��00���kE��򕘧*,��-`����T ���"gV�l��'N@��kn/cJ�i	W@�:�.��g��y���7�J8c�-?���1���W��V����(�;������{1����S�Y�y]O��x��J��Wb��Q=�h�Xo���;��a?C������XA*��6�Z���v�G�'��y�M�������o��rN,�,��g�}�ҟg��:.A��gaL�_�٩�/����n�t>w�5��aEZGe�g���;#%�SXzL�!cg��}9��Zr�z�o�AO�<q��i��z617�<�IL��^���.�]����S��2[�w���7�CF!����5���4��;�=�s���}�)&��v�������H@�uS�4+c�6?���Xx�F�P�|OЇb�Bi�ZBh��f��O<I؋	�N�ϒr a�ш��\�a�+���זq���
7A�-��`�����~^&Wg��'zT� E��7 ��\�p��*'��秞��^h�\,#��Y�֬u�.q�����_"˓2k�����VR�~�j�|`�y�m1�_O[�7yk<ߩ��RMF���)�K4�K�-d�kP9dC��ޓs}bZ�i�=`{�c^���`,ȯb���D����*F�m�������͆��/X �<���������!�$8_K�[�7ɶ���p�|���=�D�1����z���*�U�<�	N��Wu�WP�GǮ��-`�{�U�g�Ӆd�S���(�/*�v�}H���Ve���-���n5Bv)�:���@]��Xťn�wk�^���9�l�o�֮�����!5���/d�kE>�ֶ R^���������I&$��!�������d��*�Nb��D�0W���Ћa��w<fI�@3��y[���
#���*Q%���(����AҖ�Y�u��zN�>(:9h�{HmE�'0x�v�!p~�b���&�d���y"D�wSH�QɅ�A�8U�`+�j@Lc�Kd����A�JI��,�������<&�T%��r�=��O@nmi�ŋ�]������˭�����o��J§��δ����ؘ�[\%���3��(��u����o,�U�K�#̄(Ė��2>Z��۲1���E�_ᖵ�U>/� I!�z�Bi���f��+k�����@�i���w:��tlX~h�e��a�_%�&P�Y�*�9��ʼ���g�l��l�!���{FӉ����7!�ʙ
W��#^���e&������W����=�@��97�P�^�o�e�Y(�s�?$�~�.::,l�o �N�Y��Z�&
Iw�`��+'��_�n��V�qX�؉w;�1aݱ(4V�ݍ��d%ފ��;Xhb�^��yI��YYyOAם\F]D���	�U#�a�oaۏ}Q��U�n㝣�L��:Q�v�a�ŝZ�\�ε{&����=k��X�x;�<���ao��*HE:Q�qÆ��5-��!�$���D����R�)pY�ٽ�e���Dډ�&��z��Ǻ���\+��*�����?�rK5g�X�%E֐���>*#(�5� ;��E�$��M���Xs�U0�br�S�h4�$���!�����K�=��M��#���_'�g"{���O��@�Ȝ��aޔ��v���H�-�ՠz�=��j�Rl��s׫�x��&�7�ä�7��Za��s擥q*X���Lo��?F�(�����X�&|��f�Ba�E��VHIN2�Hֺ'K[y��6��SQ."Z+	�2���	���8!���6LZ�A�m8��n�݁�AG/s��	���]��bI�=F@I9{'"7�S�HM�?U�	��X��kA����h�q�������N����e�g&I��&�F�q�p��|���q���̱��<�Ae�f[�i�4|����
�?�1֯�y^ےa[o���i����X��E���j玜B�0��.�aD��3.����|8K/,T��~��?T�F�u3�������I����$ݕ���5�F���� ;�|:��.� �|R���ݹ�/��c�+A�k��$SWy��'j��a��TF.�ڎP�~y��F�tu�4�K�՜�N�7��r�:�d��M��f�Lfa\��a��V�l�+�4#��e��1;aS&.g2y٢v	�S�fY��v�[�=�l�9M��0��K��S�5�B�)�%�l6�ֿ-�}��&��?��<��>���L��<�*A��ԍy�"+ЎV��H��I�gl�e?r��$}�xL������N`�|���e�r�B��(��T�K}���U�x)�b�X�?0���GWA6�f�tWI�`�&�~���� *,���b��M%���w�N�����.ũO���S�`��H�%�S�����n��0�ˎ��T��_M��!�C!U�9�Y�c��%'�u�`)����rǹ5A���)y�ۮ!�k�gZ}�����b9���|ݍ�]���w�;��	����f8��Z�ZZ.*]]������1#���~�?�`
�y��@A����X�{oH�-A �S�B1����Q�_Ht�����=c|#��g���uQ�X��Ȉ��t�Y�љ��V0M�K��i�x��^���f�9��l�W+�1��.E���كU��fו�Ny�4VF-cw���']�$����K\j&����2b���H���^ZJeg�J<S)˄���p$�x��)�M�< C.+9�.T���
.Ї1Β ��a�m?�bS� �&:��6�15��y���`�@����cp�@���Ȇ"R�Ǟ���w��Q�g��C�j���d�$j{vl�gM�JM��N,��Nu�g΃]`����Z!�&�����7�K.�ă]C��*��� K]�|ӑ��-��-~�Ĳ��oFe3�Q$O�7ZE��$�;��f���J���p2�ģf?�~�M���h�b{���Rw(Ҫؕ���%�j؁�)�Hݒ���bA�CQ�Ì�x��&�2�(����;1�s�$du������Bu��.�&{}�%����p��B�]$�� 
�?=��q�iG���ă}>ڛ���,�{��L��|:�bjA�=y�<���YY,F}�c/C@�ýSIъ8����~�ت�N��9�>��3�����*����>��ڰ#����rʉ{6�/S�/Z�;0Sp ����6Yv�a;�g�B���(ag��ݦ;�.�ƩC<�k�A8mѦo��7�d�%}�i;��*�v��/�f=�E���|�Y����W	�!Ξ[ �7�.�}fq#�`��e�N�Z�g|���F^��T�VCy�+sDi9cp};:�y;�b/�ǔ [��p+� T4jL`��Գ���K!oy�Pi�\S$��#|əP�c�?Hېj�0-�T�pr.<��(��ы{i:5�`�Cd<l9�+��-���$��af�������S� a� �kȝaF��<�{��o��ZÝ�?S��\���>��+K?Kvg$�,�1�lW*�L�!�+����;�AR�d�)\`��ioF��A�߼	�s��\��^_SG(W��	�)T�$�!I�D�$%����4���@�Є4�Oo��,�v{C���>�Ӑ��R�m�]=�!�[��v�e͂�
�s��<�s�;�U@��o�g�� ��zfH�:Uԏ�C�h���1�F���Α�}���w�K�gH��@�����Vi��[�����&RC�4bg��[���H��*!���E멵p*�l��n��BKZ���%�::K��f	�˕j���xۤLh_�|B�f9C0!�jD]��sF���[N�F�xh�~"�x�{��8�H=���,XYv���x:����H��M�ɳ��#L�C{<����bC&�7��{Z���qQu]`Lp�j)Ö�6�L�t������h���)��v�}��.����ab�7��+��W����E��L������!��)�o�h�S:��?7!|*�� �E��DheK�=B�����xd@�q0=�(v��0�4q�%:���F�|���3]<����!�� �0�Ul/�-b��b�؎�̟^Zd�s�J{V�u���#�N�]5�i5��!D�q?JDz�"�Z��8�~JP�����@�}鶁IK�ﳭ�۳|s��d��/7>�����㚫�#r��8��D�㋓A��� �R;�U�[=d������ ���8U"�ڥZ�	g��M�:±�R�C[�ѭZiQ&Б�B5���r�7oO*�C��
�9�rR�`/ހ�s�PS�M�����J��#+��\���'��er�>�@D?�Ϳj�?ݳ��#dY��SIؗtxo�P�e�"�"�G��ɧ�k׀
69��ݷtLH�(n�1���;E�c�9K��"#�-M½|���w@��G����EJ4M/6EI��j�l3�»�R�`�ЈMAu&W���N�Q��X������Cd� 9|�fE�D����ri~�o
]�!���li��E>m��FUʷJ?(�g�I)DxYY1�U� �r�
�[�z{
w���Įӭ�#!���Wű�P�!�{>�f�!�>t2*�k��iш�Vj�v%>+�:�=(�k=X��+�ᆢ�:i�-��~����e7�mї��oF�(ǅL"`B�n�dݔ�Q����b�4�~o�����)�z>�,�O�i8b;.��7���LJ>&|��|�NG`���X�Yj�'&L�w'Yî޾��w�5�ZX֣��P,��ڦ�f���g{��R 8�3*=E���{A~��|�û^^��m�=o�;-���[@�NAGO'���sp�I�:��2�^�m���W*L�	'	8S���b��\�(����O�:�rh�P�����-y�������@�v��F�%~eN#/C��	Lw7
sd����Wg�_�����.xy��T麗��\���!���N@h�#s���N�R���^{�K�֐�x�i:�ƨ�!iP�<�a�y��!N�V|�N0gF�DS����~�n��"�1ʱ�Q�OK�-w����e_\��Pl����>!$^'A��)��/�Wx�]�"o�$�#��(Ǚ����%�Pi.Ӓ�J��Οl��4��j5�`��˯l�D�S���1l�����m�,�|s�wRg��� _-Mq=�L8lG��A{إqlhzGPZ}I݇ ���\(�i��nzTpk8�����zI�A�EZ����m%h�K�?�#�hM1t���5����/0;J@��O�B��d��i`�IN�7��������Gw����&��sG�
���Fu�,�	�S�7�X�L�O���6�����KMz�ip/f�/1�Ys����o��Fߺ� ّ����#ƛ���\�e] 3��I؋�T�<�ˊ���(�:Y�@縀K
�Y6�������7�%��+�����t�˄����,�+��>��b����va��g	��>.�G�4���ē~�H��X\xx_���Z���uȥ�B����@ �������w]	<�l��D�]��5�T8%�=��j���g��k�~g�1X���>p�
)���Ɇ8|$_�N�灠(�!��2DH�`2l��Ŷ��;J����_�b���`t��`4OG�_h�otX���,.��:e���f��К.�X�&ow��L��S� ����X��Ϊ1�<�����X+c���Ðج�jn,;6)E��<9D`��^W�9��#s���$�zSu�Y־279h��_
!�����3�Ɓz���!��������0�>\�Fk��bN暑�d�X�H�2�����m���K��3�C@�X���):�6��86��᠝ z��@P�Pgc���v4�Q�����G�5�����X$�Q�T����P+9�m*��hs�5E�S5KM��j?�b����/eFr�@��؈E������s�)ڍt<N�X��'�iH.��O"=R�aEe�e.��۹a0q�������ϫ�\l-luy8LX��D�X}�t��L�~�����X�Ќ��y&8R��7W��eRs^��2^�R���[�/�f��y�Y��6b(s
�b��ǰ\)���/���٢u�?4ф�KY�Ϣ\��6���,�}�����8��͜�,jo�'���<�w�܅�B�se�A݁�&�.Sk�/�s|X�,M.v�~d}X��E�$z�#T����ow�����O��0���o��ƈ^jadF��u��.!^�[�,���fv�}�Kڞ�B�Ś$������wa>���%�ix��W.�3�{ܡ[�+�.��eO�eŬ")�`Y�1��;s�8c�eqy�/L�ރA.Jttx�����M�SP̧b�!��DK�Go5�0ل�J�k���gԀ"�e����GHec� j�^��g&ǚ�/�p��;��|?�8m�N2�>*K�ֿX�f�=�7�ɜ�}Vnp�l�_v��b�I�$����=,�+֥1)n\�_o�+��ћS�A�a�J��_A8�Au�NM���S�[���K-~��M)"i�+}�Xm8�u��z+�3��-�t�f+�g2l�S4��u^�֨����{���2D�puL��>��,M��hBZa\m�����9�{9e�d �^��{6��a��j��3��}FX��RJ��M����xh=��4E��a�H���+���$�̾j���TV|�
�-Q濋�����A�T���q�ꛨl���)�RV�[��z)$��"��r5CL>��AXh��yޥ��G%��?�3u�����{)�iį������a���F�� Q�3��l��+�O �|�!����sݦ��Y񶒆*к��o�� RtNڜ��gԃu���P�{X=��H�L�5b!� �.t:s{�+7�ˡ$��n.v'�sZ�򶬝2YW_�E'q�~���|��,���/( ��y���D�=�Z��q�TM��4՟GX��{I�8��D���m�,�̱6DB�e�e���c�_��)��,J���H*�ҧ_g�d%1+�zG׷{�	[�����3�>(eÿ:
e�[n�|4����tΪ���w9硡K�[˕z�D����/��p���i��d�t~��o9=��M���������r|�i�Ku-��T���m����f�X\�3Xl�U� �9Z��t^[��$d�U�*�#�k�1���!��7:ӽ޺nQ�C_���ƃ�wSNx'�.��I�N�]5�"�_d�l�ˣ�;�B@�zᰖ�dю<�g�>e;3����k�׶~��͔H��
�O��3�n�
}K���]�{
�-�`��5��@uY����i@��[�Y�Y�Rn��vo�8��E�R"\��~V+삳�7iMs�Ϟ-��,�歔�v˯�h�c��E��|Sf㲴�������l=R�h��Z��������J��gp���90}(�S�;��C�3���ҷ����ҵ�oE�\�����M5���k喆4 rY�pp�4���z�v��A����Ɠc�;��]�6�J�v}���bQ��^���0��{Z31�w^��CH {6tF�|���ԛ+:�@ʨ���� ����FFhw�YFX ��4��&G*!��$}������łHu��U%*B��1	�m��uf���!I�u�鋬/LY����g;$�Q,k=����q�V�;*���N�sf��ْ*�q�H�2/v[�.3��mO�O�S��;�J^}��7P����f^}�L��)��͍�`�!��
�Ӣi���&��.YKA�jXXT�ef	� ��@Dt[����A՛���|b���Ƃ��Ez}�eZ�$(6<�M>®��rNیΗ����������}����k��
�p�ɤO�V�p-��"/Ꮥܹ� ������A�|�?��33K�҃`�s���dz�`� �Sנ�r�8�8D�MςP�}5��^v�c�T�M�wP�q3�}�Ly�Y�>�Du�1�:-��f�������J5��F�nhƺ��U�f��JR"FM ����nuK�X,׷"��+��0}Hr,�;E�� �5m�Y͘�1�(<ed�dn�v�cn#����F���C��E����%
S�Q�S�hR�ՖB��n4'#�!{�u��]��ͳ#0�zﵢ�����[K�	�Q��{�|���{5���Q��14ތ�������sf�� m�s?8��
�
}�+��,!	?%���ii��� M4�މ�%3Ȋ�$��\����m���[��] ��5�M"o������S������i8N�,A�,W�F�� 1>M@���Jw�8�Z߀����R���#m\�F�?ԏn���ф	��c�b��?���d��oo������cr�穇��J��
��~��J��!X��z�� �uB�c�!���5
̼z��+f7�ku���L~��7�.j��k�]K�6�c����w��l��ͫ�ý��H{��o �4k݂�&b��o�x���������5Z�L*���!�O���7�(]� ���Q6鵦����fX��,%2g�A�ӝX�hkS�u��Y7��7��>�$��
��YgN���r�p��N=�y�9|��l2ƼI%D�p�ml?߂�x}y���zLTt�cP��F���f�:�p�y�C|���@(��a�GB���~���6c/���]6��`ĵ����ty!@F��.0��1o�y|��z�FTLPܳs�V�~��r���s�|����9wи�?ѱ�?Q��K��WE����3 R�8O-���e?�%](g*];c�~�Eqj���p������˵	>J�#�AD����?i��OH��T}�E���P�X����a�6����2t}�?3K����F@6����������KnL�u��2u�>�T�h�얚��CȲ�@��6��H>�ۛ�L�5��Ee���x�� ��lbn�նq��&7��9���NJ�i��#(l�1��R�B���
��ok��<�>��S�C>w+����"���r�v$�u��N해�M0^�����m���e��h��4H�R�q&�����F����̸�";��k��u�b�PJ�T��T�ǾkW�l���������-�5
�Qf���?��%aF��wh�"F�Ma�V���]G�ų�3��������T��(g�$���O?��>OhK�bQ�����-�����r��1r���H�cq@�JA���y������i����.�:�����Cs��n�B�o��ND�J��b�i��*C�����\p�c!uj���?��:�5�t���7H;�I;e���"�o�$̴�VT�/�*�q�*G�g4�G�?[��*����S��d*k��?;!2�$�	NEΙ5�D���)��XM>s��6]����N��Z(Ǟ���'s������M��!��l�����y�x���κ��m���7���w��b���.QgT�����i����v���� !@�p�62?PB�**�ߐ/ݾy;�9Z��t����Eͳ���H5�����%��t���I]�)� ���G��j�5����NO�����b��b�71���9�|�
#g��솕d��0�x�(�� <���a�	����=�8L��u�"�k�ؠ=��j��)�2%�W�f�=����@EV/i�^A+�Bu,_9o�:MбZ�bcV�؏j��8��g��~m*��q��ւ��U���F5�Q�t�Z�1�tNR\p�F�o�<�d:�d��%fE�D�>�YVՠ�6x�AN4��;uݸn��������f�;�ݹ���K�g�c��%�2�!I�R4�⨔=���:T�j	M����{��P���&������1q��dwM���--lCu`�Y�N�k������'�+̃b��M��Gxp�#��q�z�m�u�L�v��:
�ɹ�y�����3��FI�K��)�U!Hu͜�*X�
�shU$���4��4\�>�Θ��c�+��t�\{oN����G9|��ZcxI<h5��)߉H���m�cq��dOZ]P_	�?��"�YKJv��FY���!�I1���_��_A�ӕHTw�#:Ν�D~��+��BNv�.Z.�h^��D���+�8O��xJ�bj�C���R�>�W��xEeu�c�=����l{\mt�HL�Gs����z:݊ńFa�uƔ�z�'�;����1�,ء��U�JR�������e4�~em�,��=D=�0G@��1�����ᛮǻ�~^�{t��|��Z <ԣ}���3�cX���y4��2X]�l]���:��cR"����^�(�����6��e�
[�er3v�q��|Y}���J~�[l2���񷩻��^=X�ٱ�u�1tfx�^°�F�G�ȈDS���s���<-�p\.�.�	zj>3���3�7Ko�4_M�p
��������ڋg�Y�i&�F&�r��f�=��b.3��Ǔ��q�D��T�Z֒ܚ��*�߁9��LFid����8��h��
������"��ߜ��K�KA�1Z"�R	�B5�Y����yQ��dxKv(I�9�+c	?u<Y�M�b#����8�0�N\@����0o�˥π��WC`8�����Y��/��4���nѸ�q=`�.�Y���$B�9Xc�!,�N���xd�����I�����"?����HG!�T� &�zw�����������"��z{v	��O�'�`��6�k���!,������.���}�,A,ϙ��=�,~=2���}B�i��bUͥ�*�1
e�����$ߛ���SY_FC9d��G<�WՇ���7�t������k���\��&�pʾ�Z�)7��������'��D��캦>Yk'7�+�ϐz�E��=��Y�$"���|�;�	Y)�V*�l�m�nbSP2��Z�̍r!X���2�BDMb�ٛ`�]\�m4nې�0�$��\|X��Yl������TQ,���Vc���V���:5�z�!<Vks�$�8�;�則S�ˋ� ��(�8��s���Hy��s���=���w���g5�~8��D~f�Tp��:&2,�U�%t�����r� C����Z<{��	F���[gcMR]go:�H{��K���������nJ�2��'�n �tb��4|�Os�&�>���a�̃��B�ML<���e�
�MI]1^1X���Ѵ�	�	Q�hߘ��O�t�F��ׁ�7:�ړ㊟������4��.�%P9
�W\.ZK�1Y'���h<�m2��B�l�Z�{�J>Rb±}��@aM,.o���\Va\d��K�0��H_�(z;v�9�N�`�����3�ϳ6�_�����d�1QG�k%�;4�"u4��{Ǵ�N�<�*;ӱ@-��怓9�T�l���&�J-se�
)�W�-����M��j����������M闕�cƆ���:T���8�-p^��I]m+R[���P�Ɔk��<��?����߼Xa�J�r3B�F���~�}QAuQ���i-	��p�̌���U�Sf���$���<�����)%�+��ف�8̢
;�p�L����>ĸ��٦�,�1M�ΰid�VJI�b��v�o̶�;�e"X8��b�A�5� �U4+Z�L��b��b�W����^�t�=X"���q�N5{?B}���`pC	���2\�Rx�Nl�W�8:p��,�����B I����%�ڍ�z�?����e�4����qw�F9l�Tkq��H�l��Q��hI]~��ST~�&�rE�Z�ʣ�v�Y[%�P������vV�������ڳN�o7�Y(�������tM�=H��a]T���C���v5F�Iw���a�[X�w�u,���e��W?���{8�4�3���pZOF՚]by���S)R��dp���b��	���ɇ�hb�Y�U�1��fE�V���0��i�gWj�G�ۂ���Y֕��\}��T-��,�É�)�09qɓ��m>���5�/�qݗ(�SѢO%�!]�B�|S>��:%µ��N�ު�ꮨ���n��V�R�Juw�uU�x��`���6D0�`Y�K�-�V�wl+yo�fOBV X�f��<j ҍ�&�}���ôg��Z&8ƻ�������n��O����D�j�g�b��eS�AO�r���N~���?��KK��6�҄��o@�D���J�_���Gm�2\'�u��h7�c�mh֬��b�D��j���⨷����j#�kԊ���S7c�b$I[�]��i酬��w2m�c� BuȢ|_�	01��U��x�l��'P܄��|ޒ�c={�4��r�7������=�8���T<�$i8�,Ƞ�˲C08s_ϓ?o���`��b8J�
2>��x���Ձ�@�
����QʴTCU����,��M��j��|�T�m���¤���6z���IK�nf��R�-"�h�4|c՚Γ	{*0:��x>����@U���U���U���<9��Yyؒ��n�N	�� {@I��0}h����9�0v�J��ť���E�󂣮�x��&)��E��Oq��֖�K�5X��S��A��hfɱaP�Y�*�#~Ũ's�9,�]�b�Y��H�>��s �y9���/��v���Z7��Y����3G����f�5ݎ.Ѩ��m+��z��(���V�����to��W�=ݼ�O��isN�B�����\W/T|������4o������ �Z�����w���x] K#^����gZWq���at��j[�&ڂk�.=Y�QV.Rr����Zg*<�`XCO�*8�t6w��u��� �;��o���u��{��������c��Ƒ!̠��3oq������X�)c�O_��C��R����Ң?�4<4�:s�/Z�RNn��=��~�.�Gs0���A�����]����(���{��*�B�9� Di�?��@�Y���	�(
��b&��Rcٳ�?~��M�̓-m�V�*��J%k~��"T<sb���-s��
n�$�nj��y2G��	0����\e�1�ɫI�I��5^��h��[Ð:�ĝ
/_'E��*��< '��%s�h�K�k�� ��VnG���Ǣ��;R,F�.��%�n
O�*N�� tA�sx�;�r���#�>���u�A@ o_8�>>�PV�s��FasN{waM���y�9�%�zr�j@��	C�q���#HKdΙi.'4>s�V�n"iUO"p���p��N<$8Yl��X������c��H�[E�-�O[{�f�����}�ov������)VLB��:=-�W�`�4̞�bW�)x�G���e?4��%x����َ��|�Y�'��r�?y��J��p+8_&�#��&�V�WHى�Ո�6�gGD�<N:A6B쐛z���x��迥�[�E+?�ŋ������+�*��`Y�G:^�|v;��*���!���h#^��־XB.~��0���k�����M##�R�@J}̓�t6�H�t>/�����M;��|�?��O�#�w����<&i$~�=�)�Ic �����"	`5�{�V���H�%E�m���hȃ�I���V�k/��>��,5�JKJM�|�	q`$0�JlVa���ƆCG���y��
e\��Hm��k���z�dyl�]R�No.�y�z���o�YD��q-q�f��=�j\��i�������B�,���RC<"��D5�&��_c`�C�)x�<�F�-9M����Z(H$��jU,��_.G�r�ު��8^�j�Fk]��FeQ۲t�^����Xۦ���lu��{�<y�;�Tz=u��oћ�����!�۷���׺��a���Ԭ�����x���|Y=G���[�e�#�Y��-����A7֫���/j�(�+�ԯ�հ����Cf��c���0��������!(���s�p_W��Uɱͨ_s�ߞj� ���.+ϩ��J�b���|Ķ$�G�Y�'��_�;Ӝ��˰;�w��"��@��Yq�B���=�Q��RV=5����=��8S����l�K�r�l�yB�:���,�)-&#��_�fn\W���T4��[D)��u�B6�y�?�~���:��`���)#��ju4M���Ud�����ߑ�ך�=�jT�H`���)x�9��R���I��֭��IbeO\k�����#�Ru��dl��w�Hj|�N�Q�|s���"t��uE�
��H3��8�Ͽ�f��V�/���a�S��bӢ_0�����(�mX�zc�!��6U�;Y���� i���)%\b.��%�:3�.R�cor�;��o���Ϟ��.�v6� ��n��>nё�T|-��g��R:��9b���%U� c�!� 2K�Ǚ{Qj�f�	y�ir��>v?ւLM4'F�1�d��F���i��Qk����$Tg0�#��z7��&�guR�<<�2��&��^a[�����Pr5��X�+h�n�~�U1�ԯ1O�ʊ%�WN�X���K$�0cr8�%GAL���� �l�.)����mK�M�+ҸR��2�u�s�Y�s9����,�-�垍$Q�Aj�<T�?� ~%��\0�w K����7���Λ�#ښ����7�o�������G��Ȣ������"��6��W�¸����}��O���`����&S�m䌇S	S�����;mCVQs�~�0��� ��N;�a��ى��Խ�.��/0�>z�`����0�4^e�'������m�ⲹ~� �o�-�sжΫk8�P�L�\�TI������n��`���v��I�w�|2��ڧ��q=R9Ybϼ<��,��D��|�4�9a�PթYn�ٛ]n���з����v�ۈ�9�BJ�7e5� %[�]S�2���>�5��s�G/e� �N~���Ɩ��/[.��η���Hv�� �|;|CM���v�!Z���� ���*�e�z.�3�Y��؏�SG<�ΪMj��3>��>}��u�'w|�-O7�� �1ʔ<}�b�'���5v�X�!��#�i�I���z��:�=V29'�S}.����uI�z����A ��އЏ��f�!��K��+�w����Xj_a�7���Y??Z��9
�A�� �o4A\���,�t�����+��k[�D΍�y���[�w�,'�a��� �R|-Bמz�Яeq��~��t��$�w]� kc\�CL�A(����{�	#}(�i�������.
<��pY�;�;�H���@=���g͵,c����������<ό��8�l{��Ol��
3������@������ �@�Ƙ���"I���;))�K�-Z��#�Y!���<��C�G�{	I~gD�!H�LS����8��Ʀu�;-��ِLck	~�������i������3�O�$�c_���B�j���#�x����_ ���,ϕ�땚�*�I�暎$s�D��#M�x^�od$Ļ�ŊI=z��yܽ�7کX�������0�юl��-X!�e��Lh8�\2<,\��[dZ��E=�ߪ�Y��f5������R"���xM���ԁ�㍧~�ˣѯb�WvI�L-u�������w���;iP�k�/d�v��+�U7zy&Pr���,�"���-�5=U��~�C�t���42�B	��?2Q���=�T�\dPd��v��\H�>_��8��I`�w�H,���\\Ě��nTkX�Py�r���uOӪ'���
M�C=D����1=i�?�vҕf�g���
��3��zBa��CM��'�(�L�U�L;~�4+Y�ub�[s5���R�q�1���-8��J)n1�Z� Bt\�	��(`*̷!�UI�f3@���!h��n�
2W[�d�j9_�*����V��������e.@����� 8*zo���Ug���FA�������gI}a9�����E���Z(�9��f��ڙ]{	8�xm渡��5������=�$���0� ���x&]�U�3�j�*�8����JU0s�}�V�0+��@�A#�E��fe��Y�Ҩ`ԼI�$�oB[���"酁�xuC�C��܏���W���^Q��n�m$��4�8�0;q�(��yDp.C6^W��(�_$Ъ�u�Z��U������l���=Y
�n�S%����H��&�[gSmI��c������l�[<d����1���J��swj�������^�?������S3�7NX?k��(m+��%֕�6w*��hV��+�*��襂Jw������x�;��/� }"�~��
�|���~���ܓ���̜�Lܣ7�����bM	��f=J���Fƫ9�q8�}I�ҦV� "���U���.��E�<d�x+���np�����%ߨ�ї����G�Xfe@�k�Z4m��P��JB�E
�$"?���]z�
(E2�O��U�_[�[�YR���g�n���l�Kba\��ip���C�%W<�S.�_{�Ӵ��5�d·�� �y����'��m��N1�����hc��=�#�2���?cC�9f���i�ٍv-���ߛm�TC�:Qc�ϸ	���W��cG���ÿ�j����\��?��=[r&т5�s~�߮0��E� ȯq��<$�6�[R���j���Qj���H�Z*�)�O�K��ܿd�)������X������M�wCT�Rm�>��� Z]
���4;;�QvT��@X��;Vx5ſ0�b
���`_� �Y�4J�Ec��sq���,�hᐵ�P�Z+ {�C��#�t���Q \�*���<}���W�X��d����!T/%�e���>�ۏ�*t��kw�G�{��3�S,����
���e���E���������}�Nq��w��]/n�Y�i,uZL���9��N*vX�}����B�-�WlO&쓯>�C���5��fGq	�计P�;���]��/��ѨS$����f�+���;!mK�ձ���v���UK��ɤM7¾�ӽ���ca��5�w�c}K0[���%C���e埘
��!jK7��q�*뮰ק5�H�"��=cZ23��R��h���������):�t��"1%��J��q�#���n�݅���U����n��x3�ݧn�9{��6�Xg�:n���+&<:��ô�x,�IFa�y���C�!H<-����&y9�H�3;t������7	�?��������؎����;��+�)
�4��@���x�m�Y��0�A��ct�.���'L���*������f�� �s���;�Kg�7���C��xE_|�WZ��7n~ҥT{��"=�d�
�%t�X����:�����=��:��^�[�}�v!.')H��`��"=	����.�l� qR�P��%�#�B?�<�B;�@9�Xe�.�yB�N�,�;v���m�=܄����djͪs.�s�hq��鹛�;���c��q�h*D�P�N���X8l{����7���c[��U&�A�x�-�i�A�g�$ѷ�^��P�E�GqL���#�>g��cU������/��G� D:�K#��H1mNu�v���d�:�	���з���'Ab��PO]���Yh �+�#aWD���񅝉��N��43$1�����l�h�|�j&	��c8ID���M�{��w#�fff,6����6�<=�	޶B#M��<(��ƿ`���c:9Z<�r��"	%�P/������=��?&ٝ�h_�!��b�~����z�"k�)��/����Y3)�yM�GY~����&�9q@�0�
Ұ����3�֟Vih����p_�y�ќ]�MXN�({���:��r��m��~�;���cR݉ʧNxz�-'}��^9?�֩9�%H������u�Ջ�`Ia�E�+�����<-�S��v���'������%�$���{��'J��VF�ሿ��GT��<��ؑ-�J_�.�����ܶa@��lS��� dh�0����t���!%# DzҢ�U���I��DG1�s����?dwuP�?o0�������C@��9=�B�Զ	S�������jߑ��f�~K���z\��:�y]���wvF��`�����)���>|O�/]������a�8e��ê-��m�J�v��,�knp��y!q�W�t��Uk>�����Am������}��
*L �z[P�0�т���L�������Ͻ�[h���Z��%=���Z�?���"�ej�)M�X+����]���Zml���y<���	��[�,0�C�J�������;EQ��S�:"l����A�j�r��4ᚅ�-�rIR���E6?��I��^����f�8����Z�8�;�C��	���c���I>���a,�
��\K�����l����1`9��4}��ܙ����b�E���юjˈ C�KU��T-��C6����jzz���a��ܪig%��=rMl:PB��0�n�T���s�⫿\�X��%NB�fF'{�BP}6P�L����29�J�`VT��G��ű�������f�:O�mٝ���z�P���\
Q��Sq3VQ�%#���S9�������w�\,�����U5�*��.��ރ.�׊��#�i#�"�q�M��p�F8Pڸ��]U`S����8���� L�i֭3�Ó%�/�㤘���?�%�\C��P�FA���S��Hr�w��*hN���4ե0P��n܌����ؐ>�N=u������1%��o�m�4���y����HI�W�ޔ�[�����J���lG�~�S"U+�=�����Ū�.�x��j��x���@���G�*�}hwj_Z��|�ug,�����j+x�U�=K󾭦���z�3KR��@{�j�BhBm����?���������+�X����+���B�bѴ�뼦�T�9�$�0X\@]ԝp�gi�����Q���;l�>�S]�1f�A�"t�O�x����~}�	�fr��X ��D�f	��e�� �9���5��+x�FP��s�NQ笃I� �@2�(D�����+V�吰�>���^<�WϺ��h8:=g�.��P��.�!�`���7&���?�e�Ù�
��2��S��4l�FA��B_���Noބ�E.����7�$s}��i��esۜ�/�O�A1�a�;L �E�p��,��p�D�V5!�<2�{���3&�ϟ��Ft^�Ƚ��p�ʭ�ٶ~�"�!d�BD��B�'�6D1�4�ȷɯ��r'���0�M;�R��j!$J��������E	�>!<HWG���r�a�h�0`��q� E������d��܊qW�h��43��B&�D���nځH�3���]}���Wk�y#�p�^&?�Ɛ2?U�H�S;	�M%��e�rO�3�~��x��('�*��T$B�~�N�pקu�U#|>�v����,�����������F�P�g+���:Čâ2\��z��T��D�m��~��G���|�
�X���d��D��lu����D�*�/��� ��VG��*p�!n�$�H�ג2���~��-1�0���/�.s���N_O����qag�(h$���D��O��J�C\m%3�E��O�͹W����9���Ia]2�����J4�9��g/�>!�tv��S�
�F�����ȇUW׍)7J��E��0����`V+�*@~s����S�H��EAp����L��Ipz��ޏ߼"�q؛���S-�jg���A���M3b2��&���?�d�?��C�5�@. �gVɉ��!u�N��o�a�3G�.�3��ʲ��j>Tw<�E���7�N��](Qً��B>ZƱ݂]��]��41K.L.b�l�xǪ���{0:}Iz��Ԅk,=��ʮau��Fe� Je�λ�~vf>�Ki>C�J�'$��"���K����5)%v�#P���S�`Z��0��*�>��E	���oL���6Q!
Q+��������_Ѹ�L�h�T��X�%w�^��Nl3b*ˢ�~�u�� �[��ʱK������>Q7��5/�u.�u̼Q��v���t��(�H{�	�Y��U�V厜p��P�9���	�����GO%�*���b��*r�b�v{Y���\�	��LԘ���,ץ?�*��F�{�K>d"?	;<QI:n4��>z�|���q���)|l�����t�bv�,4�Ȗ�Z�1�R��D�S�-�CB�m,��A�����{>Ec��%��<���=B�c_��q�H�q�>�����l'��F�N��+��\�,�����9Ⱥ�߀���쪪�K��Y�:���􂰨�Y{^��,�;������|~Jޖ2���H��R��d #�,��LiPM�"�v�֭rs�T5�/�l�����}+��������B|H��$k���l,��6J� �
�)�.�>�y�*CC�;���|�������y�t�"�F橶TG��JT��YGWç�3 +�&$%�fR��9)O�$|v5���d�G'��35L�<�G�3H�B� ����6�B��~aQ�j�&���r�:�b��fwmB6�]�h|���u_g�w<_Q�0`B%�M0�>��:��cʭ��wBhKZ��"ո#�Z#�|3]
����="��p�?z�V����<r�1��(^Ƿ�T����A!�Ğ�Y�wA�慻4}�Ԛ�ˁeN�X���O<,���w�T�}`�&�$�Y\� l�ejj9�p�Z�2��?��K�0���f߼$~�x�G��i!c���i�:���P���^���=������&�0|�5FE^��ax&B��jD��sP�Pk�6��1Zs	��s�b��Zm�a@4�2���Vj˫!7����z�� ��x�UZPeB���}��C}�2
NĵZC�i͋�T�����!k|���CA����0E��3xt%]�1���ȩ)~7�0�h��/:�}S?�dN)}1=��d:����N�!��Mf���h.��G�sWIj�&�q&��mtڐ֍�c���@'���n~�*����Ga��~��W5��Tgr$��`���wD6X+MӁ�\qs�)���4���X����3̞+^�b/�\�p��(%m���� �\�l�Ӻ���r6|��� �n��8+ڲe�As���y_�Xi�t;����Y���d�>|�p^8m��qǤ��*�{�yt���,ͣ��IQ�m��WG,�[��3dM.M}�-鱫�R]+�cdt5�^���"(�|�`�%ܖ5�.}�ά���`��I
�� K���--2�NB�7`׀�6�?��C�zkW���݃�O1����&3�k�1,8��Q���I�����u\�No�-RU�{Յ�Tn��Z�����O�Bk�:t�4����aVl'���CN#�w�зX�/(V�d�We2^bF�r���X�B�ǀu�P�#�'�l~$�Ir�7�g �uꎥIh~biUm��1�>�l��Ժ��������yfc��ҎYj}B���C������F��5��PB/����0����PW��+7�⛲�!��w�q�ݛa_X�~�ע<8�2P#��)��Tp��$S�E� u���]�d3W��r�l}��ƕ��������CvT����]Eo?�kA��	��T|V�o���䧁I ��<+�,,���7PPc�_@����!�;�W�O��ȷ� (@n��K�&�lR�rx��'J%����t�̐���͕�MW9p�n_Od޹��u�^<mW��%�Q�L<ռ�^]��{�4�R������΀N�6����Q���b����Q����U!�SX�X�������F�y��<��/��C`U���Tc�{��᭗ b���8h���Ɇ��q
��c.�h}��o_Fy���h1��AFF&��z�Y��R�z,���h�14"$�����;��<�eF��XR0k�p�5��m"r*�"��^|.�ѥ-[`�_�~�B�����>[�,ISo�G�֖������~x:7w/l~`�#
�}ag���g��#+������L�E������b����BfN�y00�AE$��IA��o�>�G��{��,6��`r���v�H9b��L *Z��ͱd]��q�3��k��䦿T���'���d�@+\I}��ll���nP��DH����"��Z��ZhF�W���=��b\�~B鞖u�1��=�,6a�9&�g�y��?ʂՂ�+���
�"�9`���0��)��ϑ�f*��?}�i���^�D�A����֪u{uZ3��gM7�R[����VՍ����v��=Ճ[Љ�ȓ�W+�Tus�b^�{��%����
u��М���I�:��> �>@�[�9������!��"�e��bU���V�$E ��~"D�xь��s^3�#���F�+7[�"��κ�]Et`g��ڑ���VuR�|k侄VbKV�UxM<`�'���uc��hH�=��b����X�X�Y�y�̬5l]
��d�#Ք���D��q+��3�n� 	Y���Z
��5�r�ɸ�ڣԄ+l]�"ʥ=��s[�%��L�5[���{S��	7��'HO*u��V\��vy$ aRal`�S�0�G�>x2D�X"V�9��k��wW�
��r�o��FJ`Ĺ�N٫���$0�1�D���X2�L2�\���c����|�z�k/.K���s6/	���w��!��u"?|�۝;�m�AlΗ�͓h`t�^_�E��#�""ކ���U�F��"n�)W\�R y�&M�x:сUα9�K)u{3>�yM�=Ĝ��F�ruw5xs ��+���gKx��n0K����
j��T��B��eM��e��ɷ�G:Q�:��!�a�{��!�C���64X�0��ڨ���j��)�^e��lV%��4�M%����|<bw��|5�d�=e���uR��!������#(�,K�v5h>St�g��+W=�/-�l>y�j禬4�/��؛79Q�7-��{��V
���Ū�JΟ+�Cы�26�;FO!x^���&dox�kZ�r7Liグ�^��Q��\�T&�^�A�c)�ڀ0�������i�<�2E�u���a�ĺ� �X����-�Jġ�D5��Z�/
A+���)Y�K����r���{�"b
)�yXyt+��E?�!H?4O��q��6K�	���o)���٣)a�6���mUe�Q���U��l�������ۛ�Ur�A��˂B	�N ���aM�!�=$�`��!��ܤ!�M"Z��J���Ӄ"��+�`�����S5�t�*kR{.�K.n3 7�:�R�,uڻwRr̷&Apo.gQ��{�d�7�{$ m[d?2����zㄲk�)[�"�6��H��ڷ�Ju��J�iD�e	a�YLe�C��<I�{�)���} ��Ns2�q�'#��_���Rl�ϡ�;����zO�D��W�p��W��L=Q%5!��1|�c<��7��C�w�R���![̍@�����0�֮�_9]~���q���®��H{�ӵ�m��m��<F��ӂ�sH��M�~��)��=g�z�ڧ������e�S��"9�Kzg�{&Ӊ���+L�K���P5��{�`ѓO�xJ� $Z�P�:d#��O�d��=�ήE@=��*�V���7�I3�v� ?��E����>)?4�<G�ں�����JP���Π�W��[��a�L��6_ L���AC�[9�� l7�n�L"NUL��a}8���[2���M�:8�|	��Mm����xhc�A��f�;T�����$ ֒?��8�}��-ō$�g�hq+ Y�,
9<� f�57`�QڡU�t^)o%t�oN����?r�h��jȁ��D��#�0���[E_�8�]��z�(5$B�<7z,\�GO.��W��Ȯޜ��t�6o��X!�� *�i@%�9��ጎX{�yk4I���[T顩�W�Ӡ�3�+B��d���%>���Z<w"dy)7�C��<��y1�Ӥ�ij�[^ge�
��x�J_e�� 
����t�<ݒX�A������ʥ:e�%_�x��_��'����«$]�Q�� ���%�j��m�nU�^��߄s���v�avi�EE�T�u@Ur�ΝGn��Bl^i�^Uk�=�����l:���VWV���(!N��/n6�xbGA<��Р�}��E���ky3h��s?��g�xo��0����
�B�h����4�R�-��� G���v؃c�Go���sჰ�eĩk�����眓_�Ex�j�Wuk�Q*.q�o�w��w+�l�)�Kns�S(3@w�nJ��U�,��5wM�%�]��T�W5���� �D<y�8%�`�sU�t��̳�VνTV����I�j������G?	R#����O�"Z%A�:��F�\���\���&BO�7/�jב-@(���C`&�:Fu��^S�Ci��h�~���N�@gC����k����
���zƱ�=�%{<��M�}mh�yI|�ߌ�y�=<�|N|z<���u����}�W��2�����s�`�k���% o����k7u�W��ݸ��%#*�{&C�.g!�㓀 Y�d��?�VA,�� �Ix��!�q���^%����z�'���J�V�����h�0�59��p`�sC<�|W�a;U>p���_b�s)���&o:2ߚn���¥������N��q����S����sN؆8�i{g�6}�z���3q����@W�.���@%\G����+�����u��)���Js�۹l��r�L��F�FU��#���Ǻ2�5T#��Do��Q�
��Fe�u�E�p�)S��Tu4��:��+�B��e-6��漼_--'��1SZ���c{w��ϋy�l����Zm��a>����S�wc�ȭ�7�O�eo�`��#�������5��.�|\�~����,,�������b�|�O��a�����Qf�E�Uc�:T�呡�<�?�z�i��య(W,2y ��Fe�\�N��i�&�d>[����S���DSz'7�/�eY�T6 �q�H�U��ƚLU*��ޖR�އ����RJ$��A��tʈ�=�đ�B���gWg��|ݷ ӌ��t#��w�}\�4[�]I��2ie�.�_��c�w��q��u�+E��M?l�w��@OQ�'%���4V����"`|�T�4V�����9;�p��9�G�?�kol�~Nmd�����.Ν0�'}�Gۀ���*����Yk�}�	C��7|̡�}ɥѶ��hj̼���z`��N�� ��3�gB"���R�}	�Kg!��=��j�0�?�c���7����,H�5�Zi�K�K>�h��I	�.,�?�}qѦ�2])"�*d"9��9K*��(堼�/���]N���X�M}�|�`�z£K�Jɕ��E(�%|v�ϭ��ȑ�ʓ�_
�S�d�n�_�xE`��0M�/Z	N!d�HiȮ/֍bs^ѹw�������S7ok��CQI��̢���]�Lw���$'����Q$!���%`󷨡���b ��O9��΃s����$��,QA��K�w��>ʴ�@:0��i�p�.��#
&�	a�Q؏R�f�^�K��%W�؎�����<�5��L��Y뢽Ϻ�t�~�����o�l�� ��(p��0���~���ń9��˟8��َ�~�NH�K��H���dЗY�*������.��(�7v�pF+xE���� 	ۤs�g'C��!���`e噆�~�ې��Ǩ0�0���8���Z�>�:�n�
�D.���fNJt�S})VJ�a���[=��R�-�z���4ـ�I>	�}["b�"��}2�$0��/h3nZ������z�h�0