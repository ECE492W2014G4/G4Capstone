��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|p�n�Uˎ��|�-��P�W�l�#�nv� 0�΀�<���8ʕ��^��h���v���H� 
�>��,����v#���Vo�g7�fh���b���g���[Nx����+�Ĝg>�(�A=� d�<�؇�;����N˅������;]疥+��Ȇ�|�J��p�!c#�d��8�h8�R��"�sR�?/ﺷ�� ������ݛn���.Tp��;~[ ��#�'�1�����R���M���6�(LQd�B������� jòǮB��kQ�n����HM6z	�������:�F��1ز�KX8c��Q��K�
�������^�2a����<�4�o�$����� U�*�{��UD{c�V�������*���J�m��(��xJ�a������P$9s��Z$$~�/I]M�\.n5E���'��,�g�j�e��t�]{ت���-����v%Cȃ�q�_��L�^�o���V��O�}�Hs9��1�`���Χ�R: v�k�������R?�T��-v�h���Xn���f��� p���-�O�c>���ϯOg�k����Q�_�|KzW�/���;�
~qM�Vw�O�7/%ޓ����wwh���<G����O����m	*>
p`�N�Q�����?m�������53�}�17�iYy����V�����4�����p�4Q|B���K>�$��}��R������J�}�瑔t�,\�}+.��U<uY�ԓ�|4I�{YNN]�7���[�	]�|L@x�F��M�,p״�W���I#���cB���t$���K���,$דHn�gA�7�(�2�ui�l Y�&�q^��gx�z������c��2�>�5�s����z�Є����@�/�aA������V\�U��#��x
�E*��V']8��شv�tl,Ə����z�A1d�B
���n�:����SJ�p[�x3T��.�ul���3Q�_�&$��]!�1��hv�W�kJ����5����pۺc1��z������sRjL�\@oJEG��%;��� ~tY�$J</kDT�NȦ�2g��Q��]�1t}�5���s=���3�2�G��L��x޶Gࢾ��:���͎խ_�?�ٿE����c%�^J�=+/�e��O��ð�o	�ݭg�_����˓8�c5��X5�yV���e�g�ʲ�<U�QÊ���_�)�Ԃ	yk]emHs�	1.icR�V�K��ǥ>�YBi.����,�	��S<�j��	�˻ڍ���2tu��d�Zs,���g���>�Cۊ�~E�6�-r��n��X(f�
#�w8@�s,�%�-�����J��S�H���B��D�~�8���h��)R(R!˴�g�b	S{�T���k�~���:���ɫ�`�/�e���A�ı-��G1��dc,{������'�m`����os��eyQ]�/�S����<�[�����RXoBt���A_d�tʗ��#�w��� c��%�T��9yjN	A5�g�Z		w/�$�A�	��@m^�1�Q@[L�N�3��i� �g�N�#�ו"��y���&�/����[P�mOJ�
r-���S���3��k��R���	��W�܌A�� b±C��~>��5��7��&6�����+�
���+!#pMU��;KfG~E�Z�L�a�D��:�ı⽤�"a�j�o�͔z��� +��	�kY��'�Ml,a�?d�f.:�'�i���b�F����2�F6���4�9�)�쩎��6��,s��K��<��eȕu�x�7���b	��zq��}oXE2���C2M�:3-���l-~>Wj�x�<$:�u�r	ʺ���Q5dO��4�,�>Qd��W�5�ou�6��Ǩ*=B88%�gP�
�=&�P������x�!F�r5>{MA'��H���&I�Vb4K~ۘ��I!pM�nRt����l�>a�L����O.{��@�yR��|xh�JX;� S8��q��Z�������pO�2���vFHo��d}R��d/G.0p@��7�)$C��i��oO�M��p���pj9K��=?������DO�����U�-�[r{�8���L�a�+��V���"�A|����՞��{�����Ga����ndW��ּ����Bܖ�Civ1��Ll_h�el�/�X!([欁�ؚ���N������Wo�����0@Y�_�tQ�1D 2QC'Ҡg�w�����1-vA��>�\�p;���՚+U@���=��Da��[���nk7�p2��g�gF� 2֦<7����6�@&�ʋEL�^���:�p�C{���}YC9q(ڇ���@t�㠵z���y#*US���BԔ�c��������%�2���CHW�x�m�M���:��?�2����#>6��U�����Q�����G��G�1��#q2�z����R�r%�����I}�#� ��NY6�{aV����u�r��w��QV��yn�jvCiS��S��Y��?F����8G,r�f���>.���3WW�(�-nH;<�����!�H��m0�9�����,@�9	#e�@��f��00���r�-����p�9s^7�h�4#�yO�dG��1#}��W���������\ѝ���G����2��S�����0��vGA��3��-@��
1g�x�.oj�3Xz�S�&�h�]	�p���C����Zn#����id���z�N��h��Mj?�R�Pn�,�'����I�
e��3�@�;�#u�w��{J�jp�*#'(��&t�U'�\��t��O]LW_��}#����
N����ks�~=�=�GO2����`��z�e�������ؒ����G�7��9��=a,��I�Yw�{�x�}�����hQ���a흿8�\A2�vl�
��6�Z�5л����ߨ`��?Z�$���'��j��6Qw��'�:�
��ͦV���鴲l�� ��_3��	����pȼo��S�`���4(qnk��8RM�{H�Hxsk�|����-J(�^8��U��ڌ��1��6��|�v� ��o������,�Y����\`'\q�]ݕS�a���5���\Ώ���� _"t�t��G�@�<��R�)���Ճ��72.�%n"9�U�3B"І+�q�օe����)�,�'?�Mh�/H�����X���l��\��b	����:��/{\��"��%5������22E�X��
B�y�E�Q���Fb��[Iظ{�40�˝yk��n�R�����g��jZ���(��
r�RN���Y�m����'wz$nB��r1��?�Xv�خ�!��qtg>dx?C:~C+m����{�/u�.��x&�c[���y����y��Տ�6�'��C�{�U�E"�5<@\���J���[P��0�I��dP ��j稸�2pdx�l�P��A�d��{��L��o$���#ۡ��.d++�$���^���	��T��9eXe���"��gN�`�ә����p���MD��Eԃ��-ܠh�"uËE^T\�=f�G#�i_ybY��WC,3�}V��v�qثn�W��n����<,�k6uE'!Gm6bU��h��A�8�}���cA�]��2Y�-���SG��b�~��І:6H�❺GO��s >T�!\m�	��K��YH�6"ҹ}��Ń���#흉m�O��`�# �le�Q�&�?���w��X/.��jF[(ԯ5,G
���{+�����}% �~$oq��LL���?U^�����M��3�i1Ȋ�jl@�
4M_�J�e���I��n��"z2n {�^a��
�7��+�v��ayWn=��(Yzl,��]������ȫu��Dw��+?��DN�kݎ��hqIJ��[��@)��E�I�v�I�]��FE�ܻ���G4>�
�Cs�:
�����_��BL�K����{��&�-��֚<���3�dE�����>l$�
�w����t�/�~"H.����c�e�yi�� �_;�=�卵��_�G1�m;E{�̣��Qn�(��c��|:9�֢?��xUe8Kxs��>����:���Xc|w��qmH��-��"�:�t�������qРwAb��&��'�n֤=\ؘa!���R��ï�]��|�
�S�g t�n��?g���"���V�Ŏ@�\>�� /�Չ�ϻ�,8�ނ��cj�)1���<H~;���%�8�r�M�����L�ѣ!ȵY�b_XBs/�'`w-��a���||9|'�(r���mï��#3P�x��V��u�؎�<��T\�]ͤ��r��l3%&f�Cze
T@N<+i�:���!��8�"�(ִӂ>˅S�ŧ�J�O�>�t(s�
C�j����Τ��K�&����M��+���swsl�#��l��jl�4]h���p�-儑6�XBZ	�攊����7�O���S��X �*�h/Hr�j�#��y5�N-~��؆�mxHQ�+lL�t\p���)"�`�9��u���ߞ ��k[=n���/�� ��P灄J1���;��+%�,kN��'���=N�>'e���2{�Ӗ�w��OdA�JY�h�y��Lu/vk�`W�D||��[r�B+H^a��[λb9��U:��|ZL�t�f�y�&"P�DVNHr��n�n���,}X����ܯ�b�qJ}�Z
��˺�>d7GH�m�2s�z�S��L��|$��9����/���`�*��]���rx�&���<,���R�C��k�C��)�*�T��B�bA��\bM�u�p�p���n�|����QՌ��� �a�3�u���Ɔ

��y'��f��ԊL+�N4����+q�I�E#�g��[��sς)h��
����<�3W1`P�K4�Ln�����[R��7��6аp"�W[^�
���<0���J!3��wd6�;�&"[��uwid�*�^�w]����g�f�5��(�V}ٲ�3���[���Rʾ�E�cJ��'�w��)ˬ����w����/��.s�F�hjABg�H��Z���ʣ��g�l�l��Q�C�<��L5��6Y��1�J��2fe��%�FA�Y 3&>�\�c+�i=�>7��QD�i2��g��<+G�ac��K�6�]C��s��l��ES�T�xUK�rEF�	�k�9�!x44m�}E ^5�ø��t?�;-T��E�+z.x�t���AU�����ـ��b<�pGp-�%�FY��@�!A����|?��-2�EWw�K��U	dpЀg<�<|�X��Gٻ
s����l��x_���
x���2�-$$Lv����7��1\�kQ�B%g��Sv������ߌ�$,�;7�!�c�}&%:���+�<�7�pt|\>�⇣�����jQ�=|������4�Uձ�E륟�k�%���; �{�m�atI0�����Qs��\d�%�یw�j�X�^d0��M+|�=F�Y��q�%���#�?=j��)���j�e����U���f�"�(�D>I�Sa�_t���[��_ON+N�<�����	�7bOO�|8��b��e����,��53���=s�k�d�
|Z��,fM�Qec�qE&��]�k�k�&$�m5�:�R��`2Z�_Kb��������.,��Xj�E6 ux���N��p�53���bшd���
lS`��֔���/\�2�TZh[����t��h��qW#d6h�~�?��{��4��B޳��u��O?���8�I������{�c2]�N �������BU�7����ɂ(!P�Ѡ���A6]��_�[
a~l�]��q�U�m��B�f�]ñANa���,��y��_)����.��n�E�'l )�Wj
H��/l�ar���1���L��Rr�P�I��Y�[���\���Oڠ�pQ6�$�{G��?���u`�\�;q��`�d��Q��l9h��@${6���$�/t3���iWi�y.�Z�]}|#�_l+���@�.�d�M�(.<E�;������E������v�\��H|����Ž�"
���v ���t�2�oL*%��u7�ؑTP�A�tt�&�4�ٿ���o�;��_&�L��A6u�GP9�h���̧���۰�����{a��@A� ������D-u\.���L �n�
�p;��
���4���,@;��)�2���d0b���3Ս���.��=S�PI}��U�wrE{�]�r�Й��@H�!��@�ɛ��+������jSe���)ck�
Sp%����������x���JFR��nǗ�@Ɗ���p�+�|���/��n|B
`�tA�6},�}����A#@�q|���	z�Ϸ��]�u���ӓo��7, �>�{ڽ,/�����{�Mß2ea�M��Z�4�1P!f���O=�>�F�'ͫ���V(4�d�<L��ݭc�@,�0��eF��#��J��Q�9��oɲl�6{��h���&T	�j���(�ܳ�K6��g'�oѠI伃�K^;�_���E��7���ڮ�K���i�mzMX+<��u��L�v���%��W�ݴ����U��;ޖ�"�EM�t��cesi�hC���WGr�_G���X�M]�W���.���qhxF5r�Xe�066(T�����s��D���2���D�Y�!�TP�֪�I<1�j�j�R-'�U���0�rTK���Wt{����̷�	��V1�rHx4�]�չS�@�y(O��B��������O�8�����q�]m���u�c��������O����X�����K�`�"���Άmj1�6L�_P-����B�D=򳒗ԾA� �цg�����6�ޫ���N^���(M��-�sj��lB!�s�i7U�[kܤ>��C:���-]`#����l	h�
�dJ��*k{v%<��KB���=�����v�#��GIk����w]��c�H��H���i3�v0�8�Sx���x]�rU��	�{�;�G�t�K��,��SH��9��x0���:HO���J��>Ԕ��?��sAqv��hlg�����($eB�X?0�H�mΜ(-�i��h��|��ZX�ڴb,)�k`��5�D�|����������t�S�5jv�=�G<g7����6˙=ZC�y?�	���w�
�8�S y�'����je�n��"e�!�����Q����S=z�YY�V�-Ĩ���EH5p� DR:������v�'���/�/bR�b液����V)��o�3PD��>,O�I4��=i_��B�A��ԦQ�(�*$�$b|F͵���Z���F;��Y����'��N�q�1v�}�#c�ua�9%l}_��瞩�� �q���a�VQ#&d5�0~�#�����c��(ROY(ݰ(,��Rp!�j�{J̄db#)zZ��J��\q/��M�\t����f5��Ƣ{`��iy�����G���Eaث�c~o~�ź�{����(`�s���V��bm=w3�-?sV�бݬ� ���8��ŏ��8�p��/�D���1���&V��p����,��W��9_$2�Y��\�iZ��	}����rʉ_�.�
�V�MKT���,�x��Sf�*�w؊�����6�^3��f��p[��ӓ.�I07'���0C��%m�5�}{��oMY
l���Lh A9�9v�c����&������j�枒�W� A:l;ྣ|��~���_�8��g���:���J�5�13�WDV��.{���ڪX�0R��;e$sy�ڋ�|����5^4 d��z}&���;���U�(م���O�%挹�U*"w>�����w<��*G��A�Ww� P�5���4*���H�����`K#͚#wذ`�h����pL��e�u�0��Zh��H�j��!��q�E�H){X��&d���,�N�d�D�� Sn֬��?6�����"��2M�Gz�.=lp�����y"�UF����uS�|Wr@�2�����G�Y�_3�αOob�.�j_��S�zi�a���*��2����fc|�B�~�:6��64���
��L�Z�W�-���ܕ�[����=,��4�&��H����j>wX:?�¬^
UQ善z�d��x����#�.�W����'� >�nx)�!�/�	����2|vK=k��%(�SK�3s�+��]W�	�cCT=0�T� :���&���z��F�'��q��l�5����<P;�j�����h���~t�� F7�w7�;��L���R��چ��<W5���ܲ��HB�����9��6�+gh"u��P��~�0蹪K���1��B��,Wr-Ɣ�!�'X�ᔱ���s�@`����75
�qeUKc�f�h�MIu҈�>�qi��ʇI͟j��qO�����QJ����׭Z���3P-L��͞��	�@�L�xB5�z��c����$V3,.ȶ�I��:iA�k�\�+�>��$c�犬��L2oGW�\������5���F�;��'�j�9a4{t����0nj��O�߰gЫؽv6�z�]��渼Cg�t�o6Hn����DR�q��o���v �3�h�Ƙ���A^�L�nC��Vh���*�'�?n3�O��gɴ�F�U!�J>9{���C��J|�8r?h�L�f��`�	������}����yi�m�%��<-�S[B_�wQk
ǀUz���b�3�;>�@Q��{�8���2�f.ey���:��&u�y�'��c�t���[���gu��=�Eg��w�F6D�M�3��Q���=� ���V�*.}��:��c[!��	��ⵁ}{p Y���gz� J�W��q2�a�(%� ���~=�w��	ߺ?�����1ioQߧ,�o�t��e
�q��M$�q��_��ϝ�첩U_Τ����^{�"�)W�t*�D�VmF�:�_�J2*���_��d��|[.�s�� +��6s�L�1�)��8s+����v��D1d~��{��ph̜��%e��i�G�sњ��Y3��U��V�p�kS,�܅� [�#6O�?��r=��]�#w�5�A�Cs�_y�_�1�(�[ c�jP��Z2��j��?�f�,t7;}�n�y$�/e�!�aF�W��@<�+��$Eɼ�xNw���z�S=��'��G��S�8�id}n�K�_P����/xH[�atj!"���E�/�]��K"���sn��ԋ�vF:O>���a�ܶ� <f��fr6=�����iv��H3��J�i�K��#���Ã��l�dy-�_��9U(WnƼ�^|��`1;�-wt���&.�b���e�Y$fQUٟ����MJ��:��.c�*������n��^X󉥖HV��݂�^`���(^��{���Xy	yE$��+O�qi��s�K#V��%�3MŤ�.���K'��27�1��2�J/�K�[b8	{��TZ������$�{V�"�?v��|�Z/����f_+&�V-��N�mW���E��C��/� 5�Ð�7��*&��PS٧���Y*�qDbC����+�u��5��*{h���T vji�m!� ��go䱾�;Tf��7�~�-N-�M���zZ���*�!�uk�b�GFp�h'!=o���C�(����,ZS~�A����T>������%��I6,�^,��_h)��WPO�7~oH�bZp6iD
N`>��_m�ʰ������ow:>��=�ȷ׮��}����d������G`�9��w/4b�����([6������{/I������ �z.��H�Gl��`ё&	���t�뺻�TV5�3��u/;�qG ��u`��T>D|8���#�4�7�ݨU���](�՟:v���S*Ѣ�Q��0��Xg��S*�;I����Yq��TÄ�|<�.w�P��	��3�Q�dorz咊�o�	
�R^�9ܒ��3reR��	� ���u�H�.
ә/H�T�P����i{�����2䬻��Q�d����(H�Q�}�c�X{�� Ka����j�'�����gp��À�}����؛Cc� 1��?��v(��W)J�Y<��K�	�)�X����]�+EK���;�2D��1nq�U� c��?��B�㺓�i��:y ��(>?S=J@w��S��s
��䅤 JHc�9!�l��dZщ
�,�uO��8B��a&݉�ĭy<�RL��9N�#Lg� M�T�Ϟ�Y�����g@ՠ4��������
]���^b:͗�˄ތ21�n�lT�a���m�FM_<j0a�ӘZ�f�Ԍy��<耲��j�WY�t[g5���|O�3�)`ъ�Ï$�he���"�а��ga`Fx�oOr��씉{�5ij%�f���n��i�&��q��$䉩Y(/��,���7C�!�^�JHZ5EZ:�$[ឧ��<�7~m��O�f�:�m��o�m ����Rv�W7]|��h
����e�� ��l���Z���)hK��~Y�02.-�f/({�bp|�l�zNW�+Rb/B;���$p�p�I��x{�����g49,a[��^bf�X��Lï�P+?�?��x�[�U�^���;�r�Ց�)Y�9��"�����:��p�[�{H?j!�� E.���ͅ� �Р�M�3-���1~|����\J�Y=ԦsOk0e���~�1�y�o>�£���Q���a�Fi�<g�0ex�+X�C+�A�~N_Y�
�$q��(���W�7�o.
�����jo?�x.籂��!��9�R�F�ɒY|��AT����kΐj���q�#���@�0V�(����w"l�/���z%8���&�MU�!�(���w�\�jS�OmM4��8�xp��ғ�jl��� #H����Ŋ�ڌ��P?#�4i�9�j z�.oB`�E�W|l
������5Xͯ��z��(3��+2ʇ�u�	Ts�'�t
�c8v|ڗh��0�!��_��*(��Ta�ݝ�"T��&�O���2=SV���SO��AS��$J|6��R���.L9�,
@�����p�)��3puO{��u���ie�;���c��,��L�x��"�����f�&Cb�5�F��f��CmZ��$���5 ܌=�Ҷ��t�?2�@C�s��j���`w�r�������}�А��{�f��f4�'w+y����C4�X���b�1�阫í"sx:y0_��櫈3�5�
�)M��Ǜӥv	�g�Wk���	B!\��%�uj���/o�Y/�(�F��4�tA�Fu��a��f��r�Ru�9�Ҕ��i�w8SZN��>1z
EbX�����E�GiE���c�{! 7�b�4�t���X�נc.��:m9��X즆Ȩ������ݨ�`B���v�i�&D�j�ڠƁ�� ��˕��U�-ly�~����K0��o%�)�7��
�gP���g�6�6��o"�E�+��T�Ƭv�����F������n���4Bh Rl���u�ƻ����pӷ!����������u�C������9�Li�̱G,� q�k(�+���ב)!�0�ub�P���ߡN�%��Z��;f1��Vq@�E�ؖ��I��ܙ*����Z�� �n�{z7��=@����,�y���wlj[���w�f'��#X�]+2��3�C�@{��=������;�x������,�)���H���S�f����%��Ri��+�A�5ˤjRI٦���|��w����(zM^����|��6��7p�RZ��ja\��w��D �s%����N�6��o3�gLG�x��,�K2���D{����]%�	������G{��gܞ�-ꀌ��y(H�� V���������������z���jƴ�5�L�B��<�����+&ȣ�1�������[�[>��	��Q�a.����~��L)�� a;�Df�ą�ɵ�ȓdy7-='��#k�k��jL�a�Sg%�7�C�A� OE����s��x]�� pQ�<i�Ca?+��C���Q�O��~�ҡY֐��$�2��6!2h��+���@��#�*���W֭)�\یL9ʇ��u�j���$�5G�+b���v�m�ir�p���}4��:�0OE+��Cp�84+� 9[���8�q:���ս�$w��=��n5�>^P��~et�0�
�_�����qB��1.y�C���K���'��L8+̛GÐ3�+�B�$~�I�Γ��j��T荀��[g��k���#�e����X���XaR�2:1=Sp��<tCKG̋�Avھ��P^�T?M�J���ыS�	�ؽ���4�TJ�͵S�!�Sz���!S]y��w���fe�I������f)q:����s��R���Ś�����O
���#,��44H�FLĸ�VЫ���N��;��!��=���jĪ-�C6X�N�٩;j��U\"�D�l����*�G����s0��!v4st(ͮRX�g۬�&�{�����s�˴`��;�S����I��z���/�,޷�?��~ejtu�E�i�0J�rA
�k���{)~TY}�_h�6f���I�k�`\��Wf�gm��4ty/Y=�����'�Ouh�{�bѷ}�s�C)6�q��ݎ�Q�l��?h����_���v@�eD�֭�'X[\r���j�2MqCW
�]�������2Cd�]�٘N~�uF)w��܁�"9N�3;Js�\�ͥV癷:�uH;w�t���8?�����T�rmw{uS����U��1�FD�`<��}3����:�{��R]���t�UI�j��|#ݎ9.C~B�[��t�/G�#�J�blؗ�	�"c�0ٞ!����u(��v/�k�z���aL�͉�$����¨'ܳ��>K��sZgK��X� ����[ڈ��F�$?�[T�vE���P��H�2y0���y�ېت�����~r �u݄�FQ�[u�̤?R<vw�4B�T*�DAc�>�Ĕ�4��tP8M���C�}�����s*m8p�:�c�asE�'�e0��;]}�ٶs��$uq���"I�Wd`��$l�q�~}hE"ŋ��;�\)a�$����pd&Ζ �n�@��Y�w�5�_����6�ϕl=��<�m�vuV��_"��r���9��B}����:L݊޸�-��8�E��u{yb"����q��ϯ���I�B�v����h�\W~�uC�"��uTc�ɲP禂�X�n� �&v�}Lǥ��YtE;R�9��Ds�,zU?�.K�ϲ��aC=e���\�F}���"�޿є!V�H�6����n&0�d	S�̴Yb�m�`�t��X���퐕��3�G�+��F���q������i����}�ظ�,S�,��k�.�u��T�U���|����)�J���ER�J�Pΰjf�k�l$;w��ͳ�����엡0��yJ�Zw-��?uZ����o|O�*�@7� ��<�k�~�E	�& ����s�k4SښM#h$ɒ��u���1��u�|��GL����g�0i���Ԯ�0�?3��n)�y@�EsQg�1�Q�F�ӕ���^����^y,�Cy�pD�*�2t��1>ô�(�JDJ�L��W!
YG�$	���J�-w�Q��.W����W��6R����4�U��K��ц�D����d�9HW���\�D ���L�=V�N�Hfކ|:ƿz2��D,�VmQ��1�i��Ŀ�G�?x���73�09rT����/E�Mb\u���+�}����U>Q�^mg���B��:��-�U�b�?�/Q��"����#�m	�] �?��f���]���W^4�u3���:{;I�PfzۥG�'������V�`9�E�}Za�3Z8��J�3症�ٿ��Z��kV���f���5�q�yF��1yF#��A�D� 0	�t�0��U Wj�-��v%�����[[,UT'�j4)c�{�H����	Y#�I�7>[{.����q��Fdc�W������w��%c#�
��[!F@ _�~T�`�m��
wr4�#n�1F`��vN�R�0����<VI�C�l�s�a��&���f�x0$!��U�<߭������S�(��d�5(�w.3�H��UU�1,?���_����Ua�f�n��*zW�8s9�Ka:�Aq/(�������Q����W����d@�ժ���@�1Ɉ�t�x)[%Pʥ5�x����a*�B0�[�2�
��a�w]G�񀦪�!���3j:@F Jq@Q��w�v�H�+�B�z��|�M�6z|�Ҩt��0�{=ՌN�_Y��b���[�%M���b��O]NW���L�dx��(�� އc����7�ҟQO醚�"��j����B�邿L��G���e��槊p��h�'��j$E�Č��0�6��5���p(���7)��^� _���[yp��;E	��f����s�����H�m^1=z��XO��{O���S��c��@ ?�m��$2��W�r�ɶ(����O��\�ͣ��xV�D؟�WK��۾�.�q;���Tc}�Q@����0bK���=��pv}�%�� �Vl>�܁� ��,��h�󕛛������V.`����@':�tRﲴ㱤~<�0s_pF�71�l��x��_p��֮5��j��t��mx�:�(�.*h���rTY���Ե�:'j�������ǧ�*]��D���Jx��E�#�G��L$�f�������a�:��t�#�'���홟�.(���pc~�%��A톡N<G#j�q�ߋeb���c���/H���>��V���o$�y�`/5�Vv\���8�#= �|+d�~�bv��a��Kp\�ij?�չ�p�u7
6�i��[q�vk�!�"��Ģdͨ|}4�->���$������,��()�v'�
v{��}{�mX��d��9J�͓���
xX��۪��j8[c�B�5H���OI-i��w@=�ݣ�%�ﰻ���h{<P��1Pz�z�����5h����0C޸��/��N������:�d�p4p�� �����2(����m�����)��!B�h_�2��ʓl�+�jډ_�Aq�G�#�1g��Ce׾�a֋�҇b���z�
���_b�3䥃��.&����rЌ���O�|��1�&�QC��iH�X�ਔ�ʊ��/����J�*����FS���2�\M�`���/����)B�Ǜ�u�/-N\?j�cr$ Nt���.�T��Irt�H�)T���-O^9	�F�׳���/��UL�J�9D
��RԻO�_�e}ZĲ�KFg(����i$��ݰkW�\��>I�2��O��p�]��`�B<&~BfE�~��IynX�^c�3T��o��y�+3�q���:�ɔHuwl����czx{.�hC�}F$y�?���G��u\�X2���7��X>�ݩ�Ī.R���ݚ*%�!>��H�IE7 6�����z�T{�G����hb}M"��vN�vuV����K�x�f����-�r��#wR�
~�5�S��r��NT��θ�Sd�W�����?KJGO���{�u":�7����oX.M��дY�fu����9�xOEC�*�g��Ɉ�u�f���H59A��Rn�A<e�Ƀ������$r�r���u�A�b��-��Mn���[��%�]� ��T� ��X��]�sr�s�6�J��W����,��<��?k�uw�dz��O�-Sx���t�L�k�t|{[��Z6��}�/#F�#E�s�aƎ3�S�/��Tvc�=��ot�zT���S@6�L�A�~�A`:!�"|�f��V9�E�q�W�,�����X���*F)�]Ĕ�⿆� �Oo�Wr}� @���{���r�o���Gxi#��82C|@������67�ZY�����'{a�5m�TJD��.����c�1o9�\���/2��A�D��$	��(ݯ3��k}�I�ۣ�"6C�N�~u%3u����������c�dv	M�#鰥Zㆰ'�q�!/�!mB���v�� �5�'a������:��ߑ��l6`�ڤ����`�;�����V�ۑ/����1��?�S���y�૧������<z]��
�&����{8��rFP�G�O��dV����Ǹj0���1o�q�vz}�`>ˈ�m�7����("��T槧���Aoi��wƕ>�:���Ջ1z�bG>OGQQl��&eF����$5�q�/��� 0�>�/G/������{�Fuho�,�o�d>R�S���_�jVî7��nT�%S�Ɗ�ϭ+��(\ƍ<�O9�_�����t΃R������و�Ͳ����
���`�W#�;rL͡��������H^FX�J�����E�$�	�I�4�{�{X��#�HW�����obF3�c��n������!mE|�E����9�ؤ�Px�	�
Q�6r�׽2�T�i	%�T-R�( G�f��hP#��Rΰ#�����J�8L�ZY�������8�����k>���#ף��*���-�P���b�O�2���
˿ͻ?7H���(��.�R<�K�3�wJ�Y��:�,�h0[��(���������\���fl�����,򖬩�?$B��|Aځ`B��)����5��1y�v7�sM���F�x�
p�K2p��	�?�QJx凅5=����
��]��|Γ#���$�~��p�r�kB y��/�G�[Vv����qY�ǽ�A��c|<j�&����x�Q�ߞ�������MY[F��^�
�Sn��xk�カ@���tS�9�9����2�θ�"���k�O�C�=v�$@��|Bs��Vf.�:�n �ʫ�t3�CY!���w�{VW��}(,^.ʜ�d^$q�׃��Ig����?)#C�p�yn��Z�����������ԇPv������?�&�:gT���Y���.]������_��3y�u����D��rIN#O9/!(��r��pu��fr�����̘J��B�|寈�|ӳQ�||Z��ӏ/����&A@��b�IAub�3�B+��+ձR[��T;����
�{��n؝Z�R�t6�<�O����4J "�
R�,l���i1��CC��R�XcG\��P஫""-:7�U�s��1��y��v�N���Վ��"�:4�fu�6���2N��CЬQZ7#ĺh���^d�p��@�R{4$�נw��xЕ/%�qXM练֥&�ԫ��|v�x��TP(����E�h�ud]L��Dy���et���{�fTX�=��2���Ү�h"J�I���.�WX���'�Nܴ'�'�Q�/+��>�}-�Wj8Au�bi��<��]�*�7�Fs�<8_�a��JZm���X<"�ӵ!�p����tĝŞ2���X��x z��4�ҍ�5���ǳ��:Ѣ}I?W'���Spb���v��fH}�ƤM�~h�b���)�@�-�$l;��,V�\`�������]"����{�e���R�w͡�(7��M%O�o�.q����Ii	7#�GM�͌��b&�H66]�����^;&tO�֓��M�]�R��W}��.J�@�*�sW	��^)=��i���#��Ve��;�D���7>��t��M���̚ѱQ�D���Od�rNJƖv�Q��Ig�hۏط|6�6��s@�aMw�-�U�w��H��f�#ۀ�̹V
n�*ݺ�2V�#�a����X1�
.Or����Fs�����U��z#̮e,G�4���
�r"�O�KCV��Z�:B�Q���C�A� n��5�첍�u�E�#l`8���Bm> �W��, \O���n[Ͷ*:��ڗj9���,�]~g~~���Cl�h������p�Q��U�|��la��RG��җ&���������,�c��N�[���A�Y�;혴�u[w&�� �o�H$�2��o@���c9`l�	��T�L0KY�Q��-B���1����IM�����~;L����h�]��غUե(�Ԋ��%$�v�.�^G��� �վ
��w�p�X�.���
3�ֵ��C�,�bUm��mAhO�s�ŶR&�ס~�M+ɭ^���X�����"�Tu@�ua��.:q�z�s߆<�<1I�I,�}4u�n�;`i����Iȩ"�c��U�G��������5m����:�we�u"�fI�� �4]B�t8	����yTv��So�'��75��-�E}qK��e-~1U���z�b���,^l�& )��8�#��}��8�LaC��0@q�ɣl3������ZqV����t�$,���Q��Z�?��I�!/�rGhu���R��DF�5NR0\ag�'M�ҫ$л��M�5��>����q���Ba۷kr���i��q#�x��0�¦ִQs����=#�q"�Ԗ���=��Azy[�E�V��- ��r��ZDޭn�!O~��/�?L�Y�Uɽ����s��ȲZ�|uu���5$�'�$Mc4aۼ��q���~N��:uL�1�El�vf&��%��-��V���8�O{Q��LU	��#rL�в"��c�3xÃ	��k��9�B*?��0�N1 ����ު����,F����'��_��|>`:|�A2���	���w64���̬�~�����뀚C����9��ť����=�u��:a^U�WvW�egj����R�j�(��;�@����źE�wL�sM�&h����>��@�l�Ƞ����A�)<�:E�M���c�WH��g�����jD��y%��m�i�ǡ��G�	��\�&�\`�?��"~��.���T���T��;1�q�߁KU�G�F���]�t!g�õ��ȃ];@HĈt
!�k?���@Oo#[����H&������B|�lɒt^{��͘��N����ި���m�<SʛϱV�"<�"�j mv�o�7f��"xm���(ر��D@׃2�����A�:EH��&�Uo}�����7�wuP@�?a�����7%> ���� �{�GS˃f�E�n!�j�@4�W�A���@���:��TX����Ei��6�{3ȗ#���q����@��h<�)�	�K�r(c�$�!t
\�xu�_A$5��m8zeSI��P�<�� �����`�OM�Jk��j���q�[�����}��eotP��%D�{�e���ن!���N�yNw���;���W\Ď�X��v2hַ�=Ʀ�P��n)���C�f)�����o|�v�Dd�eo��XC�D��K]�߻�3�ݙZP��*cE�! !���B��n����� e%mt��4'�}4��s��&o7'w[l��'_���P��Qt��&�P"�8~6����]�w��	�F��f�+;b�U�)���i#:��D��R��ꉨ��H&�BP.����-Y�,O�	�Q�`)��ҟ�|�q�)�f�{�=�n�N�:.�4�D��P	-m�f����-�U�jKzC���Vݱ��J�Õ�P�2Ĝ�O�B!"�+���.Ieu�ZfY�+��Q^�ܸ���o>�/�����7�b��\�1<��E���8�>i(�����@q�0+˜���5z��j���p4�g��dLDv�7���C�����7d����N֊��T� jN4+Z�����,��^R�&�4�}|��8{(R?�p.LRf�
&�U���v���ֶ�:S��D�瓫�Bl"�n�+�o��t��'��u5/����Y�P�Y���8����aq#��6� �z���҆�O��8��Mq������h3�
¯Z���e~�L�SU�pf���h�z"\�Z�S�<��cٝ'G%��J[�
���i�)D5vۓ���c���'��ɛ ���S�:�1��	�4����QuT̷����Mt�+5=p%���"� àQ�fC�}��������؍��J��;i�)@�j`��r%�R6}�aU�{~RX�����:�-�z�cu?NE���·o�w��4����}X�ۅ ��[����GR��|��Ck������P�~FP�$��/0�әr?�����(�q哜 �2�Y8c��1�)���6����E�pS}>EPKB���'%&H\:�����2�'Ƿ7�?�GJl��LV�2H&OR��f>��P�0\!��s-\��Ɓ�^f
x���Jr1��>[���/QN\P8��(�R �k���.�d��c��-rvܯd*��$��9@�O-Y��4��;-�Ya��`��Bt�D���F�櫅/�,̷L���d�+���i��/
��=�k�+��ӛ7DZ��H��3=s�t���D�¤r��n�d�HYRR_K'_��@�Ǳx]����^���+��;�?+��;��6���e�`˄Ś'2�C�5���C�g�g-�n%�?������.�)f۷f�t�I���W{b|ӂ��(��L�g��4 K"@���S׾���"�Zfo<<��A$U=M�M��&��K�u�kn�a��-S��{y�0�<����F~v	����{��C�s�>gطʣ�UH�:�'��uE��6J�	Xk¹�H깿�#f�0����;[��^\�����0���2��7"���<8Q�8��H(�_���̩���Ȓ�f��j�X�0�7�?�r�a�eK�UG�I���(�u�L�|4=�K۝����5��\ւ��v԰���-ܣS��~rR^�����(��+�GG_�֞��l��}���+��[g)��}�z�da�׶���[�|sI�!\e���A�f�j�xz����B]��
��ð�Z�YҾ���0^D&w�]�=c*d�[�^H���$k�hvU�U��_Ƕ�Ug���7�xN)� b\��\���ۺb.i����R���*�9�{�~��iK!��"'��$�xμ�Q��Al-�8�k"��)t��ى�ybPop�}�o���ƴF
�9�\�$6��oDE����S o�%���bF�͖��B�,p\=7��y�	�~*���j(]6���C�����'�<4E�/o��c�t�%����*��������5��������T	<J'�E6��_o���RR�a����]U>�뒌Ҽ�D�í�K!�l��e��n��>�u��9��X�t�v���Py�Dq6R���s�in#�O�W�Y������*��%j?�id��<xL��^�M��T���]�PPKj����F�A���*d�1MQ�;�o`��mR�{��MlO+��V��R`o��%��`E��ߗfR�?2e�4=�+�e�Eo����ءaPR���Q�fv%�$HT��ru��gmÈ=�/C���>Ƃp�h��k��߰ޑq���Z����:e��`�ިb]���H��=q��f_�H��pS�%���J����b;'s�+"�Z>��PT�\����sy�V�����R�Ҕm�}Qs.���P�,���M��aّ�%+-��q6Iي�M
_c�aD������
ꐰ&�ꩽĐ,��B���K]��;4[��C5��z�&��JR�YL;�9D�I]o�T��0���5�K�ڭ�Y������Nσ����I�9:���ɢ/�S�xן��E�r��A�&�I���"3rPϣ配�Լ����������9_�荃�0Q��0p��=Ldmu�3���ǵ�i�Y�c�c��@Ӏ+5�U��%x��}s�Y�t�<0�N��֖5�dḅH�g��8K�g�Ec$�(wkzR��\w<f؜, ���m$W$~���(vȒɊf�ω���i=��1/6"��/�J��}����6��Xo"��y�)gD���H��)�:�C��4�()TKE�'>e���;x2�\W���L-pW��~%p�Č��p�Du�=����~n�QP
�Y�"�D��\���z����j]�T��2%���ĭ��C9"ߔW�vC����FӀ���Iz�@Y���J�=���!}I<��M�5�r�p��e��^\)r0~��4M���H�@h<Օ�����>�L���Lo��.yÆ��{� �:�e�'�m���>��õ�����]�a{5Ǝ��"��W(ܬ�e�NV0�1V��y���ϗ"��n���I�J�/Y���=�J��&B�YDgC�o�7���]�~�!~��QW�����A[Qdb�������밑�2 v��T�8&���q��r�U�'�!!&�V��c��n��dh�.J{�>���XMJʺ�jc"׾D�wU�҉%���a~b�6��Ѹ*����a`�v���٨�*�h��³�W��Ą�q��˕��@�z�3L4��Qm�q�z��v��>��=(p�$7����-�9,��C/�B�n?�D�un�6���!LL��C xa �(��C>T��w�M���i8�Pi1Wa��RGV�1ʸ�Kj�345M���3,>3��
���s}}�1��|W>��9vu��ߊP�Ҭ�^��z�P�7|&�)p��8�.!�5����������e�@&(���j3�+��wwt�ݜc�;k|��"����i_;:���M�?y���_��*��5�&����l��/FvP*ѿk�mdMdخ["]����n��-nS��y��XeS�%*ަ�N��,5�R�ƙ�(9\g[u��9%��s�W)��L��+����q�)-���s�6�a�p#�g��[�8��O>���K���S_&�A�Y� P�e�{��o[�^����&!Pz$���.���j�ho�}�X���ӜS5��W^��v����p���fV���wO��d6#n9Ųi:�?�� �����q9Bb:ኣ�μ����/���L)�Щ����m-�aV��&�ճ��4���X�sM`�fĬ�82���t~0�̇�b�B� z��j�K�\6|�0V5/'w!T�5j�<d(*mB�Hdaq������&�<)�UY���"��mV���#�&�����������~�uӿ�'�0���ߓ���~�ޝ�X��C.��Ȏ����՘P�i��w�9K�>�"� �9�sPu@<�5 ��ϲ4<�����P/�0t�*jc�ݻd��~_�p�MԓG�#���ա2�P/f����vjs��@Xs��1l��P�)����Y�����d����jVs�����(��w���M���+I���Rp���l�E|�%r�[�
�t%q��0��v���!�;����]$v�B��a���I�n���a��1�c��V@Cl:��d���8�������`�0)�YK����Ѳ�e�c?�HP�z���N�1�_\*,�ʄ�@�S�i)����rt
�k����S?p�o��Ɖ ����S#j�^e��AHE�Q�DX�J��b"!L���K�a���q�����i�O��ʐx`D�KabV��xH�d#Լ��B���GW������*x�)�w�