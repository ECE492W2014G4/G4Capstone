��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P��v�"<ߞ��&'��k%P碶�R�ӣ�sĞ������FY&S�b�Q�� R�H��)�*_�^~s��d�0�񿀊��EJ���T�m�П~�p
��I�yu�oY��[n��{�|	T_�3:�Q��I��l��7HG�F��O�.iP�Qdu�c���t��em�M(N��
�1�+h��w��m�q�&>�3�C�a?{j�AT�4��+�-`f�����n���s͢���G�Ôp��uw@�\���L�aSN�q�1m�iE�d��7��)&�^)�K�(c�kiE/F_S�D}q��.��}5k���+��pQ�3Y�����]�O4P~=8z�{��p�O�W��%(�`�Q��XʡX��ૈ�In�
7������1V��䜳��,���oɅ�����̙��KS���7��f('M����S�	���$�5�WjY��L/�O�b܍���hÇy�T�=ֆ���)λ�FZL%ٽ	;�Gb��0��$��d;8	�=����@P>ޭNυ�߿x��QOo�P Lq�꽌�[?8���y�ȈFr	���s��煌P�t���#��/E��&�Y1�E[�w���Mc�`[�?�
�p\�a����p]n�b�m!��wͫ�*��_^'��)��o�VW�ϿQ�5��>8�/��
�l�?wÁO��4�fE�#�V����¨H���e��W;w�`C� U�p�SO��e����'��J����)Q�#X�y\5�@219���>�7���ܩdz0+���Lm2�	��CgTջ���Y7��4N���@��zx��Jt+�fRP����5�����u�wd򜲏-4Q�ۢ4c!V��p^97�0��,R�T���k	�ĳ�4@�kCxҠ�f���n�7�Gkj3X�6�v����^�y�N������;N��p�pKl�-���x�7'�����?o|��*uE�)����;�LX좵x�����a����lOE2j/n>�X�>YX`.����'\.}�}���b������{���M���k�}����Վ�{��<	��x"��H��P%���;��))�AcK�kQuA�����r�[�o�H��[�vF��,��˟A���l��?�jV{��y�:ڣ���s$_@��ܸ
���g�����q���%/�F�Z����^OP-��WɄyjI�4����g�U�����'Z�s��P6���"��G�'o<�@������2,ӹΣ��tE�`�w�c9Η��7���jB��ﴝ����a�6�f������ j�V`H����"P�4���3���_�3�����p'��_,��ο4<�