��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>��`HX����5a8Sjf�&���>�m��`K���?�]^�6�,X�B� ��dt��\�<�bT�AT���*4�M�!�c@U�v��:B®�H����u����w&��*R��Q���\���h�NC[~��p��/���']ܑ��<u�˜�Hy�����#�������D��*K�x�����N���^d�Y�iZ�)7�a�k:���M�N��TƮc�i%;�ryp��C���-��Po`�M�w�6y�R��rDg���?�Q%���Nݣ�|l7�"��Mrb�0�9;�l($� ��7���
��>�9wo�Vx¦��G��hm2
������-�?�9(��lSf�6�l�;ϗ�Lr
�>���E.���?̴n��H�/�̣��h�S����/��!�����!���J,����I��e�z�Hsa.�O�{���p���p�*�\�P����h�ճ]���4���
�`.������4*Q�Vh����2?{Ԧs��g�k5����)@�x��u��m1C֬,s]�����x��%�b�.�@B�q�3k�q�zp�\(Ͳ��)'!�����;��o�sj7��q�s���yHG��D)s1T>�S�4!���:���X�.X��F���0_w%��ַ�{�[:�2��|ؑ��t[�tgw�x$�_6� t`��6C��9��}N#&��,��Hc�}.{����T/�^ۓf<�S&�R� ���E*��	;��*o��oQL�Y<��Rel�z��<��,��b0�y����)R��d/�m�֛��]�Z��Z�9�T��ޱg&��L�g,�`tb���)��`Sj;+��L@P�SH ?.����gz���w�%�,����V?�7�9��R6E�g+#\�����1ǘ�#��/��?���m}�+;T	(Q���q���K�b�4|n�? �]L癔S��.�P緥O����L���t��2ɐ�LQ�.�d���L����5��ǣe���%�	�e��rQ	vS��k�f�l�B-x:<��.2/cfA�QhV�T�5z���ɶ�RE�j�G�8�]xФ)�O�z��lє+��c.���8�*y0��iF|��[ %��]��a��1��ƴ	�W��U�f�iiא����C�"�4k���˹�BA��N?|���~i���������n����
 �ǳ�+�FJx���M{"�0?�Ј�.���>^M���Z4ֵ�xՕ�O'D`l��F�T|�]u�p�m��~MrK�?�e�O�}�1Z� ���P�;�D��VH]�U�P'U�t%6���!VY�I.Uz4J�e��2c�g��A���&c�v)/�}Kl#eb4��͇%�k=Y/�M�؃�C�	%B��A�&_�^j�����L�o���y�߹�Q�W���T4H�.��Ċ��8���C�Г��SB���1Ŕ�l^�Ѧ�Nw��L���)��WR���F�+1~h�r�at9(R�}����(�_˝�I�7�ɶd��v���bS�%�읙\�G� )���n�[	( ҈��JKE�4S�s#�c��sm�E��Կ��+y>u^x[u*�҉��qk	Ws:l-K"�!��������6@�V��x�y\s);{j�T�QA,�%	�kU@��5\��ˡ�{LV\�7�0�jS�>� [8/���s�<�G�����<g�j-���Ȫ:�C�*�����*t�q*������Ȇ
�\8�e�5� ��:O;5y����ݞn�8�q�l�|-��%�럟�;��55
��]��iH�,-�3r`����3�$�־R�̖�4Es�n��OjD}�s[����ͼ}Y<��*�9h�,uZ��DܝIkչ�9�J�=�|azC�����3�ǡ��K�Ι����K3�+;;��rq�4�<�R���ݣ���%�^pk������4qWZ҉�<�'����;��r�c��޺�`,Tf������֑q��/�#³g�J�׆��,ݴ��K=K�?Q���gE��y�8��GtYN+��	��4E�;�+�r�t:&/�ӭNm]�����Ų���v�1S��m�xKe���oI(�fC�MW�h�;��sI,��Z���%����*��g�:��o#�h�J�͗-J��|����L��Ń�b�J��b����B���2I����6av؈_/�F�@�0��x��Z�Ï��d�J>�h�H�y�7<Y��N[�׊bw	��
�����J,9�bVVo#	�E{%�� �U����U���Hv����	� ��JR�G�ǩ��������+q�y�פh]���~�D���͒ʽ�+��� � ���z�S(�C�S'�9�.���Hp�1�����b:Px�Q�Զk�b��1�@J v��]��!�>���b���|��쓩��')GZE&3Q���LrѴ��*o/�O`O���B;�`&�?}���(����*-,������C�e�Vc���W��[?�!�Qn� ]����{����%79淏OԖ�ɍ�j!by�'����M�o0=|�S���54��[�F��j��\0�����'�J��?��fӸ�,���1Y/��O-:��V�9���	V��̳F�9ٛ�U��ǖ
�^���M�6r�&��C�����������:�����6��k�ռw�WK�"^bJ Ɨ�S��Ȝ���%�9s+��Oέ��߈(wV�ȁ�*"�����Y�0��R�C����Q��NR���@8�n{2��8��ޚ��֋&���i�<J�=}��
�G)�.�.l>��C�'��bd��Y���~�졳��T�.6�y�Hį܏���_9�T�v]��Fv�� ���/�w��1���Ԥ�U�C���Y�a�/!Y �O�3f�]_k�����1�I�[���g�����ݦ�o�]yV$�*k�����I[����Is ��;42�F�8=�9���]�z���\�����,����(L}8��y��21����78�fq[�G��@�z��a{�Eq���8����T��+�����\)iƂ��^>�gz�DOd�����wuX�����̑#�ӊ����RT1w�)�NԴ��m'���8������T��L�F��}�c����5�,���4�}�yb��a� ����iQ���ҏU�A<�-��'z�:�>�"�DSo�ٙ�$� Ɉ,��Y�)�Bo�h��ޭR4��HhK��46��q伂gO<�Rp�+^�|54�{�O�a,R`A�`�����c���UZ�-�~\���!MKx7�2m���֚u�0|�����(K_�N����Y���I��p��b��8�2����B��iu-'1I�E˙w9`��-E��bwc�^-��H�v���[T�rQ�ט���:�z��7Ώ�&�~c�@GB�*�ׅ��V�