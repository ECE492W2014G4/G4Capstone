��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P��v�"<ߞ��&'��k%P碶�R�ӣ�sĞ������FY&)XH�g�'���v�D�����ש�����Q�g��-AN $m-�޿� �Eĩ��",۶#�=�ЭS}����x �!�����#����J��7�0!>۴,D�����șصjV7��6�nq��~}4p$�9���ß��p8�Qm��{|\=v��ם�i���JlQ՟t�a\�5d�r�oz��dh��0R�a�����i7{�	���a{�S������"Ӹ�\�"0��s�J��m�O(�����p]��Ǘ~̤��8�5hY� �ڴ2X@B�q+�8�����������H�I�f���撓���Z��"̃�x+��t��h2^Zp�U�D?$�^	�q�u�Œ�L��+ļ.Jݚ�ۼ�yņ��Z���8��Y6]�	��}���%Pz&�������C��vزQ��F7�s����W��T*�|
��^b���\٤%Ͻ�j�����<����Q�s9���c�5�"�����o۽�M>�X��D�V=L��+�1<5Me7������x�d��vǽ)c�g\���yzF��t��Fl�W?��R�g�T�*j�仌q5Ib�Pӂ��򕺿�῰�6�-��Q��k3��4"����?���!�����i��]�� �a��-���#��At ����B#R��s9ݢ�_��Oe_���8j%�;K\)j�ߊ	�A݀��,ȍ|�8D����N`��˲�f���5@5!�D�l1�Oi�#����Xg�ڸ<���
л���x��[B#ם}�r�����M��������z��E�-H��9�� ci��1n;gJ���@�+�q������-Ɏr�?��-V�b�A�-�e�0$G3��-�dG�����l@;���c���7�65���}��f�V_FLs�ZB>�w��������^�%�ޮ����ԥL����pSz{u4�v�����?$�x|�����pqn�m)R�%b$٩�5��@�A��F�fK���_�y0ȋ��3�f���|Q��Pqv��3p�y��)�7�3����mm^��Fߙ~�Zs�G��+q��B=�6�q��B�`��:]	ӏpd*�����Qx�$����W���Nz/5mO�� ��"��=�9�+Էd���O=H��-:px�::-�
�U��b��I[�	>��P2/��	�Fk<0���{�Lh<ḓq!�ۡ�4!xPU]�f���QU�V.�S �v��:��e��E�P�����x��8�K�tA>����I��wV�� %f��	C����e/<�����1��0@@G`�����Φ��#qgs�>��BJ�,���|<��|:��f�π�B+9��'�U��R��@�ݿ��A�qR����bT�pw�B��1�>@��D�3��/ ��5ڮW�H���o>7�[��JԎ�7��1��Ծ_�ǣ@B�ׄ-8q�]v�Z�Z�$����=+��`��LWG���:@86X���bS�LP��Ch��l�f�P���� 	WR�||��l��"g^1~�'C��s/�@��F ��Ģ��0�hsf-b��Ϲb�Uk���"/�*�5q�F%K	���KU��RߘǋgxB,�6�J�gJN��#o�GR��Q �E$��ZI"9����rU�f?Ь�|�Q�g�H.s����_� ���y�:)����:i�j�ԃ��s�ǳ��3�G��Q�(����2p�J$Át��f2�Ԕ7�����	c��ѫ�)����Z�~&P���dDA{7������v�zZ� ��u�nz'�hx\��d�`���]w��'��8W�� ͮg��̳2�#3Av«�E�v"�	��]Z�p6��t�#6��U�$b!�$I9��4	 �ht�,��?��;#��6Gʿ�E\93"%��]�w�������$̨S�)BA{e��.��߇���9��P��/��<�f��f�pG)w�*����+�rM����i�6�0��{~WA
��w{����OeE�&�Xk��� O�S8 	T� [^ǜ�ߏ����������2� g�Ic�m�k��8K�43���'���H��&Ħ&A�Cܭc�)��)��s�Y׃&% N`�
�v]�}��q;y(It
݃t�� ڭ�>�D��fwpo/��r�_Xݧ�t�%�R�����2���HA��	����C�TH�KP�l!f#�]��|�?��7 z����4��u=��rQ���&��Ʒn_	�:����d:ɯ���2]��3Z�t]@>�O\7yA%i�i��8s��u�r������I���+<K:U"�/9���(��!�� ��m��r~Yk��g�2;��)�)������vC�8�A�jS����7K��}_�ۈ��!�_�Z���j =�$���p�������`�+}���W� w�w//�����K�&_�*]�pȤ��j,�'avuDC��n'�,���؂ q�;�T-��r��|�<�3������1M�o�|?�8���Ӌk��A7[��<�����CQTl�}^N�f�z�r��{����eW�h9ij�]nl8�wF��;=�P�kf��)�T.����,�Mݨ�ƌ���ׯ*����c���u7�kX��/	�}G��,���,��y=	�^=���b���8��$s�@ǹ�$yU�g^-bs���e�k+n�������_�5��h��\^��y��ݪ 9V׃�8���a�G�+���8�BZp��V��=�t�8g����<O��ﻸ�f��_��~r�I:/*.ɣ��'�x�U{^;,pުܹ���͐tM��4ʉ�Zg
���Ɨ�
a��$���c��ľ��QMZ����N%�"x�K���{Z�\�ү'�{P��̫s�E��Ł���I�eW��ߣ�4f��v���nd��&��!z�cM ���%���~q�U|A�X%�L�vF�(z\S3�)9�g�F.��_i&dY7q�H���ہ����2�����L�4�}ZN-�[��~U ������ܸ��4`�ū���&)' o'����/2U;�nH3���n���9�4��)�ă�`�S�����_���a=����1��9����0-������]�|���t�mq}�� '���E��tȅ����ɼ�1����^�9��r���Ǖ����{�sS�'{���Z0���h~[4��Ɂ0���
~ijB�\���_V9e]I��W
�`��Z[䜜�����#2ȼ�O�����Su&elNʨ�B��Sm���qi�mc�#��.3�A4���� ��ixU��!�~~^s�Kt��1�Ur�bh�ԇ奎�Tt��%����k+i��BN�t 	�0��$��n�v�Da����7�]ƃPyu� ���B>l�ǥ\���O�ȱ�ͱ$.a��W)���p����O,�Ymio��l��?�;�9�z��}�HQШU�e���LG0��5݈�JSK�o�-K���xA/⧘I�XL�i&7E��B��������T� 2�A)�OCn��gaT��`��L�D�ޝzy)�lw9����\ݳʣ������4��7|?���0uCN��gnPpE���i�{b-o�[������E`���n����b� ,��*P6���T��6�$���W�t˜y�5s���c{�/M*}�FԩP�	��k�k���3�@��v��\�-؃p��H��I��n<2��[n����L8A�z�1슳�t�7q�ODK��?B^X��u�q��ת�sj^�f-������� ��I�1�_~.>i�H��qyp��(@�r�i���ڟ��{�������� q|M�=|$ ��aa�+]�������7A^< �_�p(%6	�PG��Kv��LGTv�N�S�,Ĺ��Msp鰎$�C�Ӏ�+ez�YW@�M:���{3�3�I�JA����M�C�%Hs�۞��J7׬�=
i�q>�jj��jU��"`j>�N)�0�i��0P�]?�.Iv}�x
��*.�W��HO�L�yN�����B����Le���$��J�J��������̅��TD��Ω����)��lh��)ӹ�f�K]�k$�%J���9�0O������}�� >hW�}=,~���Pm�H��9'��Q�h���o���4��B��t8h�̈́����|��1f���Ե#�@=v�Q3A��[�M�s�����fJ�Q�iǌ_~�_��������S��y���c����Ї�D�y]@�yuR��2t��y�F��a��{�h?b�Z�f7}ﾘ��G+�@~-Dş�}6�c�\ÀT��9iݪ�0��o×�m���2�ʤE�>��i�'��j�̞M[�(��qֲ�R��~�T8���9@�nZ&D	8y,A�v�O��	�n�C�\U�̳˳���4{E4NG9<:��� �d�`�3�TYu?ޭ@��]>|�P$����"M_�!u�'3�q��a��>����o{3W-�<H�����i�@^�lA]��[`� Њ���s�v�����=9����'=��0��Y���b�;3''��$��t(���ݾR��D�׊]OD-O���Y4�����Wr�0��U�Z�����n"B��W�̇<@
�s�U��_��p�K9>�]���n'G4���~�߰2�vnAy\o��KY�5�!v�FS�Z����4\�|�n�2��v1 "F��c��5��Đ�or�����י��`NDq���y5j.��������3�Ɏn`"��
c���gu�>.��M�i�
���`},��e�0H%��r�N���������顭r�W�O����b�W|�E}C'�od��=�����?��O~q�o-F ����u#�`n� y*+�?�;%�V��i�ph``���"*ֵ%��	�;j��	4�_����y
��l�j�x��k�|�pP}�	c�v٣��|5wnY=D���{�-jf1iLcK�u��H�%sɑzL!���O��e��#R5m��MMyn|>~(��f	!�9'l�����wY@T{���-����t4��s�)}�-V}�#EՋ���x��Z�q[s��9)���C)���唋+[���nU�\ALLL�F+��:�T�o� �&o��jRm�8-�t� uI<&^-�\��Ԃ0&{O��������CXP~��	�av�p��So��a|�h&�T�&8�xa�iB�����y��