��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|۶��-�Eݒ�s.P���ޢ';���SS@;t@��֗��Fp>��6�{������(|�#�����jҜ.W�DA���><ugLb:�	�bG��7���S|GA��]` ^�G'$ƪ}?KT�.�<�<)�rX��}�]X�a��dp��	jN嬓i��E�~Ū�n���4j�G�c��t���x38��A���g>awFP�ZSYxho�� Q�b��k�1FY~��u�;8s�O�,
N��z�m��Q�ҝ�d9�0T�-�z+��_~��_��`�����n�坆�꧸Jɾ��A�=/��b�X�g���4w����@A��ח�˘��qt&2�k��u�.�������R\@����WA������/���$vq^*�)L����`=u�oDQ��{��/i�����������s�����@-s'_lZSrD,�Y�"�){�� ��+�x��E􁷽������t��mX�z{;��C�s��ʀ_)ب�n���U�k������ؔQ3�wVBi(���	'�s�n?{��Qo
� vz�/xk�m!�L[���ɲ�F�;/K_�;P'�qB�o�� ��r�w���5��r�����TL��kI$h��0d�j��hڨU9�t�dr�F�)ѓ�w�0U�3+ˇ��j�Ȳ����q���mo�|��ő��9ļ��e�E�}���X��hQ�jEȃ�|�|H��1U�D��#zM��	m<�vܭ����&��eOnv��/��s�d�%<r�%��z=�䯁n���fզi�V�Lbs�+�"����~��Wp�vx��P+����(�T�y��#� �Ǻ(X�+��k�|{����Hֳ#���L��u4�@�t'��{��YaI<!����p�"Ĥ�N��R��_���h��g�G`�Bp�T��a�K'7��c�Y�!.�F9�\�F9��x@�.��\Nˀ�3��i3o��y��8��yTE��<�`R���IӼ�$�����f�o��ϯ9uG�oO��@���⏇�ٰ��]�~�A�0i��ӭ�\G�y�4��������Q�G;���G�ɑDx�NULQ�%�d���� ��R��9��b�-X�A�9@�fEZ��7_���9�. S'v2x���Td�I,3F�4'0�C�l�ʹt-KC$0rR�y�1��Z��(�@)��@p$6 y�mRXo������\}ӯ}�*�Ҏ���\*�=$�r ��vT� >���`��;�����=j�
�Y(gM����9:\褶Y�r*b�YA�y4�Gx@&���\�F5��h�(zd�-��Ԁ��}퐌��QV��d� �1(l�7�48�F@p��T���q���^�9m�����H�:{Ė�@�x���Ƽ��bs,2��Ψ�h<r}�;�l��@y@�|r�����Tw[A0Ͼ� ��C5��p�G�L�p۟�{	!�֜Pu��aG6H��3ut�K�lS!��N�d,��M������s�i?İ�d�HM�d���ˁU\�Wq�޼]S�E�0�9�5.T��[�/��0��MFb�)e���(B��3���Ax�L A��t��>�D�V�;X�غ�<��k��oO�Ĕ�����:�xr�^2]R=��[�y��2#��M|e�~Ts��4&�(�ć�%�h���![W`�#5��
T��	���1{�z�̩�;�m1�e���+7b&Ⱦ���Y���:Ћ����.a�/��7d����@����9��u�� �4���.�\O���A4�u��7�K��ur����-��J�Ve���J��1J�7�Dǫ^�hs!?.���C�]�?9h�'wdXpP�it@JC��-%w��Hl�;]1�&�7}�Sn帬�:|�0�a���ښkJ�U�i����ڷFY��ܰ[T��� n�r�V"O��+Q5河9��x�J\��G�Z���xS�ڂ���q�m���1Yw�:Op��"t[�]y��jQ\J�ס����MD�̴�[�$,n�]�����<;'��vv4~��-�):tM ��K���O�z�}q�d��\37 �?'Vz/�����A�z.�]��(/&���Dxcl݊X�i���K��Z�(@��?nD�s�y��d��sf������=�9v[8�1yBL��Q+ \O+dD�7�z��v�w��\g���K*�'gj2��;�$C1"Jl�
�ll�MXl_��� ��4Í������,�C�'lj����פq�lT�GrnͻųWhO��}���߹��q�fVs��*�IA�K�p��71YJ��!�ق�r$E{f�Aݽ��M��4n'��fg��mL �b�~┎ou��Al"����#҅NY���(ǻ��2�-Z�6*�s�� ��=�ls�--��dC�믃W�ټ>��I��
Uč�s�]�jʥ�}���3���<ו�>���\�5�3�L/�c"����{�A�3�6�[� �%�ofSh�>��h5߬|̶W�(�;�����*(��LW(�n^��]6�S���PX��)c��g�	�u��Lۿ��zi�D���~\E�zS$o5�<2�r���fm��#�@�4�(0\�T��o�O����Ѩ��ʽ���^�ǣ�_Λ��L|�;I��jr�Y�}6!� 
H��%�{²e1�łzӠ�Xi*{���u�����/�	�����P�s�-��kV�I�1�[�bSeӊ���NScm�vYk9�! yI�SD��W(�WJh��4���u�̇#�q$�A�`o��U82�8�=�/������X���6:q�̳��>!oH�sX�=�I~	��)�w��Zu�صkN%�f�_�$��IT��Gp�Ly�U��������e��{�4"}��̠���\�-�[���H� ��f���l4�@yjj#'��״��(��v�hZ���5�z�l�E���W���z|�hx���5H$�=E����Q�W�%;����Ü}g�S���ؐ���p�2���[ø���]N��,zŇ��9��Q�
O �D��r=����7�B?lxk4�l$E��i�&mEESV�q�c��{ťQ�'�Ǿ�Ol6��7�2h~��QR`���mi=�^Y}Y�O!�5Z��mWL]�1��ˈ��1�"s׮�D��de������e�"�f~�T��6}���e����`�փֱ�n�j�7k��x�G]i�C4`�6	�"Y�n��sm��s�JSf�!�����ز�t�T�&X����\�
���!OI���0;h��;݋xDY�'�gXhu�9y�H�}�4Q��RUF�kOQ� ��)��4 =*L��m)'}����T�T�����������
C̏\a|7*%�F�Sp�s�Εpb;�"����%�uP�-	�I���Y��C�Ͳ��b�{Z�w魤Wծ��ܔw��โ�6�������yCD�O䀲����VZ-�<��/�&�����R���i��4؊�nؑ�f�-�BLl�]y`
@Ty9��J�����<�,I:�ӹ�$@���&US��F>]��\��I<4�.���9�pۼ�D�f�%kq���h����o��P����:r����w�iaZ3N�������E��ƍH�Է��A)�ܑ�>�43�mf���Ĉ�;�����UCV.�j��������8��Tԃ�t��	!�U�D�:��tؗ���T�.�/���d���$7������%k��	����4�8 g����'�V5� K=�p/R��[Nʿ�J�U$J!���Sp;��,��>��v[��QT�hP�F�jw[�fg����bȇʇ�I�:��4J��4cQec�y �D��0� �W�8Q�\�Y�K3�S�F!�ᐐ-xc6�D��h닳��v��$�/��d�Dۊe��(��ܧ!�|8�D�ͩ���BC��8<Ԟ�o񣖕#�M��<�x	�il&cex�6�۫i(��<{h����"ղ8�o����d7,��_�I�7�F]BOb}-�\�~��ʵ�]ڤ��D?r/Ş�!��=���-[��Bu�S Ã������-���1|� �g�q׼�&��Z����ʍƗ��)��"JW~����,�R���	�ZH���i���X�� _n��7����_"3S�F}�=�t���J �jAY�'�^@���wM�"��^��+C�`���;|7zھ�e�#�/��v\���di3"Dj�UF�njchEC"^�'#G �D�5TSV_59p���n�v�D��Օ?䥎��;��	/��4r��c�L���u����y�y��[����= �ģ�d)��?���;/22����l�XO�=h��쫌u�o�?fW��aE~�ACՇzȊEºI�$'���P�׾
��{���(�v9��\L�2����W�u�I��)'�J*h�u��e[^b��)�c�ʄq�%�����E=|��Pak=�=�����/�BY�ܘH�U5����[h [���k�ö�^���?Ϸ�)N�Rݛ��,V�5AٞK4Y�L���uΤKV%`.W�q*�C8�D�s�1!�)�y=��Z��Iw4x�u�P�1��� �Q�o^��,�p�8E���3�$���v[� ��MD �X�:�+��_�Z��}�.]�|�o.Hkx��J���|������֧�VR��ۛ�$U_����v��1�q����*��녡�"�Zq�/�b�0)���W
���ҝ��[�m�.���W�B)��6��]�J�kj�ҟYf݇���1!�}O�e�-�Ly��O�rK�wfl�NW�vQ�z��]���>L��:[����Ѡ6�~ds>��o�RI��.�һxQ���w��c����m����oz�K�f���^M��d[�8�x3�9���������� �����h[� QF�N �C��ώ�ǟ=���g=���S�B�,§Bͽӎ��x� b2��\V�V��(�Y�W�������O�
��Č5�0��7�o�7���
M�%R(^cyy�UD$4d�yb\9k�%�x ����E�;�+�")�(���/�����?���l[�t��GM"�.-٧��0IK��V���0�A�r����J��C�hp>�w�Bi���uLd)�z1��9m�_���vmF�r�����@w�!��0F�Ɉ�r��i�1�n�ԛ�"����'3v���Eh('Pb����+�Z57���>o�pO��b�}�Y��,�~�f7����3H�4��"w�
��7{�������6�!r	��܀�-�ǒ���r$�k�a6?�¶.����ZDe��^�~\e:���������ЎK��5MRz-���Wص��C��r��o��g Q���n��)&��(x\f�\�:�Ю��sg� �B�h?t��&�_����;�㒺й�[?�iU	�
���'�ueA�ȍ��x���T���k�� s���ӌ4K�k�.����U��\֓�� ��g�ff|����	�pb�	#rR���E�Xv��UPH)�m��3{�t��T��6B���L�(M���ve����U�L��8J������ǡS]����s:&�"��; *jU���� #q0����qh5-�rL��S��>�%Kd/�q��
��᥾�m����b�ݕ��\7�r�N]�IG�kC�*YBi�<�ve3`��{���C�[KJ���{%��ѣ��yc����sy����&2d�(���*�.2�Z���@]� �l�^�!�7�@�F�.[o�AY��2�m�0�H�:ە�w�vc���֊_���#�}(�-�"��ОUf'>�,���VT��.�*G�����i��d"�KĦ;/dp}�[���6� �?X�%ȅ5�6��i/����V� �Q��k���NH(��퉧���v篑���
��f=;�p�	+��DƽK�X��[��QAp�a�1TOp��&�^8�6���S�	wW��Y*��M��� ?����!��Uv�������I���/����3u=��vz�0��A]1�I�f�wqy K��s�F=C��3ҝ���v
(����! �M:ɜB�KN�}��ƾ��{^�xM�{I��k
o'g�>�����o�i[ �?t��U���j�B�������V�6HN�%��\H��uU8/�FI�v��!��`휭;P��WE=P�����(���vA�	��>S�6l�#�H�8k�	����UZ#�q	������d�%��OG�}1F�
��
�[ώ���$�Cp�������,Q Z
 �����fΧzˮ��g�e�/}�q�B��`j��-L��`.��D�w�7˱�\L�4'�߭�و�[Y��_��9:��~�4M+Q�\����i���DV�c<b(���b��\f""5XO���8Hd��{��;
�Ҋ��G�2�\h�|�%o����9�����1�1 �C�m����?�n�͐{�0 Os.�u�@�n���@��"�����������hbE���sB�@>s͖r�o���h��.�NUr"�Sܶw��=<:	��3�l?خ���,;d��7��nce�
R݁bVSI�A��`!Χ�`tTH��%0�����o٣k$�$W����0���&zWZZC�}yO|C�S<<�k�)|ǧ�2��k��'�G%����H��&.U(H�?�Cҟ�Ku�&���Ű.��R�A4S�؟1���yt�}W�؞���&gx&�����[�IF1�l�󯠊�^Y9�v�N��� ����W��
��"�@��J�X7�
z0#h�L�t=�3#����C138�A��n7����|ΨH6��O���v@�f1V<�-k{'1�Gd :��,_�u�ݭ2W�uB�:��"�M�{+[��.֌��%�S&ޚש����t�f�VM��A5fjhAc�׏1"��y�}��N��a_|�x+���[���w��ύI�= ;��X�d�Y�W,��4ҙ�)iH��q3��Kx\�7|%�ebWm�KFE�i�(��YCϷƈ��Uğ�v� t��a��1�������fP��q'�Z��a�#��f�~�%֘������C	7�خ��9/����/0轛p���8��o��2�e��	Ȝ�����u.�����R0P��uhdI j�7��yh�D���\���=MZ]8~+c�H{�J&z e�W��>=>�����ϴ�j0��.P,�.��_�y���e�H�?�:�I����b��F�k#�'G�H#�ժh�JܘVL~=F_�YS���h�
ҳ^	sh� f�"�mw|I0��l�{5�[S���7���q���[�7ٚd��|JA@�9�+<$tu�w��q��T�̞Ӥ�
E����!���"���WRU�M��瘫Q8��>`>��mz��"��qƖ����P��]ĻUIOR$��A�<���H���w��G�y���"1W�[������:�q�;�b�i����N	+�mdfYSA�m�Ӹ_�-
=��8����3K�T�'����=�^��qk������hmO����.{�����v*�n�00�@�*p�@��-�a�	=�d6iKW�2i��q`͞ch4ޥ&��'N�=�ЕQ0ӯd>9�� !�3��Sk�-�I�'NF<x|8Գ��P��v�o:��T�,u��o�?�H�tՊ��ZdAb��_�L�"Av5 I�j�OŜ���-G�ɪ�q����:��0���;7`O.�_9R�'���L��@��������- .�w��X���`��_ �՗�(
��?c W%d��~]���)>r��Gt<xZ7}���,�.�a�9aJ��l�e*�+=�}�ӹ�3����K�H�Ȧ�c�R�XC���:�!�?"��k�^��ָK˹�	$<��Rrl��=�~e�H�xU�8�#��!s�N�{����C�����9���2�	z�!�&�|\Q����w]�~8�'�G��b���ƽ�rk����ML7��u����?P�����iGNG�bu�8I�m,a�k]���2�"�؈G��#}�}O���C�l�#[��ȵ��K*��8yvbCS/�����]hOo7�9�UH�{{��ՅC��K�bRW3*�Bt�o͟���XC��ɝ�+����[�ѫ���j�y�$!ҪA.�7���A�.�#�<�,���y�ã��rG����ao1�\���� Q��Tj9)�5��Qͭ���1�K�@%��q�(���>�'V=G.PP��������CK�[s�1p�CV�Q��4;��:��6�^	er��>�v�f<z�x����B� ��$$X{v����l!�Ts���Yм�ya
ߛe�L�).[��������Z2 z��n^yd�t>HC�N�(W-6N�xʶI+��3������묡�v�ܙhy����g���Q�<T�l�E (�%Oh�k��1���C�s7 9��Kwv��@+�E�a����}�7�=zR����G�V��Z��ٿ��woj��zo�%@�,Q�ok��(�%y�˦������Ἁ���d�G����n�γjB�%�{�%
��aӋq���E�4����8�uc]���;�N�Q�҅�0�o��u3*�g;����9�����~>��������ᙣ�է���$A:^���'(��^��Lf����O;+�Ľ�+��PNs=uw�F}��ՁH�L�4z26�2�x�w�p!$��ƣ7��ͼ`��<L��l����.�?��߮�T�]jV�~�q������u�J��8�ib��N�{�u�o�£{ϖ]}�^4�7T������{X����p���Y
�c�S���:*���c�͎#�pĉ��i(t���PN�1ᑞ�ӢR���/�N��#�{3�7g�sOu�d�YL\��4�>���n��v�R�WNYO����҅����8�)��)�u�M*�M�w�/���*���'��2/�ʉ�{h.L�-���;>a����v���	��ծ��Js��8`�S)�Ak���^k�'O$$wT	��2�U;�35�A�R����g'af�v4�S4_�튫;y1��.�Z�wY��Y��ҩ5�c�k��	s���l��)9�������e@0���?SO��{H�kG|$7B��Q2���A��};���n��l[OR�Z��wV���h�&H�ȵ
�_�T�bV{�U�`s�\ꅡ����I���]������'1bT)�Y�9�Mi-�M�����V:���0 ��*��' �U;}"��_mD�<�D��_���_�'E)bz�<��D?�H��4��g�x�h��Z�y��!��#wmQtm�,ڣ��B4���O��]=l+T�c�Q� AԱ��1-�@�6����W�c�3S�U��/�Q*
hp���nV��F����k�x�g/{`���<��.�ٺ"m?EU��u��)���ʊ��`'-�b6�{E��<1��OL�Eh��%{�o�4�A��fk?(I��)ꂖz\�d�]��9c&�B�y�,�p��?�,�Y�m��I=E!g!�����7y>D�*|m�*�"��I,m���^�M��$��ȘXq.Xd��Ӂ�W�4��aiT�Y���-�3���>�d*���ߘ��§�N�����3����:0 �/��hE\�
�~�K��#��ݬ�C����ˊn��
��L@�4����i�Sm��T�9ѕ���)���p�oӟĞ`�F� �v�f��<�_�Y��g'*u��x��yYE�������Y�b�����m �.�m����")r,���Z�a�@���HL�;�n�5��~�����z*�VOh���p�H�K���]ur�v_}�=����oǴzC8i���9%�l�]+�XI�l��2�N�e��C��89�0ߛ��-k��Pt������� �0~m}W�쏁w�������\�E�p��v(�E'��E�,��ɈvY19�$�H}�0p��a�ju.ͺ��t6z�\�����vDߘ��T2�t�u�,���y1o����s������}&�JsmZg����v0�<��9�}W<��&dp���X*-u0���A߹j�ɹȳ���w��R�d$	�\B�}2�٪�xB�V�Gm��K�8gߠ���[���Z���~]�q��҉¢���u|i�-�{�`1���~&�0��cs�V7G+Yxu%�QE�j1�����������n(Ն��^?>��3����� )%���uGK�]"y��k��Gn��P��c���������4e䂔�ǌ�����iE�)��M�]�0dė���4#�j��.������$5_ڵ@� ����E��(�,���u��d�KO���-n����J(e�df��f2$?�Yj��B,���B���64a������h�8w�鳖��m�"ހ-��ŷ�A��dS��3m0�qZ�"���s��
>Z��+��[P{0I��T�7����.���a�j.�'��J���l�U[煦'~�C��rU���Pa�����&��+1��Z S#�0�m��]�=�Gu0[���͊v~��P���|��x���B�~��i�,�	(X[����JK�4���g}M�2�6��6�yE@����|�/�+ae+)��Ҷޠ�9�nI��*�_`�?o��X�5Mz���?_�Y���Y�.��x�3{c�Y����	�G�\�ׅ��$:.,� ~fG��bn���W�E��Ѝ%x�H�U�Bo>6��h��>��C/�+<T��u?���_!e��埼�\H�ظ��9�	���/,�p���E�jv)o��ĝ�����b�^VLp�fB�9)�I��/�R/>L-���;E�J�����Y/���0����_}�zԳ �en��9`U�^��O��}�.H"H�,�|����}d�V��Kg���u��"}nH�U��hଈ|��nU
T'�����Y��/Qnᐅ��ݗ�!"]TQ��5���RW��� do1��(���9Y�<�����l?�=��~?t�탙m�7.C����f�����z"Mb�W'@�:�yQ���2\����ik4�(��DVgN����.�C:��� �tn�F�-~i��;1���!�T��R�֞$?�2{:���eF���eA'���(^�˿S�V��P���JԚd�������Pl������epu��oM��'���rkx�3x�;Pz~��0_Q_�)��P_LRd;��1x�'W�v_ 6�y�[�#�)�	��t�E�a��7���l�<��"�&^��#�	@��S�+ ,�<��}����/;��}5o:�T��Ƒ�y+��<S��_x�5	ۙ�#.8�P[���C%�ߘ��_I����Bh�7�ADhc�< ^�neVg=��.CD�O��[ ���b��'�M{A���d-v)PIZM�#�+�q���[y��aϗ�p�����@ӫ����p�S�T$�(7�R�d��C�º��i�ci�@.^Y�����8�w��K��\>t�;%D��!Sc.CS�(�?P|I�^ų��b�zt�Mx����m����}��C��f���Ho3�������$�3Ļ��|X�>!�_1��k]p�ޫ������������5�#hBŰ�(���+�k�3�S��S��YW��{��ly��~d��/�!��g��!gަ��C�T���Y��էn�Ґ�h� ��6��$`��y`�S�?B��5��+�P��\$��[9��H¥	�e�.(0	�5�ց��٭�Fc��ח�3
o=��7},�n>u�C�2�f�nTQ$?���:Ro+���f�	��m�H\[$N*#o52ೈ�I����j�t�"�����]� \�֝	j ����&�<�� Ӛ߃�\���LH"�r8�S^~-��՜
��!NY�	@-���"S��|�K=���h�J�R�A�5UB^� �Mxzk^�\�j/�Q�׻v߾^S<߆� �K Ȗ�N5I�X�6��!}Z�NTgMئ��I�B�eH�
�-�������,L���^k�E=V�n��OZ&�zF�n�3��N���#`J5��@d�e]��H�_���8U�,��.����Ж8r�e�k�8��9��|Ph9���I��A�F��Q^ ���L��ш�a��Z�
d$��BR��\n�vA���jR	�Ck�< �_��T'�Q`�wY���RhES�^~��^Xgo�f�؉+m�� sh�xڶ��gC=C�]S����j�/�/��cد17�T�LU���0T�)����'�H�S�ُ� ixb%E�����.`�W�{�D]� F�-�v3�|q|6V;�%6|��'�Ŧ�I��,"#�����I�o)Tc�2��Ϝ�53�ŭӔ�	�/�Tl�Ea]�����e�CH�.�U����ۄxp�z#��� ���pPPjW;�� ǩ���pEU�4hj��>�O�ב�0��F���z�jtg0���V���>��3&S'������'�\�'���mr 03C�Ћ��o���-��Ŀz,����ډ�Un�g�����sO� �6����`}"��U=�!�/q;�ak��?r
�/O����n�qN�OY���IMQ��N@Il�;�|N�k �Z��@>[�Ei����!�'`�'��s�\�x%�g�xL
\���B��5�T�[VrWh�r�o������KĞ�{K��ڀ���< 5B�"Yw[7�i�_	��Xٗ��5�1�L�����gj����������Ʈ�B ����=[��>�jH6��h>��ߖ���b�R)��y�9R�8n?*����S��&�l����p����-=[�r��w@T�wP�z*Oͭ����6�h�;)��pT���Q:�~�T��W��<������6˼�rh|5�Y�D�YA�ԒQ����UJ6!0�k[���Qz����W9$w�v�;U
���	QI�û�M�G���)䳡�4X����4<��B��L�JP۬�>)�.ou��q�v�M��ds�D��E�9�Z!�JHp��\}{�I^���h� �{�u�,���i�V�#�|B�<_AB� ��JC��[��?7�4t�N�J�T9oo<��W�h(�4���j S8ē�S_r�WDc�q�jaH ��uM{���i���T5w2s$�f>�[0j�c�jP�?��'��g�G�ذ��||��s�8X�4���u@��c���@�VUo:��6�@��l6��}���H��B�fV��A.���S���7;iOf.e�y����Y�:ꅘM~��F��3-BS�5�<{�7�42��we�2�m[e�Ң���E4!R�M��w+�'�^V��şW�Kn�+�_٫�>8�%_�_�g�
Q���7I'w΁��*Y(D���2�2�=���(�T|�x��� �t5>�3%��!�E�2T����"�������,�n�==�6��C��a"��7�45d�[0i�y�ڇ����>6#Cؿ�x�b6��;|�e��%�����X�ث|  }-��&����jJ�`ȄJ?��֑^���������p�9&�>t�@���tu�Ih
�Wp��ō{׵�u�܎Q_<'c�V^���WpQ�c�q\�o��5��i��S����LB�g�.y�ws_ԯ� �"D���bu�M��a8�:�V):	9CT���@� F�V��pޗ�����a��bx�p�+E>��	^�ˊ��JIX0�K�BV�Rx������T<�4_�c�fƮe��P����)��Ih�{˥?Bﴟ=Dʗ6�A����h�2��+����6c�Sc)��!�����,肵�[^����� g�]%�G�!2bk\���m�ؖW�9���Y�1¿�e'tAd�Zfm�	��׹�-�黗)�ͪ�VÄ�a\�2ÿ�:���2e�&qe8g���>��:\�����l�GIn$r�Dv-K�&K�a^���G9���_�Gh���Y�M3�&(�[� �w���������S>���3/�� �쎈��.�V��괲9X���Wt:��)���V�g	k������u�`�t����-���?n)��o���,?���w��g�7���bZģ�J�b�?����:߂/�R�����H���T9�����5���ޭs1�q�[?�a~K�B����R	��e�v����̚�R�[��ଙ -�#��n%�?#|������:x1;�}�����F2N��K�Ͼ�Y��1��K�Z����.8((��*��uS�˸���5���� ��c��?q��TO۠8��T�ҾY-���=�q ;ಘܘ�μ,���.��н�j�1?v��2!W�ىk�^�K�>EC���խ+D@Q�&=����D�e�����!���͡þ���U�z�OTC�&"���P
i����9�}��]���,QB���?Cb��9�5~���6ǩ)�������0�
�a��3#fq�]�*eB��0u��3W'O�iā�:P��7_%�&���@�$]���V�l5ArZp��d+����6�=�Jl�n���*���K+wް ������JM�a�����t���a-�n��Ɉ׎��Th-��J�
��9�·�^�'��E��ȋ=�N��geL]�I��,���i�E� �0?��gj�RFZ^6}�������80�7Rx�����7ߎ]��cT���W��qSV�*��C��{! b�af>��n���"P����Z���=�4s�*v��,P�~i��M%Qg�
qSKP��}9��}<�iʫ�'[/ >�� DZk����L�7Q��볢;)��ģ��@/��0��s$?A��9�Q��	��^ٻ�7�S�TB�dݝ�;n�����;�����S�����RgԊ�I�]:�ag޵M!`�N�Q��wp�_�3
������=��J;#�!:���%�%���դ(m�~.^�uB�P��B�sN���oA�3����
������%\dB�\Ew2��Ќ��܃M���c׮�(��hQE�-�r�F�6��EQ`g�D��t�)w�s�t�S�͐G;^�>�ʦ ~SF7#��	/D�]̏��5�ʇ>��hM[�P	m��b �k�E=���x_��b��U(�k�*�C��Y��K&X����� w���O�ڒ�e�1N���db���@�$�y9l��n%� Mb�bf�0cW2e�q���y�sZ��>a���Ǆߖ�-f�R%�� ;�?C��j�!H��Չ��YJk��=Q��x���T���W�#�8�ذ��6���X�]:I��=�:I�g{fSwa p~9$ǅ���B)Ǵp�TxN�&���w��t�s���#��Wɾ�	��G���21�]�~x���qJF����¾���g��eQ���2OXnD��tS�����1�`~M�3�O�Z�Ee��C����c��S���[�Ls��7���������C����fEgy�k۬ !�i����	�o
��'wKP��f�����i�6~dz��̶z]��}w}|Y'd�ciwME��r�m��]UƼc������sk��_��UG!�8������	��Vו�%(`��.�$��q1P d[J���p@���?QKXp�ֈ�ܯ�˝[���ߍs48��-�����׏TBMw�����bc&5�%2g�mL��p?�)����x��|֟W_oy��Y����R����È/V����V�à4����C�h�!^V�Z��]��W�{Af1;@1jl�HIm9�^���#`�����	U�����Ƞ�Cx5Iר¤����c�������@��+e@+t8��i�����ҵ�;�@D�)�7��9j���Ke�QF�䢤��%����3E�?\@]b�8 �
���_l�C�+�kU3��T�K��)���p�V~�����.g�T�g����%&�T��Gk�`a"N�׃.|���?;�C����^�NOE�Tkc+	w�W,���k�)�E��+�fL$l�xfʅ7q����~�ZԦ�|�0e[���=�;��@E�/1��,�b��
ꆾG�8�d�u��F�~	���<.���*@�[�~Q@#�֎M��8�O���,�/U|̥�
a��K���5�P��Ƽv�R��kl���"B7'���!�jk^V��W��!�4�����[������W�b��	u��R������%�x������Ȑ�K�`����G�S��
���ߠ�V��r���-'�|�.���
��T��sI&��癅�F%^$-�dO:E5r�b�D���=
�sl.�7Ar�3�e|jr�0�E��q]��d��|�qDՎ|���:0��t�������5�����0�SGvy憙���H1��hJ����"ሡ|U��#�S_J��k/��*P��m_W�1�W@I��6��a�Q$�Sg�;fT��R���S"�����*��}K���#�ʊ����_�A)��f^�?.�lj����%�ym�G�K`��Y��	'M$�01�sȓ�]f�l<��4�36ܿ��e\Ha;	��,���+��e^?��Џ���X�V����y꓄
eYq�	p۷s���m ������5{���8�_j�����V��/-�h�nl*��ɷnvU�C[0�?`��]�^��GΝ�Q�\0f���l�T-h�q���b�4Lwc� C>BKЖy�.��S�2��K)Β`�� ���^��2�E�}�e���X/i��.7Vɍ��6}�� �vC�v� 5�:���ua�'1�/L/�l���Q�������J���^�z\J,	��t�l�,�i|� �
��ͦ��h�,>���<�7JK��Nv^�ױ���g��I��{}�����ץM��'wP�J(��o��N�q��4܋� ��/,��0d����˔5�gӪ<�8���ux"�������~� �\�B9.���-�N۲*�Ա��Ҩ���o���K�si��yy�s���3d�~!z�����a�wQ+��q`fx�*R�I϶N|Iژ���.P|��i�+���_���O!/�=t�=O�JjuyU1){�)!ݍ���Sa
��
�K�+�%���,G��ma��7>U�VJ��![w[p������=b��i�X�R1�+x��r�8����B�{Z���� ��!�LzM��}�0� >;��=�c���lI����/��뉁̀��ρ3A���|H9\��0�+��I����O���s�F'��k��=�ږ�/�z��ԉ�p�z��>��0�6���w\^�� � ��r����S2ό�"ey:��7�/R�|(C�-�)X��L���VK��o����PX�\~6�����^/����Sp�d�Oơ����泹ǿ'��o}�\~���z��?1pr���7�>�A�Dit9#��H�T�N��oKO�E#A#ͫ9�G��KM�f�y�gH;k>�?��hۙ0XQ��gd���s7��J���<b}��+�ҽ�;?��G���ۈ~ҟ{�3��}'S/�e���
f�v<�ٖSp��q��Ն�"ٛ���<�T�>�� �]��"��L��ъ��'�cL��B���si�Y.&����$���HT/�9v�����#���ih�t���kK#{z���n\]�;�ǥ��Y�I%:�.`)-[�7�4D��|�X24�[�����kZq�\5���03�j���"�?���gWi+�e.>>��A�ў�:�5{:cf���`Q.���'��78zd�j8D8O�ul�sS�����R�y�^��X�q��č�5����ڽR���:��̰�@dS�rD��A*J�oV=�$h50�g�����0��RF�?#SG���;6!�.)L*�ģ�J�jEt�˙.�\%:�f�*�2{�;������/F��'�[�O;����%�{�;���~����K�V(e�D�Ȧ�d?�Ng����Y܉5�Q(�eAdf��Ldd�3���a~��)䞓�d���r� K�Qßޓ@yH��{I��BS��J�t�3pP0�ɫ�~;�(k��3�>m�?�c�Uٯ�,����x���彎?���&��q���!������+'��m��vk��,�-��^���m�z� rP98��xY7=&��>]�����Br�]獅m�)�����Г;�d�a: �����Z�.��$��-O6�0��)-Z��'v�NHE3j�Vg�R̋6��7���K#˼%�B=T��̉���f��ݶ9U@�66|#�D�U��Wdjms�K�=������1�%r���M!S��Bְ�=: �kdHJ��}���,<p4��'3p��Ly�tl_v!���mF���61_.e6��e0�RJQ��9���җIW��8ߤ�*覤�؆ЫW�f���	Xe�fY���M��8S����(�Z�Y݉�֥(�� �������Ϭ��HG�O!AX�h�0���vi��,m5u?�-ߒ"�s���K���}���/�j�]V�c�S�o+Q�#�&�!Z��W�ڄ�*x�C���� �M�����ɿ�,D�-L�����Ns��j�av�1���	"�,�\m���H���x�B]�Zִ��H��2��w�K��=�|�y4�~D�2��\���L;���ډk>l�Y{UU�j�f�۫|�����/��a�e����0�P��PCV�m[�ܣ?m�E����$��JC�l�dW;[�}�M����ź����W��]+�e��*����D� ��:��t�G�_i���0��
E�S(OOZf��2�Trt~F !�ù�9�[)�$��Yp2�)�X\�6[�kH���������dI�h7!����@�P�*f\8'�Rtb}�_�W��A_���<%)D�$|R	���C���ha�a��d�h ���w\�Z��2�5�k��I��q�����M��z��k2��z��u�W�FZ;�oj�s7��9 >. �� B�L<G.�����K�/	7	�~Fp�A���$!m��HЂ;�k+j���#��Y��Fp��(�Lo:�����W�r�MU�k��W ��k �W�&��VمO���:���ϗ^ƈJ`�"�?�I��D�id}�O"��;�^@5�l�rm��|�@N����
b�<>s�VW�c{���50	���.,�%Ʉ�Vb�Ymf�F�&^?h~���=^��r�*��p	A�{��k����� 2����G�q׸ ���z74���'#cӭ��)�L7��R������S���@�����_Ȅm}귅 Q��s\Mx�OFv:}A1�K�����]�T��Z�RHjb<*sl���� �x%��Ia:F͚T�Ub���oa�2�n�"3��aPΌ���rN��ձ��od>1(	�����u��2�iv��D�\b�4���kmgUR�0�O�0b����d���h4~��/_�/ʢ�9Q? �Y�B� I�22�9f��(��>��3���
�����3"O�nu,�'�i��ѱ]Ȳd�]fiLN��)cŸ].{�E������ɘs�/Uq�����T��`Y/��������K�_D��\*!���	�������M$�d�CN0�"H��D�"��r.�o<
�	+�ȱE���l�;=��q&�����"4�.W7^V���HK��'�"�1mԴ�ŤF��31�G����nY�!�4�9D��26�|��A��Q��u�)8#�w_�F%���x��ͺ3������<��$��
�A�#�t��b<�-) �1�����6�)��0��Z���[,ٌ|�R�;��(��Wj+[ ��7es}�'%�QFu����*�H�!��)�<�_ �0�((�ϱ�N��Ɨ�j�R�6ud��O�t:o��e=S3S�����>7O�!HA��!Z~#ceĐf��C/E�	Llg5��<Qm�)�b�ָG� (�R���q=���ѩ�0t�]��хF�/=�n�e��ϡ���YR�I�=7����Să�/*�	�n���r�P,�a�����D��eD�De솫�����/*Q�oV"����n����]�a2!�?��W���d���E��ɳ�^�xYq�A�!�B��l�/X��aS�����4+g�p����&G62�G��]w�ej�(s�x�bK��Cx���|R��C� �~s��ǻ����9h!u%?3�֐�ӟ�IJW�#����,
�tbR���L��;�/���	�rٗiݗ�Bpi�[^(����򹀞�R���� +�r�����M�l�&}Zcx��QG�[� s�dp����h6�&�kr椠0�XD���JU���#X��K��6�ۂ�O {g���n�n8\>����N2����@�����$K=��/�����%���5�����m�{� h�ghՠ�(9��&�^ێ\Y����=s􎹜4��_��	,����}��/���o$����]7�9�X�#���A�<X�$�r�=|U�>��0�>�L;����Uܟ��!��ceդ �S��P��W��V�`+F�����ӻ��oN
��h�d�˳�jHa�x:�F	���<���l�K��&�Ѿܵ<IExz�A쵱��-{^����(�n��bc9�+~}s�O�%��V�N�{"�|��%:#|L�q��} ��]��=��H�h����C2Ⱌ�������yP��ys�ik}�z����9$����ӬU^�MR�C��g(^Mh��/�㎃�!MG�6�/���A�QY���?�2���@Yk*G崋��4̈� R)`������OY�Ċ9u����g�Y���ߨ�Z��D����D!.=m_��vɁd����ϴV���t"�B��T�=M �N���g����lfk?B]�1E}���@�,$�N�?A�y Q�Hi~���$C���J�jH�M�^�+
�`�/��v}f��ŗ��g��~�0���˶\b�pf%��Rz�^L�Q���5K��Z��ל�f�y� ��H����n$:16JFL�,E��oЈ�M��H�RJ�I��+�^���&��q;c�2mL�2��i�J���CRYN��L�j��Ӷ�R�"���aGP���&ve������1�v{�=��m���
`ߔ��!�H�S�c��zI��.��.���r
��6�^/��YUG���O_���}�{�%���5E���{��:Om q�;y��d������P�A�增������qűϕ��������U;�{U�(iq^��Kh/��WU�}� ���uMBa4j?��2u[{e��ѹo�q^�"8���M�z2���������T2�U��U\��%��1���7�|��r۔���~��4c1�}6��%q��ބ��s�y���������~
,Ҹ�����܌�����$k�t��.�Sh����PG˼(Ɏ�A���p{��7A��e��u� _��3�C��Lq_2��!J���>j���?�zf)c&���ʪه�<��8/d�RM�v3�v�*{B���_��0��MR,�t�ln�i+��3=������]��&G65�����@�}֕��0i��B��7Q3�4�!�n'���V@��K��B�C'F��n?Q洟����I�*Q0axUY)�L�����!K�]�k�+#�v"U{a�u��H���k�C�1��n|�����i��7�M�Ũ(������&[JiɌ��������3����5|��MD�<+��x\"f��K�$pG����BŇ]p3�A��Կ�H�:A*l]%f}VX�4%�=ܯ$��հ�bƧ��0m���'�Ь:��w��hI7��ߢ����Z�'�)��N��n��JE/��\֥I�r�>0`V�IPIߚS������]n��m�B@���TV�Q�C��
�H)��8yS̵H"�K��]�Nc���i��O�����U����9�µ�����:�9d�h��D���4�>��}TZ=!1��Sg��J���d�"�F_1\� ��Kb���n� ޶l��.�y�"lUh�hF<_�����=�eюE�2�s�~���I��BH�	�b�ڝ�Ҡ�+yO����Ѣ�JS��;�ǔ.s�U�տ1�iKז{��Z�������mF��6�I�Fw(��*t�KoZ^W)Kl��F�c�*��B��c���A�ft�pr��տ
�z�@��02�n.��X_�p�P�c��w��s�}}-�e�t�0���"�9}��C�3ט��Ņm�(��{��m.�87�e!1ÂR����g!��'���T������J�r}���C5B�[��mQتg�a��8޽ѧؐ��O���d�ns�$r��٠����O�`�N�R}%Y����g@Tw��Y�]F4˘�Χu�s�|C�7:%�����O.����������r����Mo[˲��Ϥ�_��rqJ��Vi���n�0
B��)I�?\?�:�m�4g�v������d����F��1�4�^h�M�!k�k��^�dȑ��ە�����N���i@��7p�8����G���R�#��R��U[.6ALMo��Vٔ+2�X�G�ú�3ο���yD���rEڊ���G]9��,����5�!��\����Fc�P���z���wFC��x��zhW�*��HC�规�����,�p�Ƹ�6$�6Rݛ�@�@hO?>u%�{�7�L+8��$h�����k�:��I����h��ٴA�?��AH�QwH8��uNJ��z���1�5�Z���R�
edqI��A�&j�
8C�=��e�-�lH��VGRa��{b��JK�'�dҿυ�S����W������&����v��n���|�쏮�����|af��fW�$c�mj�C?����T�� ���VE�&+=�<>�'���`�C��c�B"c� K�B<�.�=��%������R�˯Y������¡}������kj�7%�"�'ـ��|��8����Lo����Mq~����,�c��VQ��n�^��,&�̽���+�Ou���/Xњ�T?�=�)���7���Z�KN�)+P��OfDPm*k5'D)
�߳cE��0W�Sw@L@(��6���b���ko�nH89�|�Ik�l�z��S����pɫy��=C�TL�����>���6Z��(��	�����hB���N�1�Jxs���ɠ&E�o�N��*��Mq��H�����;a������E�?�IU[�����'�Mv�G�~q���t����{��Q�'�v�޽U��0�*�xytų7̆�D��S���}�/߳�����όд�%��q�V�w��O�-3q��S���nAv�#\�u�5�%J>z�Hj��6K���K��'��J����E4��e�S�MԄQqަ���+��r�r�b��N��4�čbi�f��(c�F�շE�@�nNn�o�[�Sh���`�i�t��2kOxA^�>�~�P�ShlL2f���ah�؃�����揑[�Ԓȣk�����"d:�v��|TJ�y�������B5D�BH�PG��
Q��Q�Z|�x0��=�'��z�S,��\^��]��F;!Y��r*�x��*/�~C�<��?}Y%t�t�����ļ՚���{�>� YN4P��]�/k� c������T�ʑ�_��2� ��9v���
&�
�+>����*^�TӶ�J|8k���C/EP�-PSkk[�H�n<������@�m ����mR�W��"FЯR����7�*�φ@�������'�|��n[��_�np�"�X`{;b�g]�������t�Ju��v\�f��M�]��o�H�r�����y#V����f_�p;���f���M����>1X�|eFL�-[
�^�7AA�<�2��O�n��]���m���@���芑���� 0��Y����q~�U~�Á���h�v@�M�׀j�͢��;�H	KyΚYeEg���Y�O�>pMu$�/a�#�4�|�mG�QbEY�x�����Š�O{O=k�4o����ԟ�����n��ϫS�*��Jy�J�&u�z>����~�y���S��v��L���=��mB뿤!VF _����(7�.�W��>�f=���CF�8���e��
�=�}��j��'8<,���z��R<Dc�B�.Lj���*Q��Ԑ�a���^�ѓ�-Cm�Z�Q�ز����V�x�}�|���y��+Ab?�a�q+EDl��>�*��?�M���$�� �W[�5�2�f�g���q�69�|ǐ���pW�`�M�?�b�^��`UY%��R�]=w*N	~t9�Ȃ�誸��(�5/����}s'�@-�)�mL����
�4Sk!-�;KV���	��C�1������K�d��d���3aq�&��˨�kS�Kۚ�DvP�H�@V�x��$ �bo��V}��g�Ҭ���X~��;\��Q)���;OI<@����+���'��ܙyo[T5�bbKn�w2���;Ye�f��3�\���m��X���U.D��D�������XT�e�k>03��M������p�O�]T3��
=�����p��Vwx#Z�?̸���n��w�fnLKg�J��!�ŏ��2��vܗ.U�hE ����W��Z�W1�Ju�|2�M�D�fS���T�~w�z�.疶��g�Uu�G, `h[��=���R\���80�j.�|�rT!�r+��x�v�l5/�}�_f�x�1[6ǒ��h�H4��ie��L���/�9sG&qM����*���k�Ϫ��2K;@���ܛ�n�4'c�cV�#�p�}��!�����D}si�{�{���Iɇ����e��pB��<�U�O���5IYߏ���b�.�2�&���7���7��p�(AM~h�ړv*�o�MG]s��-h3}�����c�Q�cB|�k�>�� H�����$!�aF�4��q4��[	�짘2���%��yϗ��$9�r�.SOB=�rI���
�æ�g4�1�w���!��e���3�Yq�+:��ӵ��&����)ARQ$�Dzu�wk�2\�������6�v!����/��;g�z��L�[J*���}Gz�����N�vW��,�i�� )s�����\+�����I���w��3�n,^R����UB��&9�#Z�,{/38���$�o[6�<���zC���E4��y%���n��[m	��bhË� �g�!A�gM�	icۣ�6c	K���!���{�	�[�V3sTV��!��@TUD��J����*މ6��~��"U;�w�^�����������Y�Őod��LD����4@���`��ű1̨x�6�6MU+���É�!�����*������}@v?��>Vz���L~@�&$�!3�ϛ�0���i ���?�b�D&n���Kų��^��~t��O�O�_�;>Ԍ=���\���h��;s�(Ʌ
�6��9K�ny��Tb�u�S=�M����z$>}_O�]�=�xs+�֏x� l�:��u�/뀷N���a#��>�x 	�h^�@���6�RU��s�k�S�C'2��������3���$�1)i��]v�����r��r3K���rF�6�ި�g��s�Ω�5���,K\�r;�l�7��h���e$˩��T���"�jI|�Uл�/���6\	?�a-*�Y=�޲�/����iZ+$�{IȘ������La�^pT;F�+&L��z{9�G����܉�F�1Q
�Xxl�Bp����Cu�9��D�F�{�=� [�(h���� IG��@f+>���Cq��N�����3SI�s�ϐ&
Hzcs�+B�Mo�&�� �Y#�r�fX�[5S���س���4���&���U���õ6�D��`Q!Hw$B*S.�S�"�P��$׳/����~*0}��`�e��x�9�3G)A�����w���Ux�ۇ�n�)A�a�:90�ӿ�%�����2r@Y]2��0�v�u��4!�*-]�#�:�L��Y��I�N	�;��-(2[q���~�7�����?.g��qR���^̊���:#������sm�Oq�@�s�I}���]1AN���R�2T,o9���/�1mF8����A#����%'��_>��r�S׌v��Q���-��h��m�K��������ݓ�`���f* S��W���:z�0��L����5�����S��ck�����(4�GC��Ĳ��%ѡ��}t�o�{�Lq+��xP���eF��b{I �������p������7�S0v���5/r��(�!]� ��޺��f���E@�,��%8�榚��Q9�?U�Q���0|6x<O(���5r+J���u�)�4��'N��H$0�e��@5&aT�O*	%ǁ�v�C�H#?�`�64"��3�gvi�,��K���5��k u���zb��c��E��3>�?{�re���a��I��u9�º>qvj�:�z�~�
.Id7����_�=R�F����P��Kƺ./mI%BQ�@�)�A�.�>��ݤ".]�{D[�'Z�35��-ë�s���j�Q���D������.)���`�5�e��G�㿏ȱh�5��|I!�`o<5�� J�4�X1���dw0/V�r�Z���~.4hr����ҿ;e�º0�4<d�u�~[�����]���~	Q�^�K��Ta�+�}|"�ig�
hYywxiK��/����C�n/\9���h�2���P�s���C�i-�iY��9�I�&�i��8�kZa����|��=@3:���0CID��.`�������h��I����ƈ_@�Je�Ohw} '��S����Z�R�z/&Ο�m�����D�*[��zE��aP����C�Ѕ~��%3�ɗ�P6���R@�Sҙ�d�*�>Mw��$��:뾟��OC�E�<���������\i�o/��4H&����ߎ����G�R��u1��L<tz��0  5�2�0����m�0����VD�L]Q�P����)�f|Ԗ ��� Zj���II�U�C�Hl�X�<y�T���#9��z�`��&�ay$�)5s�C�@55Y;��؊B�CO>"Oـlˋ4!�~ɢ����/u�f�?Gk�`(�����1B*dI�qCSJ+j8�)�םq࿲֕�ִ�YJv�:���+)���G�￩go�
Z'_(�~�v9<��~5�?�j�Ȓ ���˫�A�TA��\�����W���(�e��/9M@��e��U~*7����I���9��q�D�$�q���*�v�$��ߑA�ry\�4/�:������]���3�+#q���nz��%�O\��UmN(���ne<��������!F#H��P�0���aVtЯ�B��<�zȆ�vq��i��n�>����x�T�4�J�%g��a��0��lP5u0�#���h��5� ���O��u�ec�����#����@�%sWP�r�X�NG�@���~pZYyt�hKQ�T6�5��͆��}9��E,�9V��~��&��C�S�z��ִt`��X�f�!�qBy�����URqC�	*��,�ld��4���O�}[<�BKF��q-��!U��Tϕ"�H8���J/?��M����`Jc�7�+����3���ߜ ��n�{|�E܂d��������8x�2 �J䙃�?��o�fh���_?乚]�
5掗Z�biB�u�7�����R�j�1�H��5;:U��B�1Nf~`��
ˊ�S�T����R����F��O�~��yW����f9���GB��ؘ����.���K
Ik+����'�U�z�a�1sV�x��
0 �k�����(�0kG�6���2�
�GX�t`�,�o�TS	7~�����@ø��v
��Ǒ�
��r���\SpJ�}�����ܺ����F����YK� D*��4x�>yjQ���Ӵ�<�iR:r�Z�_K׮��y��Zs.�7�������AW.(Mi�/ny�f�J6d�O�Ɏ��3��'%рDk���7���r�{��¿��v/b��7�IB����W���7M���C��FU��Q���`fAJ�%9H�~MX�r�f�Z}��*K�<:^���I��#lG\@}�K?;9 �A�/9�XK�����iy�MncF2b�(���fqb�@�����l|[o����v���A׆z�}DsKa6i�0�Ѝ�$�#_Г紋�3�ݓ}��70k$������`1%P�ko�+!����w��qֿ��`�$b�d����m"�]#g�U�%B��a�Jm���kP�X����^����/�q^ԿK�2C�T��!q��������&u�%�t���S2�/�7`���7u����5%��0����%0���]ת����Tg�&�|�����
l�`��Ќ̶�ܵ{�t�w��
lN�/g0襳4U,��]86d@;ٝ�ӷ�=�ƹe�v� ��k����z��k���b�_Wu������RT۴�x�h �Z�����,8�u�����l�?K���B7zbx)S{r��Q��)�����2H����u�j�$i�$�ZV�İ���2�
d:�u�й�_O�\9I+�I,M �v>#��/�M_�ٹ$�2/�C^������F�?
�d,H��oDcY'n���U��N���g�KH����B�\7 G��zN�+�y�.���蘉-�l0~������Z�xy���i����p@/S�V�jA_����q*zu��t�p�:�� ���%<5�y���)�P�uA���=�p2����V:m�ޕ�u79�f�λ�]���sw#w&�"L'"X`�q�!}6�p����#Y��?��f�V���E:a=��N>h ��w4�F�d����$�".eˌ6H/�g�#.h� ����0Ȫ�D�+ݙ�y\ɘ�v
����Hʲ�fܥ�=oʀi �z����o>>�ų蓗
�O�%<W$��<tM!uo|�3_��] 4Ԩ�������!�ca�Ԁ(�f���N�/����(�h��!���2*�Eb���B���3�hd��<Mp	@��kJ��R��"�z'֗K�/��
�(:���T4ջ������ӰY�%-"?�o�%6�p��n�zO�v4tN�v����`k�L�0ω���m�Дe���z���r���������E��$`�U�}Vn�`�
.����]F4�`�*4|�z#�h�P�$.��~Í��>Ǫ��T��'�{�[6U���*-���O�ԕ�k�dE��s�	਎�VI���|�ku���ʏ�b8V¿�������>g�
}���ɐ�j��m2�r�Rw�8��k"E��mիw��n �Q���q�e�5�t�9�?�p�I��`2��$,�3��*������>3h���{߿�%�~��T]Ζ��H����jp�P�8�+=l���Y�-w
!�Wq��)͛X��ڐ2!����3943�[7*c٫�\��rE/���m��,��	�Z����6!�-9��+�j�Y�dR��c�fo���0�L�c����nD�x �L�>�����*�*���+�u�4ƺ���N���g��c�>�_ǖF��\�[�([r��$)�T���%v�H�+��Iz����9n
dP6�DHA��P�3kοl'�D�����FZ-����7LI��z����.	W��*��eL������p��jxo���`�s!O��ú������1߂��6%=w���z��Ẩ���t� ����L҆b���OsT(.3������W �Aϴ3����0-���bK$.�iY�:@��x�<Oz ��n.�'��֙J0�t��?}���wQ`�
s��YR�"�Ä�E�V3�gS��� �G����/��	BB���!嵨[
w�7����Ym�jDK��١j��]�s�ğBfJ�1��)7/("��9V}[uK�tn�r5LeTHj��V*��;RXx���G�u��t����(U�Ed��R}�Qm�ȑ�W;�b�H�:G/�*�7��<�lM��/|�Y������U_�#�/J, K����Ĵ�F��-�X���/��{S��ȉ�4G ��ϋ42�b�s,�rXky<�sD�kݬo�t]�)��x��UQ�8^ٱ Rȴ�I5�r�=�a��^�-�+��^`��/Rٰ:������A��kE䒣
�4���s��T��X�Mo�,�==w������'�;��>�q"0�m���n�b��h��P0I��+eC��(�mj+����o�G��t��<Qj� h.�rT6�?4�7A�)���e��O̺V6�w7,������j{J�_j�pG��ŜQ�B[k�'*�a�r0&�q�ҏ�+��Î��r4<h�}d��Uŭr��*����F��B����x�6FH$~��eg�M��=�R J��G�P%���$*X�C&FH� cv>r�W%�tZ[�.q(�A��ay����-b�0"x�i�N����t��$Eb�{!b,)������eX���-Aa�g�޳
�&�����\���D{;�)��TDgoQ����� ��W/�Θb��L�C� �C���)�\��d.
�{"Ba��!�*� �E�"����S�t!$_�Ѿ"��#n�0͐�]����+{vx��1��7��w5�����_�(9ǐ��o��<���xur��g�������eՠ���MB�L+ɝyB�Rf�*٦t�r�nV@J���m5ُt�Ȣ�3����C��,�+5�	��ݶ�x�p����.��y֞d%��+��� �G`ؕ>����`55���b�����8��
��P��#9�2y����؍���ǆ�horN>L�XM>�������g�<�>I�Ѳ;;�3oL��Gq<�qq�@F����G����CVfx_��k��.9�\�A_�~ݿݐ��!ʡ'��m�W�d�Z�u��H����c���6��M�}So�mPJAp�^�I1
���H$�@}�k��B�Pb�W��k�J�����M�:�!�"KN����&sc�iw����_O��$5�����!.']��孾^�����.7�c�1�5oD,]r��<�?\i�n�7�N_p��A�j\Y�ފ;P��v׍��ƙ�OGL�()W+��F��v��끫V0SR�L�N�gGGkg[ji#��"&'��,�즇�o'���x��5�b�D}@���߄9�V�Z��4O:/L��y%��[n*�x��2�)6#��ћ$\��1�l�z����>Q�j���݆+��Τ���!�)7�uWva��V&}�-���B�jxIB�s>DT��]��qKZ��bͽ�&��;��1�/^�"�� X���<F�o@��uބD��P����`RCE4e!��SgP���vaD�
ց���i�=�����O���R�O�P�#����O��ɏ+g�=������wɜ����Օ!_u7�4��$�J�?�(l�Z ����W�.�[��a��^�È�da�2�)�`�={���U�ˡ�U��NG.@+_v��h������!Ә�{��]Ez.���N�*�^�^h�l~nɫr,4�XD�������D�4:��aM����s ��@� �m@���_g���V}�p�M��ɞ
i��+X�Uo��=C�v)��]�ZD�i��W�^L�n�%P{b�2ǁ(�^|��u(Z�B��%����]�^?��{��R�e�~�m.6�(�o����`]�r���vc�i��+�W�j�ewh��c���C����U�V��1��1�Iӯ+{#v�Q�.�.)���䨍� ��<0�R�l� �f������ׂt�I��R��I�j)Ģ��R��r 	 lܨ�i_#>`�篹~��v�yċ���E���
q����.6�uk�� �ɐ~���M=��C�{��w��I~��Ho���KRw���y�����N!�ePi|I����J1Vۏ;|�oȲ���E���<����8P-��nή�$�<���a��լT�O1*`��	tuj�, O(	]�
~;!:�u�r��C޳Hl��\+�lty�9���	��9�O�?	^oA<HV܍5�����f)��T@
X {�2!(�}���Y��vS��Е�,���1`¹/L��1m�+�J\>�^�)�W&U�W������V�ϬƘ��i�!����9>F�UH)�?f�2�)�z��kM��Iհ�ɵƓ:�8��|E�Z-\��]cu �)���23I�E�9�u�?�T���<Һѣ�ܰ������SO�_ȶ��y���ɺ,Js`�=�L�ڔ.�ս��=+Im"��D�|o��%99��_��i�1&�>�ԣՏD�O�EPCA�T(}m<z"�t ����ǁ��#.����%<y6�#��л�EC[��?���E��b ka��JR�/�OT��n=�Rt�ѯ'���C?a�����[�h��D�Q3ܝ:N�y��(��d�T��*Q`jŅ�x��W��`��sc��&����`�����jG���ձ�!��2
>���<ĳ��62<��o<Dto��*�d��nUk���Đ��i&"�K^ �\<d3.5}ý�g�l�y�ݼ���ۍG�����x�n�qB.,��AD@Ԉkz��=tO��0��Y�^��Tހ�wU���Z<?Q��I�s%OX�������<�@�'�~'V'�`��QW}�4�w��3�A ��w��U��$):+L4��Ѭ�	h�Q`ݾ[�UB�/y�
�ϿK����#s�uL!�Q७I� ���Y���}�@����<F�F�=)�@��Eˋ�8������l
��Ɔ�é��<�M*�>�3Y-�@��Bb#;����A*�є�`����A�{�L�§ͱɫ��v�X����H�[��W4p�^ⳕrb����!.��˵|#}�?0��&zri �'ȉ�,3�h
 b�r"P�=^�]l�2Z�(�{�R�
��u׮f������F�tcC�Ma����f߆�u�>(�p96?#���4��f����ކ�΅A>���	<&Nϖ2q��RY�a��4^���9�7����:�d�y!i���|���@n�j�\�~q�PlЧ���ÉE���}@$s���Bv������S��i�S=g��s|�	透|�L�\�r�p����_U1�#8�&��kbM��
�p�<'�F�@����-"�h5m��v>⻗9��~(���bg*7@�I��3��5�����^(��x\���9[p��Եz@X2�
���w��68��9�۸8�'���_�W�#�	59p����z�L�Z���.�L�%p���qzÚnEj�}��+h7���9V�iCk�~T1�i�f?��o�1=�~I�(n2�
6�h�"P���cK5�9�5$�|�C`)m��'h�:6�cR�cn�Y�{����`�.�n҆|u��jb�v;s���>y���ȥ�����E��@�y�O�ʟ�0��;����J�F&Uj3,}�����p�	&=���^)�
|�Yۅ���v/�������3n��a��5T��E�B]���:9�p�f^���|;j�W�rD/G��1.�W 'Ƣ~ꡆe�[�������������y^w��p��|��O۟c�?%�����E<tHU��9������M��}t�TQ?�tI�)s"���\e��~m�))�j���^3a�0?pފ��[%�=�ȟf�rh(+ɤO���F��k�1`X�2���I*����`׼�@�	�
�ӿ��U��C��s$$�q��Q�����O90���V}�w'1W������3ؒ)[L���f	~.���j��H'�By�ObE~��V�֖���H?�quE�F�����B�pR���\e�����u@�A�+2�K�܆6��h�g�,�1��F����RK<�[��"��#����?B�DԂj��s��QXd�G�Y�����u~Bf���hHC�)��A#6²O&������g��N`�)��O�����L7Hw0�qϫ�#� �|�y�1�~�������ލo���H�L�j�j��*V%�co�.��=E��Evq��=����C�.���V	~�����*(��u��S��<~���I�ƾf����"�=��*={��9d������n�r��l���t��LY�|�?8:�h��&:�'�!���{b�ɫk�"z_"*�H��-���g�$W�a,i���q� b��Eɏ�
�Vُ��؆�9�l�0]p�|晧�O*�[7_�nqˮ������{�X�#���4���]h��M�Jj�&��k�0�'2,�a��g��w��5
B�N��̊U�0M���t��N�C�a��.��Bv\+Mgw����X������,:-�J/B����Ȯ�Aw�t�\���"R�5��6^/�����n��<F�O�
�j����ǅ>#7��E��F��o ��e\J�����Y��1E�
������p�w����?�Ȭ�����_� _����|�N�lu��`!�LG���%Yy�H4��MXß
@�*���z�հ���bbE0���66�%&F�Q�~>�c�ݙ���9���I�J�L���/Zh._O
J�=PV��3_��tpԁ� ����~�z��fI(&�"�����rm��F?�����O(s���AR���ow�����' ���w��ȱBݢlQ5�Y�=�;]�
9(B
��v#9�K���)��5��D�Y.�*C�l�$�"u�V�X>�
����P�%��ˮV��*`��KK[�������L����N����D�nY�W��l��d����$���<�O�7[��x��f(�׮:	�\����ЌJtű~���u�x�Y��c�ˍ�����.���I@hҏM'�~D	A����v�xpq`ͯ�E��T"H�Q��Q��l��N��4�H�PPc�N�A��t r6t�2�$�1Ƌ�~��� s1>�}St̨�Q� h8QW���� �ꦆ�Nj����x�t��4mIk��E�x�Te#����U�7s|����'��DG]���;r:��%�Jܑ� p�;�t�\-QV��D�D�wZ��t��h�!��{G�����+�D�lQ^S����_������Pes��1� pf5
��;y��*#D�$$enj�hZ�~�!���:g����rM��lw�Š��mD��������L�3�Hs��՛𬕭�9Y5E���G_� ��A.���0������\���O���-ͨ�oY2K��w�"!"�����K�6�	�y�{��Eň��̶�`���b�8F��R�t�w�_v���z'W�B��7J�d�c��c��f�/��<��\Q�L����4D��������<�)������,|t�Ma"�l����I����������uD�	��|������/�XX��d��b~�vӇ�.'��j5�d}�Ȥ�q��M�����O�ʎ+�h�t�@�|j�w���I��=�4ScC���Cp
G& #��#)�N�e�C�ҖH�$	zi�f<�h�I�*��=o_&�MWh�D�>�,�N5����Z�W��5��C�k�Y��0G�Н-�I��y�K��rF�����ڲ��a+�x�=��q8��7B�U�;4��2�[�`�)�"��f��Lom.���T����vxW����ڭ��R1^��Щ\�ZaTΜ�:6/>���!�Y��Mg!"������R�ۀ\1{C��v(p_/E���]�{��l$f�+�n��_���%R�s3#"�9�[ �-!4�f�8�Ĺ���uU��>��I�⚗t�l�I*{�+�}�U>ꗄ��>2�V�`/���-1�h�F#�~��[b�8���ٖo��{3� �5� *YV���Qj�֚9�^�N��r��ܕ���t�{S�)��r���(�y�78�rɴ4��kI���W,fvyB���b�o�f��(�8�g��y-�	O�%��m��j7�"��C���qV|���E�(e:P��'1�-f��|��<���B�5Y f���%�/iG��-���U�F���8୸&�#��)&ˤ�,��sii��[�Wy�E�b1l��6T����6����b���lp$���j�
$��,#��go�*��t�.�D�5�ED�y�n�X��8��Ŕ��/C?4�K������m>ߴzB��aUK+)�F�I �1�^�����Z~�nC`��%�����)�P�c�J����aX�;���G�E.��Q�'��
��r�%�\�|�A�L�u��f�o�[���xjD���1d1 �VyӺ-��ic���m���
�w��
Ș=ѯ����7�,�+Zˆ�����M=5C�� �mvh;B�k�ֹ����E�&(�Pqs�ȳ%�d�M3�����S��iq���%gC��Y�]"r�w"�U�/�%��t��+������Gu���
i^̌���-�����xSY�� �DLEKk�%̣zbɵ�9E�u���i�2A��IxX����慢h�0�w���6�VsS�ǰ�K�ϙA���HU�{�i���0��e�*|��:.t��#	}�27��U���8�U:<��єA��U<���F�kwƪW���k�Ry��c-��]�Fk4�Ul�9Q b)@<��_��`8AT��I��>���l�cB��j0ifrX��}��)/w��n:e`�2�����z�Z^1�B�>UuJ�]����� ���um:J{6}d�'������Z�*2H�_����I�a8H�c``�Խ�T��jԇ�L�
��A�j@�FY���XP  ����H�aUE��2���0f�Ñ�"��NZP2��-�Y�P���Q6��52+	��G'ޓw�z[����n6���N�ԫW�B,�?5� �\���4ZU�?:lj�3��{+��lH�z���Õ�ARը�f_���E���4�%j�e�2������;����"ŷ��fS�!�9��ı��o�QK-����.�	O,�\�U�Ѓ���ˢ��9)g�C�_�	��~��D��v� ��^ef�S�2Z�dmjo����#�*�l�|D��:��(p�K*V��詯 V�6t��'P4>Ա�d곶����l,p�I7�<(NۋC4#|�'�.�#�27�;p����+ͅAA��P��^g(%r��]ȁ�،�\Y���-��.�L+Wt�x�2o����Z���ܲ �v	��	Ⱥ�涪a�pa�g
�&r����>K��n�Y����QR�eu%�>��$C�7���<$������m���.� ס�\��%��d.��k�3$.�E�������u�����@~��j`m�ml���!]�a�9��ʀ�BY*P�zA�*4���xt؟��Q�X4v�3����-�S��Cm��ޫ�������"���p���q���^�N=j�Ùa8�TX�yr��^���>��=�sY�5zEryD糩�&Ǝq���?��{��"��N��抸��;��w��4�4�}�lĒ��/�YE�����g�f�U��bԩ�S�0�MQ�H?�I�3VB{���C��Pgc�E�q�ͼ8��@f�,TH�	w_�u��Ș���������b�&�eڨ�?����.vKty��,\����J^O�!��Ԝ����^��ב�%2�,[�~�"C|c�m�hK~jZ��E�E����f	�nAt��[h�2��GO�����nE��pa��� ˬ1��D���ь� �T Ǆ<H��x/&�
hMۇ��B]�E0�M�gٿPwV�C��XP_.��ӛ�����D��󦝤1f�T��.�I�$Xɻ)%�RDs�o/��V��7�܋_ǄQ+��I�_�9%UM��TɃ�_�)��:�!E7��I������v��g�g{�nS�C�'9�q��*����[�Q|�<t��R���Gӿ���m���'G&����bQB����=$��noĨߝ����Wb��5cUT�,���d6L�4FX9�H���x�+���OC�il�m���g`��n.s�yn��d=���l��D���%���kb��z��P�
���ĩ����N5��-�=V��X0�>b��L�|
��+���v�2~;Ȕ]!��V��뻇d�$	�`���bDN��I��Ŋ�H��Ϛ���ŏ��M��E_|��|�\��"{���4��$�#�o��:��O+K���dS�S��Kmm��V%�~A��Qﺃ��_��l������a!��C����3ב��&)��i%�_�rEș{�=����=϶�f�]��kx��	���n�b��Eq�ېY��	��vRb<V�W�K���;�ɛ��d�d��D	rI<�8��#�:;6qUKg7�c=���f�����,�#߱��1���jLS&�Lp���aN�����[�B���BCp��7!�&�c��U�Q��6˚��A�R@�G�HTS�C�/�'��1����ZD����\���DQ�H B��4Z\*����OU���K{��zf{�ؽ����l��#&O�$)���~^�USds�6(x�T��5��$����{,��߆I��i���2ܼ���=���+�S�F�;-��y������{�l�ݗ��-����Bq���qv7�ьbߒA �V?.h(�S_�����P�&~�U�Ln�k%�J%|���U����bQm��Y2ܢ����n㻴Џ��	ɻ������{(��u����B}i	�!�y5"/�����$���~r�p�����IT�5ͣ����_�ײ������#�{�T�5�] Dd�V? ����#.�$?Pn�f�!���d4��f�Pye���'��3 �=EkA���������>�f/3�&�GR.J���{�P��QĚm�Q�wk�D8�d��8$Q�$�@��U�I�������K�Yn~"($W���c.G�L5��uí����6x�+�|�)dIQ�'Er��exI�+Ebw}G���hL�ǒلrP �⢯d	�}��]�U���6�_*AQn�5�I`g�eZ�\�O����SՄ�<{�`�	�1�41C�R���)h	(=��~UֳV�8�����{� �.����šƻ����	���$]���g������k��������2��Y�W���2։@��`NM��.��6�n$��$�6�JS��h[��y��#���0ہ����$Zm�V+��[/�����Q��'��	h�+:�FQ�c��7�Yn��P/��a����#R��2| �w�(��<��<�_��[7�
�2��Z���ۧ]��
���	�!���S��C�}�����`�7�#�{�:B[��(k��[Qi �Yy	�pƘ.����cf�{��)H|���H���6l���gP������=������e�[��l���#s@�����ń�}a�ȩ�k��b���J X�5Mdl�ǗЎ"�
��a���{N8�B��Z�+lj�R���n[�D)�Z31�fMwq��LJu��Do��TH����`9z3����9 �ImO�:����R�42��;���P�%��o��oUk&�K�M�T&?T�2�?�2�^�;�R�v�_��y�K��g�b�Eb�#d�����S/�}9�@�ŇT�#J�J6��*p��(�[Z�K��t�Ir1-X���q=`y#3�?�}f���'�dr!���4^�k3?�+�F�
�9�pA8[qH��N�{ٛG�V�K��;�Hg�	Ih#�?̡�}����Y�L�;oז���j7c[7:��(�̑��eݸG�+٫rC7���:_�w���E#���^_Ⱥ��]v��|bH\�̭x6B"uÄ+���7:~��b Y��W��j5d��Ss�⬓�5,�bY��p��X�+�&�w�$�N�i����n�B���M�UX*|��v�c�x�s��[^�S:|�������)|;�Mr��MOܯ����(��a6?v�J�F���ӒW�%u�#�ICFsC���-!F��]���(�^���i�f8�Y0�͝.2R��)��#�dk���/wR<SG�V}O@���)pS