��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>��`HX����5a8SjfSު�U��c<�`|�g�J�@r��c��W���J2iO���7���d��t�#����3 �SF��%u�l�×ElM��{i��O �cZ c�R�����+Qn�޻�yv}T�m�O�D ���@.u� �[���@�+%9�Yف���y����&_����)���JH�?��mh�If�o��(qZ����E�W/}���&+�� ����F�ɧ�a�@���	��S�/���Y{�!҈�2�>Wh��������O܏ݸ1o�&� L���By��;�0���ŦO�E�5��Z�P:rJ�
k f���1�Hi�<�jfF'��ے|�]#^8�x[�x$z��rn�h�[�a�Xv~>�@��� K-y\�f��
i���Z����4f�n�O��'3[���u�:x��#���-����c��p�z�!�J���"�j�}!��Z�b�,���Q�z�,�'wFT�� �g9W
r%Yrhq)]��`,!�ep������盏��/���K'��L}�:�a�:dl��#����-B�������BߵG��Jecu�Y�IV�ԋy�G����'�P���ٜ:y =�
��ǲA��`��ɤ|֋�W�%Q�`��t{��
�X�O���v�_�h�B�����б�;B�e���@�n|b<y�}�����.q�3K��=��9��D�e��<t6��ibq�܋h��6O�@G��VE�4����-�|����-ul+���a��1._m����4�5w��C�o���c�P�-ϱTrT��`��p�m|�S8N� �Bޓ>�y\��9R)
|�m�<i�s���>]{eA �L&ǲi�8�&��܌���b�]Jr��:�h- ��xs=������O�"��ݜ\E5�[�	F�������#�N�[��;���w�E��_�+i�x�4����BE�_�������H2<��x:�GC�(��u�N���Q���J�W;������m��(~VB������6�r�$On`�7�9�(�̫���8�Ġ��L���>^CǱ�%Ƶ�����q~M+a?�_��?�<rf4$��us>EV�6�D�9RMf���~�G	����1���0���^?=�Ȯ�4���:�8k:��B���{���t'|g��!>*5t��#će�F԰&�Rh.\�7�˲i��fJAfR�O0���}�g������@��-�X��H���̞,��$���:{Mw
{> \k���V�I�5��Θ�-��QC�!���Zg��j(Z��yۃB���hE��1i@c����)�d�G�ib��V���EX���c�**��fl�*����4ca�����Ť� �;z�d.G��5}�[��-�}`(hДPv��z�������CE�mh�7Ayg��E۸I5�{
ϕ��{A��8�ǬXː]�a¥#}��ה��ҭ1���:����j,�sC�O��:�BP-J(��.�B�4͸����t��N&t<�#ܒ�Ɯ��<7��oIeT�3)��t�z�����bm�7��D�:b��^�FÅ��T{���L8�f�A�-�����Q�
?�g�Sun%�`&�#�V�����}Я'�K�^"��O��jomu�h������9�z��)���S�Ƥ`�pй��XT5�
��'��s<�O�]��5e	c�]:џ��&�6��;��TkfW��e�9���Z#th�C]�T����q�U{�o�� J3�;`C҃�u���@�{��_��M��z�n������6�{����i��NKjW��W��@4C�v2˰tR�T������9-,�b�K��'���S��v}gQ	��T8lǏ�%yr��4݀T��sT.���N����ݨ�3�JA�T$��+L�|u�	+ӡ|G�����>M���0]�Ԣ�E���"���)~���XK�|¤8�]
?|����Z��~T�����{�3�	5i]��yX�Jf�	��'xF�¬��C�}��d8����ޑaXo���c�J�eod�I�=h���V��m������@W;�&Q#, �,qh��YD��	��%)X2G�W1թ����2�16TQ�._�Ʃ}_F���PY��!e���|��CN��:%HE]����!Lt���L ���n����n!����$�0�����{-�x��Q�����i�i���z�U(3|���F�8wC���Į���g��s�����n�f*7p���qK���sz�l��cI��M8�����Qj��Q�*�x��o���]3�We�6�:���h�)if�X�5	��GO�0�v ���0Vxf义���=]zM�'4V3<���K��a莿�[2�T��6�n��N��H��|Xg�>�<K%ȯ���9v�����	aӳ�R��EX�&���W�+����y&�f���_Ji��ko�t�,��'~�<��K���s������-MD	��W�1��)�����5/��XD����<�����g�pesI0Ff��k�0@C�����,H'52A�*��HCt�(��VPM�zL��H˦̨��&��Y%5���\o��H�F����By�����7� �	�ϻ����h�a�#{{�]�.�S���������n�|�p����8J�&��	S+���?��rO�$��Ad���'均�q4("�/�e�U���>W+tڔ�K�����fJU̺��x�4��zݤ�5��\�<Eӆ+��������HO��/�����z6bs�G��;�\7=��o�`nd���zpf�vEu���S\��!�;-��ޕ�u���=0���6�Z1&���j����OB>�u*��g����������@R#`0�ӛ�s�r�_����_��뫈L����x���w�=�و�~^���Y��τ�E�l�C�h��9���a
T $"5�4]<���bo��qȵf�N���]Გ��D5�b�,��ت�lc��-%��Q�啛pAў�/	#���.Wï�OɼM���A��I�L+��˦������򓯶�H�l�`Eg��]��U9�EQ��h��w(3�����B0-�Sʸ'{!hL�-��0X���B��
cY�!��$��ȗe��R���VF���_i�R����d�'��:��8/���	z n�5j�=_Nz�u	��a�h���<R��������-���@�<��FrH�`EX�^��z�O�E*o��;S,|NS\S�Ñ�C����'��sD���L��p�� ������.L�����,���)cq��ȹp��}����ϥu��;)���A�
"F��M]��'Z.�*���V�E�������N��X��қ�V2"���]�-�!U#��9�jx��'>c20=-�r2?�� ��! *5��J=��'�4��{l�j�G`f�+��(���[U���m]��+.����s xݙS^ԥ������0������?�lfV�,N�{h�	���*��#F����<y\F�H������=�?L.�PeY(�f�b^�C�#i	z�tUvk��W�˻��^�բ���1�U:�L��a4n���1L���i�S��l����I���ֳ�5�b��?�mmh� .�ƶ�V���$�F ��5&�m�.�x�Y��k*g]���c�����e� O_ݦ�M7~�B���7��>Q�U��ܻj)%B��������z7� 3'�7\a��w|���`ov���q�i[f�4� �M��u��ã0��`9�|s���۵�$Y�CSငt��x/6��
�!:�&Rq��;G��ж�i���t7Ӊ)�n��+��'1稷��T�_���Cw�� ��(��h��J�̗�j��:?3�i�����r !�B� �A��΀�·�a��s�W�!�u\Ճ�N���� ��~����B���F���7��V���/���|�(����=�����ю�F���J�I=�٨���k�-"��^�&�o,浰���|6��Ԭ�mu7� �������YM))����.���P}�<�
^������zY�s�s��u-��J#��,i9q
����kZB@��L�%���{
?����G;G��rL
���[��\M	=#C> �qƘ�ٖ��FT��D���|�УF��{9Wa���o�r�f�dR��Ο�Sw�Ut����ēzdJ2�b����YCtpŞ��<ryI;qяQ�T�'t�f��M���y/����I,+�o-oq����e<O��1lER�/_��5|�3�E]�LV*�+{Z�j��� ��<�>��#ߟ��Q��0{M�^�ʡ,�u�T��J
�z�0�)a7��Ǒ��$��Cu-��~	U:�{%�1�I��ո��ϔNk\1�l��m/|
�79���)��D���^�9ZdV/tE#oA�C��r���<׮�o2y��Z?�~�\=��bK[g&�����1ytI�k�Z/�xpX)O���C�*.S���J�}|tT�P����|��͔�U8��#2��Q8F�i�6��c�_�,nɏN��� OO
B���e����!~u�JOC����LЗ�oA�M�i��X3��DsD�����wV����>���}I`	V��ba�7d=�nY��KG�b")������fɮ�M*V��"� ������3`G����'��Ur��؁z^G�GΝ0a`�iٕ��a���`�A�/���IuM�ո~E�w]��Ñ��i|fu�0:�G ���{��1H
�:}&�$���������h��.\f��X ���\��7Ё�N&��y5��;�PE�l뚇�wd5�4�vNg?����V~K��/��������LU�(Pj*��L����K$�E����)�CP-871�~� qx�3�����*kLq���*��x+��Л����0��so�I0ɖ�^���J-��n�wh�.�DD��1SGJ��a���k����Y��@�����>����]g	�A���J�yVY�v�+���2�x��@�R*�����AM��k�8������=�a���nkǤ�d�����m�À"�5�HZjn�,t���@�BBf�\���L2RƋ�/���琌���jCZE��ީ��v�,t��J��S,J����N}`�ۣ�\�Q��\(�HF� k?Zlkr�8
Blڐto���qM띭J��,��wY�1ɯK�Э|_���8�2Ң!V��AGdl�����-a�-��D�l����-5�&4�<̓�c�<��bf"KݖYQ�#�|�.s��*��W&�+�@�4��9�c�%
D��{#�B/��|�T���<���m���aGg�EtT�!�M�)>T�]�R��"��Mx;Ιkw�P�ď�I�Rsv�3�@Q�X�I��j�(G��m�Aȟ�IZA�t��?k���E�����@�zt�2��Q �� ��I�jf��%�X w�@���	-�[�v��U��͘m���F?&���Z���}�����
	�p|O|�|s7e�~�ŷ�� f|n��V]$R�_
^M���Jz����s����{ӕgu�b��D��������K�>w�b���c��������|����e���ɡ�4('�D�g�l��M9)�y���*S����P�z�C"��|��aϫ2$!�hlN[(͜,�9�LsA�nI���|�r@?O��B���ұf�K�}�[�>�F��d�~��=�tH�I�������;�.~e7ԕH�[Q]'km�뭋�5����D��C��Uja�.�%�ñ�R�����'[(�:�t�S��|��}��"����B�=y]���B��a�a���M�Jn���l��fUe5�Y\\��!�i1���iձ�Y>�:JZ��-e����J٤F�D�����[{b��1�Cj�nw�zO#���*�:�ۻj����
������y�y5����"��F����U�$�B+J�B#�f�a$��?/��ɳ߫�E2�1s�֪å.�T�'�!�X��AN}����gd��u�:F���M�%c�ER�A]B��]����E�0cu���>�k�#��N�0d�hV��,���]�gY�o�Eh��W{�a
�Dq}wEM<�;�"��[�j��J΢g�ٮ�yA!�3���`��_E엛Z���O�QO���{��rd:5fIS.ę�B��}\W�@�LH�
R�t�6)��NJ�θp%W,��Ғ��g6�ꓚU�՟pr��۽��<�G�0��X��:���*����v>��
M�ɱ���^�3^*��D���ǰ��%�(ӯ��8��-Z�v.���Y%d�-��%Uo:u�NW�mX?L��-q}�!�F�	��k�ET���kDf&_o�� ��\�ڐ�D:����u�N7�I�e�{���%C�xXdl}P�/�TQ,�L���mO:�Gy>�KXQܷ{�%�..'c,�G��.�
�5-��O����j����ۂEO�!���}�E��&t,Ÿ�wH �01�����!;>��(C���I�m�`�j���쑓
����n9�o��Ѡ�������;nvf@��͏Ɯ�
���"1�����k\s�J��Y
���4����? թ�t18�~����[����1ԙϋ����i��_Ոc-���j�P�,v�V9&N��k�E�%E��χg�k��Vr�����h'<n�й.u:;�mыth'_E� m,L�[�KRf�H�."ɬ�Q|G�p�c�U��Iҩf��������dT؛��؉I�μOy�9e��?$F~��䖑�9���f՜�U�kYgCPj�	�P���A�ꄞ�
<�!�Z�T?�]�4*�W�A(��F5��Уf|e��w�jU��S
������,ʧ7ں��	�����E�q)��Fp�>MbG"M+�C@�ZY�-��
��6^![h�QV�%�Z�,�Hq�EJ8D�&�J-�8��h�gC�O��e;�L�LZCd�1)���_a%�ͮ�89c�J0><]�H^P��>j=z{eٻ�h+�BC���ݔ���!���ᱞ�� �Ӄ
�)0�5'_���Ta�[c��YE� ]=��c�G=o�/�E3ȤA�K�f7�
.�,��V�5Eж7�xg.)����d�@�rl��r�E%]o��G�N��6���w�w�J��""�k�k�j�5�2E�COW�m��}��i�U�ט'�2�R8���m�^9�l�N�^S��gN4�&:���v�IU@��.  �Ծt���i"��-��(шa\��~���Cl�I��x��V'^�=�c����_�ک@l̚M�Lf��=��L����eˎpE|eq��.��"}\_,��Ê|�{#��(�j����(�̍H�!Gz���2ϫ�)�/�G�a�e@���k�sQ��,��}�ņ����[o�KAh�ח�Ij��J��Nz85*䠻5�<R�k�� )�lbW���"��Ҝ�B��F�G�se����HՓ*�jI��%ȮC�������EǮ.��;�G�z��.I ߵ�'��\u���@�<
�x�יq7O�	@�F	T��wz03���0��%,B�����CXMݎ�m{�}�v��3b��Ϲl�K��t��Ѥs��o|���dI�q5��ΰy�>�]�+zW��t�>�m��(
�_�e��D�f��]ɼ�Ud�p��%��l�e�Q��|ڙ���H�v�Tr,��BkƮ���8! a��wYW����.é�-^)�C�M��*hp�6�i;�7��)B�ԉ�e0��B��=�1�`�R�FK��;]L 3i����O�l*t�������O����R�q������]��w�5���ӏ����5�i6}�>`���&�&?���q��Z9dV�~�t�:5U����M���o����=I���W�ݠa�*�t�\����W)�?�C��nx��W���?��^YE7���^�:�H{TE	?ɑ��?��v&�.��d�����}��ĚR��O�'>a����G��"<��#ū�����K�P��1�
��Φ-M�a]�,^R
|8(��T_�u�)^�C4Τ�*w�#����׸\F��2�� ��7k@�(�"�}�{�ךK	G]ÚI�?�a3��hKƷn����mW�<�J�?ď��,�h�:񌇬v�k[G���;rh�W/��D��L�UMȁ�&Β)J�V^r�}��zWphy�T��39{�8P,st$#�ur� �T�������o�\��Vl9_VgBE�L��ML�����	#)}���噬ø�����O�<vX�<C�(�׼\�6ﭓ$�a����r���	�,�.b��q�~�a�\&^
���_���ެ�7	�td<�P
AizX�Xʵ��u�"�g�%�]`3.�����1?�>�,B(�gܵ$�t�H���K�\�������5y-\��>��%a�l�m��M-�	X=GIK]�)����Wq�rP1�p�)N�]�/�AY5���d��L�c����;���*�jR_�kIȥ�������b����-�������<�ʵL��R�gC���@l�o^�Z�:���ܒ�z4�N/��<m4Ȣ&H��1�U������˅ܼ���,Cj��&�25߈�ʾ�Ŷ�����N zSH
�����܅a���-f�6l�h|o��c"o����H�0]gY���xA�Fa�wQ'�j�f��M�#��z�x^f�����E��A���Z��KG���e�64�����FP&8|S3���o'Y������/b&����(���4�'�Eղ��﷞v�z^V�K�o8X������WP7����d� apn�����^-u��,j7}��Ȁn$7�	��]�S����Z����/�W�O��G{B�Pj��(F?����^b�T�j�	��7K!�T�:T��ŭ2{���o�0�%7yB�����K�?�W�`�;B���Ÿ�f`G�G��Z ^b`��yң��⤿pj��tE-�1N#�PC)0v�����z��6�P����ԁ$�+t��`���A5T 
���v(Rf\��
���Q���wJz+V��U؎��v��׈�q�:��uqZ��	D�����\r��7����ԩ>0��NE5� �M)~�Ea�)�4���	�T̓@/����2%d���Em��2H�P��73X��~��{��45���3�o�	�57P��Lu�\��T���ح{GT���v�ԙI#��&��������:�{=��~�<�j�P����%��&:�it��DG��������dxRH��0\� )B��+�Ũ(��m�����SD�s����Fx���0���������(IXI+�0�v��e���I�t9o?��<��Ư�
�:E��ut�#ߐ��#
��r�*w1�M�a��Q�ᴈ@*�D�1�@V��� �˯>�����a�5�:�x�>�lo�U��ӛ|��4�v�rP�1��v�L�+>�����R�{�^�CE,�M$���/2iۜU�@�s!/�-�'b��;~����&D��H��R��J�٤�B's���˜�g�1� �|��*'��t���woD0W옻���-��b�8~`���@�����9XnK��#j��Z �8�PPZ�X��o4#����`�P���
��J��PO�mN`�e�5e����S�Y@��K�l�}?�\��G���h\��D�Z|٢�?���o[o9_��2���SPk��8Ҷ>���g����̪,����;_r��Yw79^�z����@��Y����l��郴C�y�a z��Q
b�X�(U�zO�<�;*?�%�����)�_)
�v.?V�ߣ!��)�ndNm[/G��g����Ci7�\l�:�1M�����H�O�dF&�Ϝ���hQ�
� PEE��������H3�ʎ(�	�Ck+xl�{	?G䚐��ܢ�]2�
�]��*)��(������@1|<�9�(����g����2=Ү�5M���`��J�ET�=�jM<ΰ��2��T�6�`�3�/ŕ΁�qp}KC�oxh�7�i��l8�?�&3c	�A�|E�FUE�DB=uEÉ/��/h��R*�2�`�?�B�M�t�kaa!�l����;�����$���Hθ��:5z]Wjg8#t�!�<֊�(�8��)h���+����m�p���a��Yx���S���WT�i�XŢq�O|M��C�'cݣ�W��<vǼ��M��ɷ;]����	a��Z٬�ry��^�.8�����8��_`-,q���I�Gͭ���O��� b�9�-SƄ�@�����B����溰͟��a[��E[��9��?�l��0H6��d��&�2Ƈ/Nȼ�0��b_:"U��pi�O�os����,�4����h��*ȅ	�=���l�:��aAl4ֻȒC��߁������#�%8��p����w���U�oH����Ck�z	����Y��>ҫT�v%�:��XY(�5M�B���r��xm"���Ua+���H���!�w@{(�+���u���X��TwmWL��������H���i�RgB��GM�\=3������ �t��>�#��)[EW�T�\�B'�H���|}m/���\0��B��վ%ȹ֩w|���)l�&���G��-1u��R�e���(�����Q7iCmh�'�ŲN�0O����emM�G��s�0f�g��@�a�O���MRof���+�J�o��JFh���m��ߊ���5'z)_����e}�/�����}E�8�|�I��(5@�%N��P ��P�,�ѫ��D������
��́���<�	�[��#u�,�:���-�LUˈc}�u�+|� �<A��jr@�ͬ�� �)����ǉ �����G��I�)|6]�J+TN>�7�k���\6�����X��vhyTH�����9%�Ѩ�>ϋ1�����@���!�;�c�2���V{.���ϽE���dϚ4j��Ѻ��Ï��df�:���c��+W/?6�	Ӣv�fE��*S�
T�8q���V7V�`�ԋ�c�T����z�X*��ד�W�>)/�E���Y���)`��@�{�=��lJ�3C�9��g݆�O�fg�WW�[��X�P�����K0RFc�);��K��˴>��`D��KI�	����.�u��g´>Zr�W�$�p��(�t�.C���
~�bp�Ѣ����L�P5���ݮd�gZq����U�����^ԁ?$�(A�ʒ�ʢ��,�^���%[ʄ�h��\N�� �W�$��0!���T�M�2�%�Ԍ����s�c�M)uΧ�Y�R
5GVlF�A�'����Ոv�_��Z���YcD����aSA��
�Ȱ��^���������oW�j����e��K&�`[�v�̓�ȭ�N`�'�SE��� S[2�t`nf}��'y,V!fg'2o������pv��iGO;��Y./L>%;I�U'��)O_ܒg��v����s͆�ƚ�4��+�m=�9�V[���Ȅ5Cdb�4��(�]UX����|�!Vc��J�O��ʃ#%����\~i�Do �H�oL��Ost�i��&�:0��a)\)XZoW�=	�:��+��f9��R�NjL2Ov��Y )~�X29z�k����4aL|Rc(�-�f�8J&O���Π$�A����$|�9xh�bvW�� ,�����K
�?ِ�.����k�G�F��ڨӜ�����c�������$Y��6�,{X��/z�7dbՋ0�X�m�LB��V�7EA��n\@O��_4�l�:z ;a \�(����s�-�D|:��;�ϰ�� Tu�7��'���UnNa�Պ,R�ˈ�'v%=�c�^tV��p�@�/�Z�o�s��uy���ѵ3���,�c��������ʒ�)f��f�K��|+;�uu����a`b�Q��.�r�n�s
�%�(�?��+Y��k�	ȭ�Y��E��+�L�?;�H����	�����j��K$#x�儵���_U��oWb�v�H>�g_ō�\�#��s�q�biǆd��x��"G�pgrV�-F��<Y���� ��yx�����3���k�L��,0p���.�i�T"!�*>x��(�a�[\���<�|�$��h�������0C�.O�$6K�m>I��N����������8!����(Q��Z�-�H������;�ˡ�>TN���p.����~�5�!ǓP�|�br'�~@��R=��9�9�'��斔N���Q�eo�N�����F,����kj]���$����U�9�#V1���E�37��2��`��Z�FFp,�)�,A*�D����Eu�L!�p��o��t� �A����,Z���}�����.l�SO�z֤���T�}q'D���Î@\����k}C����g��PC)�F�/�P��K+}O%I�Q�
��j_��D�S�����-��ᓠ@P�q������d��̓H��d�v���~���W܉�����SԔ�&{�y�lq�����yQB!P$2��!@�x�D3���=B��S1�S|�x�jY'�z�I�M���}t�e�h����p���=��w�F�N�cwpע������u�Y3.}$��i�7��$�0��ܣA�Ҭ�Z�����B4V1��[Zؽ�ƿWz=OҰ�eܨ~+�\�Y�G�#q>B~eR��eM"ԑ�������,U�|&{����X�q�[}���a�W�\���?m����Y�*��m�C����u'�>�7�Vmb��h�7.dF��Bm�K��i�
K]�R���U���X������<C��W7�G=������C���u�윻��&ڤK�vV�jخp��ݭ�6�S����sV.J"�����ui$N���@Z�r�+P�l0�Ƭ��6ۚ�?�fN�����P34L1�F/Z�Σ4{��<�)���gգ��qڦĬ� ����t�S�S��/c%�OpP�z=ٞMf�]�:��N�]_L4��p���K�uqc�d�Xɨ�f��,/~�'����tv��%�ܳ�d#7�Q]�v����j�^�n#9��咐��R��O_ ��Dv���\�%&^�TW@��"�p��5��EK�������I	Qa� 6r���-���d�=�S��:��:�����SdX��FкID�7�)�05 �-��/��(܀v��,*��'�Y����:��A���fB�- �)�s��'\�STM�����tB�:z��s��PB�����Ɇwi�{�%��`0��1���O
r��C�#\��U��2����
0�AhV��3�h��&!(�ML�0�Mn�(�y�͜��>�r�����K�6�6��k]Q/F�|�
���o1x�Μ�R�>���D�ހּ ��c�� Gi��!��4Z�L�mALN`ke�s�����Z�& ��H��laȩ�\�b*q/R�*��te��D�?�q'0��~ɥ�/ʭ��NC��2�1��p�t���+��u+�6��:�dXh�&XW�p�!D��g$�q�����J�'�xM*�ѫs��n�mr�w}��P�u���H�����IKZ�Q���ҟ8j�:�a1!$Ϡ�q��w�������J������yL�h���z��I�������V�B@���!�
�^	���'�b�b�([#�k��vF�U3����Lޙ���Ć}��>�p0y]y䌜)tT��`?]�����j�����9r"YȄ�q�f�u����������r>����>�����u!=V�bD��D�v;
��X�ZՅd���׬t���"f\���f(T_�2< ���b$�L��(@��H�����=���E"���J�<#�bj���yB�3h���#z�sBc���L�7�;���:�Pfw@�D�/ǜ������M\>p���I�ä4�P���p���u�=D.
&�8�,��ޭ�>'��R=xk��>$�|�p��	$���]����'Z����Há�)����Np]0��ع���nt�u��0�-��F��SӘ�"|�s�o[wQ���s�^G#f͡�!CONᣗ�%H��)�D� X���-�%pw�o��y��*�M�ߧP%0�=�$}ѳ����{�� ���]DF�gB���1�v���'�̟�>v#k1��
�3�0��(������ ���zⷨ�����> ��