��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P��v�"<ߞ��&'��k%P碶�R�ӣ�sĞ������FY&c�W��f
d�i��vo�� +���	Eeҙ�k/�}�Ms�e(!�V����v{6Y�����,����/|0����f��w�����R�殙=�Dqk��뼱��aI�x���T�k(����E���b'#�.��-���1��rr��h�o�߉l`�'�u��8{iL������?���z� y�9�C�J�J���Q%�k;/��9�~}�QC�b�d��p�z."�������<׈
5�h�O�kgo�G�ԟME����q+�Н�Tmh�����^ ��:�+�ii�|l�ի��[���R�DW�=4e�7����}�.T�B4��+M:*CN��R�Q�P����ɜ6�<�.�+����}�?�iԤ��<��5UE��?8��*c{Z�Rd� F�-���q��R�������,��VP~(���{4FC��X�|�e�5�nz��3���J��b_ ����"�|���3z�'[��=X�gU�W�:��ΣpіJg\ΫB!�u4����JD�'�"~�D?�X-PF"�u\��ָ��a��L���Qwf���߰�u�0��}KER�&�Oi<^j�	��ٜ�����81�̈�k3^�1u��>kI��3��'�����5��%j�ZˑI��2R,O|O�8s>挲M�;�cc�E�I��W(�m"0�"�L�2z��Nj9��L�<��g��~u�AX�8ht���m���Qu�~qk�(FBg|/���3v�y�(\ϒ�M��c�����{7F��QsuTD���a:S���I%�����\㙅��.�'��}�CgS����/��Ƌq�n�x�:�����V,b{Y�es�-�)���!\�g�\��x�o��D#52��5pE�([JŌ�̈́�nĳ��i�tD���RS�ݮV$T�i!~�چl�[u*�ߴk�.F��aTRj��s��c��4_��`Z#�;y>]2�g5y[�������]g�y�'��K�%�=r�?B>	h8<������o9�̌{������3E�
��Vi5�����\:tO������m[i{_����j����-E�^!j��B���8,K&&��4��Å�q0��_lq�
��_�'��k��*��C7���[���|]�f�I֤�?4����5�|�l1:�C��YG�;�yC��2�h��=N{.]9� u?�����c���,����X�mIƬ�T�M�NG��`�c� ���Rm`��w��	_�?Ps��0R'l�A�|7��\\/��eCbϊ���%{�ٽ�r'�ʿ����N�OÅ����W�Iz�E�`l�IF������R^�VF��R�$����cX&m�H�vK �TВ���Cڄߍn���wғM��*V�:q��D���X� !#,��	�B���`9g�G7o��۽��W�Ok�Z}]Zӌ.�V��EWFW-!�s�.��	�?��i!D�.�=��ND��Ŏ���bnS�/	,ې[�H����08;dG�#v͜�~t3��H�1���PgF5B��}��(�r����W�O��
|���4���^&��1�q�̴4O�o���������X8x@!�ՇBE��*YϣI�Xs�
����|趝=��P��?�����v% Z����v
�s����c:{8)x��x��}
����f�5�Ma{|�%9�,T��k��pj����^��5�'��WayO��a�آ07طF�<x�]�$�1`f|O��E��Na;X.�;�_a�²m��ew�S��r�g���`ÛS&^�R�i���dW���C2��Τ�F�lG��='���:�����}�fNc�)q�W������lx�Ŀw(yWD��Y�v��!C�D����6q�Mc���pA�5>s77m,	clD��:?�`ʣ�DA���u�V��[��N�t�u�
eJL���prh@��Nj~@�������[�&�XA�NPxB6�#�i��E@���5�0j�rͤF��"��CC���6nM�k9��"
�o�r���;g��-�`��';qe�e�#����s5�7L�
["�[�DMD;`��tV<��N�`-Z޿�����]����ᄨh]��7]©��w�B�����j|��k��\��5B�]��%�Md����	j\?�p��dD���R6"Cy�M�� ��j[�8���lS-��E|�h���X.k�����G�>ǀ�	�����Y�:���?2�W�n.jϥF�X��> *�0u4�b"E_�^\��4�a��6)�{�'����a���r�Y0�Z����z�� �ׂB��4��8�՛g����m`�e`�5�P�c~��)`Ŷ�%w�Ω������Q8�v� O7�u����D]x5j���(�eĕV�*�;|6o�	�Dmǈ$=��$&����T�((�MC�+�w��)�M��X�eD)���'ƹEˌ����<�2W�c�"l��D��,�ŨpW��im3�ؒI0�B|��Fu׾F�$�Ar�;se�Zv��c�#���Oշ[�V�0��E�#�^������հŎ��ZX��}���+W��$`)�v��ǚ�'4�L���G��y������Ǔ
���qϭ3vqx��(� R�~���*g�d�~�9H���,/�7�}��2U��n�+�j����+G#��8�L2g�R?Vw���m{�j���h��$&urE�
��g��~:���D*�9�vh��ɷv�0	�mĶ=VP/��w�#�[�a��r�0S�GRb�Z�'���m�V�V���>����gF��@��Hx�}բ��g�J�k�2���Ǯf���� TG�_o�i�����"�8kߞ�m	!�-�q���*�Jp8:k�IQUP���V��h�P�Ӄ�AX��r̓� ]�G�}��^ԍ��hvP.���1�4c`1�)
(��Hh���L�w	�����|;�H��y����y�"�n&[3���y}(7�c��'�DÇE#�|K��9E�0o���h�p���QJ��z����R�1�K�%_�ft�b�?�U���D��֌�2��)���Ǽ�B��鍆$��A	mc�@շ]���|-�u�w�%�k� ���C��&�h��%�0��@AXK7R�+Fj��ZVY�?���j^ �]k]�n1���m��U��F���>��@��g��h�q���o�JU�·�`ll��a�Q��(/�V�ϼ�.�X���(�'��ē��ģH�M�"q���2I����F<�iCqE�'z���������Ч�X�`2� �'uQ��Ο�.g� )��w��4q�iZr���w�uS�]c�^ZV�o�{#5����I/˵�x��0Q����|��=�mJ5ftȽ����6OR���;��O�KMK���&���A��N�1���Uݤg�4g��*���C�EW��Ħܳ�������S�j*ؑ��A|�#�$���7�{j��&�]Ж� 9�scW����-�|'�3&�	�ͫ����s#r��pXr��e?_��P��	l"��Mnvs�1?|�kf#	�Mz��R}�͑t|k��2���J�����)���9ْ.�[��:o�S��ʋ1���65ݙ}5�`m�]�-���A�i��O�y��9�`X��;�9n����O�(�`0fd=@�&��P�Q4�Va���0�������`8�Q�;d�}���܌�f��C�i�:�I�b��,���+�W�&j3�|��[\�7�@��h��E��K� �vD�G�}4��?_B�?� [� �4|���k�g˖��R'����	�;���(c�O�J_|�=�M�N(H�U�C8(aX4���4o����^<-M��#Q��|l �x�2�Kz짘$�_O���in�>�b<?�y�mSG}��?r�s?��*���4I@�Yն�U
��KkWsT9�q�����@!��1İ八�\ g��������xg��؋�h�>��l����8�%�g�:����9|�-��c�𛄺�{G�f�R�H��u�8�<R�������M�Y5���$0R�ԣdr���]�_<�է�7ơ�١3^��o��ȡ�����ԟ��{_[��+A�5���DL�����X!}b_SX#�'A{-��kpP�MN�BB��K�bӎ2:K����p�I�p=as�L��i�.z�9�O*A.��1�nb��K����eþ�+�<d��b�T�\*u����E��`W����P��簓,��UGޒ�G3�����j���޴$ޡ�<`4��xe��~Rg|������y#�5Z4@��L $�8�Zk�tۖ��[�YUb�5�@���F ���������5�\�ElL%�Lx>����_؍�~�wa����:k'(��Ķ�O�旊L2���p~0��j�c���d�^ޗ��'��������&���/�(� щD��ݞ��"�$�C�5Xa&8����nY�*��s�����b�а�?�m�KY��T�N�Iә=��c`Fv�#e���G��͊s.�x�1������G��(A�&(��],G��k���A�Z��s.Pz�&�����]��W	@ִR;;��D�(�����sur��L�p	�q�9c��h��s�;�b�vU��K{�m����;V�
�rOI()T#sPg�`���v�:�� ��8�ŝ�${z��ǵ3W�-;���rhK�Q��G\���Ѹٴ5�l�g���󌻫q?�t���)�޵�I�Yb����X#;�E�m��*�3+��`Y�}�0�a�_	��Ƭ���W���۷�]�Fn�������QR�`���6$)����N��I a��=��+9�������=���2B-�e�j`� oW�e~2xGK��]��$�	�\�]��]���%��P¢���o�+@�oZ�g�2/��^�|Af��7��K�oU7u�jN��B���a��Ѵ=�����8Wq�y��0�	Q��o�=+�r�ҥig�̖��(0f%�U�m���,��B2��ҚY9g���g�!�t�W�V�+_��1����b+�F0���/9�6_���B��L��LT��a������MEw�9[����f��O!�> ��C���Z���6y��DT+ �� z^G\C"��Q��<j�������*"u������Y ���,1
[��tI��<��-�)��Ǵ��]i��JT�{Du��zey��&Y��N�ǑsLz��R�e�Tz���vb�k��d˛���Z�==T�0�9^h�F!��:��T�H�T:���EU��"�M`J������Ǉ���px�KШ\r�K�FE5u
�b��D}J�����G��/��T[�YiGr���x�3�K��cNl�,ϋ�t�*فѬ�p=���xH�Ge���1r��50���k1V��vBF�1�b�ݺ�G?A���ìŪU]s�u�59��s����q�A��.@�4p1��1���]��h�P��(�{h�Kx*X�;��C�9��q~��{����r�SZX�m����60]�y��W �O%'fl�YJ
�˾��/Z����n:���Yx����,�Z��L�<A��ކ�[|���n)�6��^�cQ�f��c+n����{
 g="���a��<bW�g�`��g�n.���C�2""���ݮr��
��!	S�u{�Ȭ��R��"<����������������?P48 ��\�*zR�t�+��7� �$�n��#_˜���h�(�L�$�*%�S8���;��={��>��bP�B6��c:B�(����3n�Mu���y��K'Qvc΀�n�#	�dM&Xv@�E|�F��ֶ���QiD�o�-\�k����u>;�|j�>�w&u�I���U�֏���gS'����+��{��9W��ʋX��&R���TV�%��
���yno[ض_ȥ��@�-�rٟ�Q��p�_˶��%:an�z�vj�H(u�$bAq�EV�QK��%@F�e�����د����3�l�T $Z�n��XK�ɴ��f}��'+b��NV����G������Eއ"0��j\Ľg�@%{�&�ż�;����G��s��٥&t���<B��3�M	�����Gh�	<�������vf܂]ʟn��*�L�#_6�L��t \��y]-����EVsT�]$�W��p~P|z��]pO�Z�α��G�R�`Rn�uf���g����W��r�ҙHz&Ǡ,~��4F*%%�R���Õ�n;aO�?hL��\�H�s�7g>	$u�i��)�������,랐��٢k[XN3 #(q7q�xy����(Xԗ1=9��"�X�.����LI�V�M$.�g����.��c��9	�j=W��Yɴ~����y�L.o"T�ʫ:�}a�hs'���i�
L���F^x%��Qkf���C�A���ŨӘ�+��	���ELV>�S���֙J,n�8�X�t�p3i��B�)f#����=>Sl�'P��K���������J� ��G��Dj������ȸ������D�	Z*�mA� /�Hf��yt�"��e�!*�JX��SI���q�>$�o�<���LǼ� C�1��
�#1�u~p*D�afU⋓��?��S�o��m7rc���+U�Jgh�>\���"��0�#�g=jގR�"0��� ;,�@��Brwu��5?���i��0�<��a��E�\��x5u�P�ш�C��S_rC��#��x�|=Aߝy�sN<L��5�./4X�;�R��s�2�G-��/�i�5x4C����)hR�����^	�%�w����{ࢮqy?R�_���1M+� J2��~/�1lQCs(;k�j�T�{��yk� F���.>�k_G��I��`��,]��.�"*i��y�8B����
f.����)�g��~m^��3��*��Q#���k��;�Տ�Ng-h�S����U=���$�NiE�ykf��O[uȎO��N�Nkq�k�n��xv>{? ����h�e��C��$�R�L�>AfG�@>.&�k�'�C�����aj�YGE3��p���Q*�&��ܡ���Vw�1��N˳�Ȩ6���r�'�v!>]�p�1�=b���>iQ�
5Į�G�P�tV] 2��|欄�P�f{��AX1�Fw_��8d&�EEKL*�p��l�3����͒1ch�91����;����a�H�h����J݃5y�u�yj(5�v�j��K��[`�7(/Gv_UT��L���R��X���j/�{�9jΆ9n�ZZ�+�[K������M<��p�҇&��y��ϟ����?M����27e)�:ć��.\";꒎e�j��er��0X�x2��"�5��Z��7�T�E5	��VlS���!� ,*@�@ܳ����{-I4k��Sl��f񛑃.<�K~��h��+����2�h�5DW��j�߇���eL�*��:^Y֡$�0��Pt��=?~���s{z����8�!��9�쎰��"H��0�Ve��%�&�v;�F5����*_�0�&��u�SZ��7�/�:Q&��X��y�ڰu˔�u�(�2`Z���T��x�?r:d
�pc���g3R����>�Q��}���5żJ��oJ}j/в� �>�L�k�X)2�9��D�����neltM؊�$���W�#��{%�\� �;���
����ZUQ�ȴ�S�!ٹ�XEqՔ��'��lɞs�"Zb�(������a�:����&��9s-Y��2dx��qv9�7\���]�W]��;aí�$�T�!�Q����b�OǺca��Ob��)WNVm).�*��!�����)Y F�`������A���۵�nIP�w.-��9���6 M�(�q�;̼�\�������S��'��֛��D ��C��ub�n��:à�k�C�"�6Q"H�AKe��Y�¦�y^N��ġa���
���_�W��w-�=0<Jzݨ5-�����a�������B/��c}�����犖l��X���	�Y�V��O� 6p��L3��9B�Nx�}���\^���>a�wB��7�͍O��?��:K��Us2 �v츩?��D�_X~m���~Q=on�.�� ڲ���E:��ƚR�fO_<f{��S����nn�f2 xm�gDק��~�5>ӻ]�"=��tC�w��"�Ƚ��/�wƥ��¨0�D��2G=ܸ�o*��l�Si$�,����/PE�������<�(B�d�x#2�f�ý�+��Z�0���V�\=��w^�&<�? O�x�5;}�5n�l_*���.f��M+s��@��\
+"}"��N�M�ir��]�2=̏C�]��^x��$��6�{}}�9��1ؓ7��N�f!���6��>"�]18;�������%�A�F�F��pt�e�'8�*	�H�^I� ��\~W�E5~ ��AuG������fy{-�N�1�QXG��l�����^�^����Z9K��r5�:5M+��5'�C�����dB�ח�z��, `��<d��W��ԭ2ʞ4N>۰c;v�"���e��#��s��S��$�z�%}N$��:�o��t�$+<�㼦$�MW���żv@� x%�1�&�E׶�Y�*�~F��� �>�즨,R���9�R���3�)���r�g/�r_״���M�<�^�y�~���%��ڵX��d�n��R�'�r7���|�\�SU��9 ��Y�K�����5x�4��̶}�yo�'jO��B}/A��d۫��<���a���@9��ʂ'{I������dî�Pi1 ��<a�