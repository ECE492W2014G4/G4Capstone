��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>��`HX����5a8Sjf\�|Vv �|�
���ۇ��������)��T�'�L�3*�51?+"�W������7���׷� Y�[�}nP=�PyW'���J14��qKxW�୽�V����+)Ό���-�o(��Q��`�`߱��H=%]�ȗj�u)9P��?L\�Y��rq�+W�||ꅡ]����Ҿ�G��=����`��	�*d��y��z����'ݤ�ֿ|�TI�7x\���B���挪}wNlR�p����\S�l����&Fǁ�`>���Z��K��EN
���4�ȸ��2�^������o��$[�5J2��.~��\N��r�8 3k�~E�F�%���p���:��:H�%9�χ�H��SHg�7Д[v룕�Ɉ�x��Z�S�9ͭ3u�.d/�0W�͛�B��U	�Tq0&Lxs�aQ|�yk��8z~d]j�V�}�~����@i��Y���"��t?��yz�ذ_b7)��Ar
���Bu\�J�9k?cY2* |��Jw����0s ��\�l��|IR
K��w���V6����H�Z�!���r����&.n��Z.�����L���d9Lmq\��%3_�E�ڜg�b��u�l���ez��"�4�O;�E���*]hҞ�b#)��9G)�H!rX�(���e�+
w)~"c-��
F��ݣ@aߥm7=`���S���/mŔ�21���%=�vL���e�T'T�8���j�p*PA��z��iob���o������C`��� ARR{�_���x�%�S��u/A�G8�Vf���T�Y2�����7�f'_>����E&��G�x��׍:��q�S�%b[�ٱI�W(y� �m>|��%3��E�t�|D������ל�r�C`~ʶ����dd���"~��){[[����T�to�Q�
�Ó!�U�x_��M�z�!����1s;)��<S.�(�T�ѯZO�*�������7F��.��x ��* eʿ$H�#3Y��	��J��k���N�\TZ+v(�U�);��{��<mg˖v���}"��F|Y�V����G���u"R�ԉ��g�Av�
$n�C0H�c[p,ٗ|�����e��?쓪jG�p+p�rif���>�Yd
�)���m�#���07fj�E+�'����,.X�l�� }����5ᆪ�{M�[4?d�	�S��"vW8ƿ��Oz�?N5��±4���?���?���$�N���B$�	��Wu��+X�8eK*�>>,�ū�i�q�ȗ��(��i8[-C�J�S�y�c�z5s���QA/�E�c��I� �O�d��0��/"� �c�+��8Z�����Z"
(�����q ����/E7;�@iY�X�^,��N[ �?����R[ذ�!���03����S.�nq��D���S��a��]9��e#F�%�����p�'i�$�e�L�Ũ_�"0C�H����-xX1�!��6C�x?^��6@A-~X�Ŵ@�	Q
���+uq4�J����pj*�B���l>T��TC<�OBI"On�st^����7��Zy�bBmM;7�	����5��Ǌ|HΖ��~IDEss�ML�~��c@����ҍ��+�)�M�]X����T4j�O�3�-+��B�F@>��r�lE��:V:yE���4���96�������Q����y�|��e��#x����b����-�?oa��߭f[�� 7)��iX��V�7�rBN��Bb�阣�i
|C�c2х��<��^Ͳ	���.H��we�	3� �����n�p<'��� �"!��Z����"N)��oD�lPU�ѥ�s����R � {�b��I*��͎�����CdIהh��M?������[����i�p�'��?ދ2*_�ߡ5�����`�I[�^�eɼ���4~�!̿��+��@��ץ�z��I��A��4�`��� �R긷:d��Q#�}e?� o;�^`$/@2YJ�5��;Cz����Y%6��V���Ou}���i��]"�(��SB��.�Ė���H�"({��Hb�u��c�Q^hPWm�(�jd1���ыٛ�A<X�,��!����{�J�szD�)wV������mo ���N[Q�[C�����v _��JA��L��Y�-,�$�[�2a����NT�7����_��ð�����=k����pN%u����W�x�$Tn�涥vUg6%�/���Z6��c����l�Z�C�ֽ��I� 0R�]���uSڂ�����%#-~�Yb(S���Y����՟�G�ѫg�'�O�����}������=���i�t�.�.nP�&V��=����bx¡ez	��&�FG�|K-��M�u|���(,��;�n�����`��޵9�LS�������a��9�J,5���	'p���o5��<)��4�\�d�mUuy��2�梢��=R8�vl�����p�w�9g�y��H�/����7�Be��B1��e�O�:/����Bl�RT/o�١8U���f��b>��G�-�j���5ƫ�^+�~�W���ϯ��=u����H�P���ָq�!�[��tuW���>����C�1~FICZ��Q��bx@4}A���R� I e����q�)%Èp�c� I���.D�}*@�|q���58��[:�3��>3lM�tjvZ�l��^2'Eg���QLm>x�)������&̅�l	0��b�e�y����)�ŸhΞce��Z���龔��P��L���A�.0�0�V���&`����X/�h ��>;�F�M�wT�Z�W�?��/O�k�ʙV����n�c�e�����Wޮ��o��IU5��%��40[��gՊѽڴ^�q�\��i�-���62��36J��>T�عV`T���X����7:Q��u�H��Ӂ|��2N���:+?Q�J��ܽ�����B�ӌ�Q����������#Z�P�e�K#�~N0��Th�Ť������ݏ�C���X
���9w���>dsAÒV{&�����X���L1���j0!�?G;��]��q2C]5̣��k�{#��NYf��Z=����{�AA��mT,�e/�����SaV1�NP��ɵ+���,���:3��J�a�О�^����?���TO��>`ϕT�Xu�����	��4�V:5�<�x%�$j���h������(v<�&��)V�����N5�F6K�>�M��3c0��	:��é���Y��9 �2g���T�j��8�� s�[�Ҷ�q�uh��x����)��l�hO0� ��� w]Z�O�=�qے����?��5��-�4kB��#ֈ��-'�ۼ\��K���m���u̐Lt�����S@�M�	aN�e���y~d����b��\j��|C������{�2ZK��!~�+�3b"�D����l��#������7��%����J��X���#ϣ>^k��?��<���/�/�@R�0��'c�.�`�j]��ւ2�p}�)�~�u��Z�2��p0�f��������32����m�~;�.4�������C��9��j�[=���9W)r��l�����KGbp�]�/U��x'c#] X5�1���TљE>�D�Қ�g�����)3��}�����Y@�E&B-��п��E>o�q`P�l/܆s?%XJɅ.����J.6�|E&S �u�b\��p�i��3/���8&y��� ��h�,�{��+�a������a\I2
x�&k���{h�gP�5i[+�y[�����@��C��o���C^��ٿ;Y�}���m��'a���!�]�֗����z�Anq,����u`U0q���-�_nsgb^�>�M�����:��S���-=�D��`����I�{�FфC<�Ƅ)|u�rz�p���#(���1ۋ�e��<��x��C�fh]^ޘ�"����Aa�$u�1���.���0�2�4r�;����եAD����Z4��R�LK����(XL�z����d�x�~븚U�	sj=��#3��/~��Tp�wBoO��ŵOA\����;�I^��W ],�Z�6?<T	w��ۯ�[R�����г�~"}o�����/ݔ�j]ѣ�)N�aDN��g	8Of���x�Q�׾J��o��$�C�T�>M�A��t{�  f���H_	�M��햧޲��F���V�d�<[v}�Q}j���4(õ�\��aǃ�$<&��/��W��|j���@yը�'aO�$�uS}�͝(AVS=!V_�
yx-(�]��$�k����B����]偄#�J3!���]L�;�ʩ�=.?�-�fJX��Tms]���/ ���W@�ި�v�V�4���_L(�\�t3�y}7��Ww���*�P�n�da��7B�Z��E��+�2G�w��Jo�߲o���'����ٗ��rq���l��02����i�m�c�)���&��tN��� ��UT�|����f=hS
"!+��ۆt[� � (����z�J�[Ni��j�s#r޼��9��D�������&��f���B7�IyI��s�^���[�EL+����	�^��?�E>��l����٨2ء �4C��	�_�<dr#��d�M��1���D8T�����U�ud���.EkKd�)-�b_�d���(W�r�@��g<c<�t~�)
��G����Hv������̩gk)�s�g�ը.D���<X}Ч���: �wUxb��IIO�����% fR3�����#���K;�NՉ|8z�[JCHU�h��B��0+�{�֜+D.���6DUě1]�a�ࢮQ��3M�� �~��_��KB�7�?�)oT!(���<�k �����-S5*\+&V��qh�U��6/��qNx�<p�0�Z�7�M+�[����V^�7��p�YG������h�v�TU������Y�ONp���l�$�F��emY!7.;';+T������^
/$�
hd�������C�2�L~tX�{k&%�����Y���5qZAd�����-�H5SN>���{J�)����h~��>��	��� �j���Ĝ?�����	�Aم��{J�Hz��Y��x̡��-��SV�qTRg	���nr��4��<���r|�;�7�����,̤���p��˽
&�'s��Md�_��b��9��u�����j���QF=��u~�{�`��/�_P�}F]�w�Y�$�Bo?
>�ϕF]\�A�U���u3p_��>�,�9lo��	�p����3s�)ya1��������j�e3�9���aW��XC��I'�b0�qU!�L�+:����?:�l%��;�Ǜ��ƾ�~�I �[��uٿL�; ��ɩ��,�K8K��,�"9�N��x7g�v�-vf"��=aSD��T�����|d�)�J���a���3>�;PJ�&B�*d�8o�D�S��;�� t�\�@DA���x�R�m<�f��$�
�R�5F8H⦪Q(�e�����$1'Q���<�s��O�nR�T�XO
W��A�T���R���G�k�6zY�*�\i~�����.��1�S��VT@T�f&�8��:���4����z�Ē����d*R8a2dGç�6*�HU��$Tch˓�\�6Qj`Q9q��0��񺊑{�s��:F��e	�i�B��&}��+ %�(�$rm
��20� 	h��Q
�.6�ǲ�B����Z��2"��F�uH��<��]�8σ����`�K51���'����ޜ�F��(�4[���]�U�֡*���tU�mU�󎕢ZQv�����Z�0�6���*��]oͭ�h����e�#}��Q���Z�ue������(�5��FWW^������r����@*�hN�Szl~~s��B�d�G'+�0����\�Ե��`�C�V!!*ͻ��o8�;%Й��n�Y��ʿ�Mb=�15���[���nP߫%�Ҏfϻ�~�^�ۥE�r0�\�����dҺ/����v<���ob�E�>���f�[���ǎ��zwk�W��U�6��P�>4:�	Ѹ����2ǰ���,�J�����t���Gy*��o-G��DUh�AL��c�.~p���T�t�f�^4�G���I:0���rQW�P�W_����9-�O����Yk5;~�ϧ��5stj7��Q�(+�X �sIv��l���V3� r�$�g8����߮@���eRG�`�1��x��?6 �xȵmا��"E�$֏�?�u@v������n�z_�z�S�{�}I���9Z�	A�����_$@�7=�DZ���zV*��=���{K�&�J#�����0p��U�d�W���b��F��D���\�0��(dn�3؂R��I��.�t��C*����n�K���,�M2�[Z"�k���T
m�R�d>^S\�D�C�?J��׫z���!'1���V�|1�&! Lp��R��1�_��]���K���H����k�3�M D��x��U7�s�X+�(��Fh$v4���� ���QIZ�\H���N����tg%0��Gx7�$��G�4�,sȄ�>)�!���4/v�[^�I}��莚-l���*I�ʠ ���=���g����Qmu�h����`����_���Ő��*�X0#X?Bo'��2��7rù5����uk<Zq
�q'�61�bt�;\MPXm��@s]�}�N�K"�Q�{�,9��4;�)�ݻ���`d�nv�qEK���Y6�(������MA_ST['g�����0˝����RQ8b�461�ɮ�"�0����*H*��lW�=�Ѽ�]U&�2��o[�my&�H,��ݞ�礍'g�3b>L��;�>(�^�o� J��E=su��������3�=X�5}�S�
�L�z����P�#[ڍ�������5@mQ�ਡ��(�B�& ��LK����L��آZ��u�ى_�@
�f�;��*	>i(�FT�W�?a,�ܴ5��t_K�hO�(�K�͎�d|�6�#���ۆc�4mь�|C�[`n����|ꁧVG�ղh�'i����Ӛf����4yUh�=)psj�ǔ�T����n@̥@,ܰI���{�-�	+kݙf0[q�BՄ܋D���h��,��[������.��M��7��v%���*�)�R���T�l�hG�hb���}Z���W:����g�3��7]�d��荼P'��LX��V�&���&Ĩ�<��Ԅ]\�:h��HT�{�.�<��� ��R����Х�]�\�d(�)�?�%ӐG�Bׇ.	B��6�X��P���]�����ˡ^�Mq�qE,�߇�:PW�e3o͗�c��˰P[�e��C#�*�4�i!lrf�O~�GU�ݮ�K�.�pDtj��n~N0�]��q��v�}ǽ:=;c}�O>b۷��HD�u�N%(�yvc��[��l&����%�A5ϜJK������
p��(^[.�����=�$7*|��Ve��_Vͨ��s3X�5S[!�_]��"Z�Cpt#>@�cV�ȡ$��gP�^���͐���C�HygD�'���Z/ �4�0�Mk5R�uh��4#���cӪ`d�����{+��O!���iݮ��m2zU}��}D�`�F��g6��k��k��j؜��I)ϋZ�E\u�y�(�j�� <Qr����^�r�PhFԵqj�hY��=ט�%����n�E��AL"�B��qYgգbH�4����	b��h��yv���h;�U�Xj�F��R�.��Mx����M���2�K�f'oi�@��N�=��q���6�����s�ibt�$F2C��{�4a�A����m]P5��u��έx��ߍHȫZ�S5�X�,�J���,?�/=y)�ֽ)�x�a�ۣS��Eֳ$�F��g�C�Nh�;YeZ4�]J�vQ��8ֽ���VNvv�8�z����NdB��gkG3��%�ZnC��n��!q2ʳ^5w�	��a
c{t���o�߿v#	��7��H}l���Vp6�/���� ��$�d���5�PIds��U�S���l�ذ%e?��k��mG)���Q���'��N��.SĐ�j�z0r�\ǳ�Z��T���������!���-�K��SH���+� �4'��< ����F�9��]ćծ���~._�VA��"z��z툺0���$�wKj�:ccC�5՘72.��UJ���.2�������?a���˲?�DFW��h|�Kn�$|����ݙ�_�H�t�a�A=��*���]5���Ŋr@��=�M)�T�AT�vnj�v�]I�%J-��T��W�~U 4�̓$��,.|�P�=�#�M�u';ˤ@���j�p�$��}!�L�vAz_��'���J#�K��g��;m��8gU�С��J���X&Y@	�]�A�%jc辪p5�th�ՍayBw�.�1�U�.wx�:��A%|ǅ�Մ�tٱ�>��%���*q�?�n#t6�՜d���P��މk�#D�Y��
��F" �'�����p��aFnyq�x�G�&3W`~�ډ�n�p!���WjJ�d~��A��|T�|_�K%d�'�n}�0#tW�Y�jx�۸�1m��A��9�����p$���3g�?}�ӹ�-^V��{_�d(���0�����vRUZu1sH>�D�kSǆ��؋�RaG�E$������4��ƯME��bǶ2|Z�\���^aq�H��4=�_�ϣ�5L�q8������	#�ҡ3����"�od�<�͹�S��Æ�]D����%�G�s���a4��t˂m��ü�*�%rT=H�� �b�2�,n.�p���g괯�z8Gk5���~�R��/��*4�@����������G�� �,�P��T�i�^�ێ�P,��E�'7s}84��%��J'��^�jj�f�
X+�<(-͒ F<����uK���,w0�.���H#D��WP]����Т��,���x�uo�� ȁ�:���\מ�x��'�|ʜZx���uh)�������9��4��3�'m��Y�Hva��w��8��Q)1�z����,}���3w5�s�d�������y��!p�?�u��w1%P@���m²o���ϵ������S�����hѫ�p�eun O=Y��_$��g�r��l�"����!�j0��`���%j_T�xT�M��q�.�N�� �"f��E�X�[��]���#����1@Z9�F�I7!�{�?��?s�n{N �~Pa�Yzv�ՆfU2���|�:u�:�&LԚ�?����Yd矧E��L����_�R����6��~r4�6����G���oƷ��X��t�=�烊��-������iiʥ��NM0���؋��Iؘ��w?�<�
������2;{��u�{b�Dn�V�6�W_5������~>�-5N?�����h��?ѭ��up�|B>���|Zd+8�2V>p"u�s�r3V�@� �`���;H!$_e�ڸ$������/����n����
�tW��}�|0Q���:�+��l�]>�*<m���e����C������4�M)A�̬p,�~�@�M�M��I�gc9���+�v@��=lXk�3����6����>G���&d���~NM8�.�5?�c��}9���o��%7�g�M~6��Eb���ӌ���1����6��+�#̎´��'�H� �Q >�|����D�f�i|��fQ�����n��t���m��%=X�#b(��`��S����X_X���W'��B�채��?���H|�P�ꠃ�#M�"c�x$K �vH㶜IC�xv�$�����U��e��fH������**NT�}�����83'��znG1�0��ޫ�����>�m
�P���1�E9�ޖ�#������@*���O������y�fc*'�3u��I���9�Y)Y�ܽT�;n�M���s5�{��&H!��6������H�����f��}#a�������Ӗ�r%��ê������?�7cz\�Ѯ#􋇞����9���� sY(�m�3Lʤ2��/������eFʜ><����N��&i�=%J�/���F;����h���V*�¼K| ��\rd%c��#����"Zڄ��Q;I5� ��2�f@�~�!حRI/�'����P���o�σ��n)����c��8��_V@���U�������9ȸ��<b΢�|޳#���m�kA��/�U8��	�fbE�^��#�>����ѫ�b�T�KF%�C���+vc�LVá�'�'sl�wGy��䁔������xSd���:���:�;�����E�Q��1�P^h�<^�/�w��Ha,��B�:�}'U��� 6��Bڐ�>�f__��+�W B<Z�YY��N�g�.��{7���Y뭇;"I��9OZ��JgYSq���yj^�W��mzl���9���^;H����&�q��g�W��y�?Q
�g�*�.&�q*Ɯ�����]l�T����#�%��o :�U���=�&i��4�Ĉ��ƪ@q3���'�Ռs'��t��) 	� 4��� ~��?�#[=%J�\UR�ȥJۣ��z ]]��>׻ێ�� �w��c��Dz�9\	�/�FC���f��@^��q�0�D�|��W�c6e�9�c�9<.C�}�T��2��:�3�nB�p���1~+�O'�Z����h(l3�0��9��Kj'����<K_m`���"Y���{Rx��Ӭ�M8zպ�m��wҠ0�3���6�{��(W�
�� :��E>�A�Oy�\�f���[�kj����:�_��D����Q�6'F��\�}m<�z�y�ױ	�3�	�lQ���nl��/D�g�
�`p؅b~�:��7���F��ض=ڟ��1��}�~���)H9 �I�X��su�!�k1,���S��5f#j�J�-��qMp�����_��KN�P�|)�������xe�W�8���z��[S���h~��S	6"�lvp��-!�*jڠ�+���#��v]���������IA=������;���TJn7m�S9+���+p���{^{ϣi+���5�|2'��$��Ķs�����V	�w$>��V4�X��8��u7x0Ռ���$P�����S�1פcEAn|H��a�C�)�����Ҩ�
*��<��}i��z��4��D�����f�@��h��$������R�6��,=�=����,�9G"������:jL��JT������w�����!g�ca�y��]|��˼� �t��hU�z�O�~��R'FO���֗V �aF8�X9�|�&ܭ;!�\��#��=X�Nq����z�a�v)�!�Fm!�<�{��4�I�k2�}��c�q���/J�Pҗm�4�H8;?�U�R?���O��pA��l��o����G~�h���[����m2!� B�Xw?��xV%~%/��ѯ�3>MO�R_����}�Pt���EV���3縛W=5�$f�C�i��}5�fij=��`����η�ьq��$]�)dA���1��m�ϼ5��������p��u��t����C߰�#��(Y2wj8�C�Wu�|[3��!�q6��vh�5���v����t��m���jm��
��M&Q���_-��K�_��S_83-�{�TP�a�ŇL���扒{���>�?I>��s�/1��|rP~�U�"+!ѫ�") "��c�nިP����.�
a�P5NLGJ�w�۹�4>��t&Vj���N��^1����#T�:�����b�V���Y�D|��Qx��҅���yE2�L����RH'�jrS���O��Z�A��Xa����zp8���Ͻ(�H���A���czh�Y��,�GE�eg��⼬��g�v��-�/���Za*�m�e�^gg�3{�9=gZr��xb$0���l�Ğ����r�M��&�ʤ�x4ޜ��惻E���R�z5�����ux�}�������~��XmoLU�.p��.B�5����ƪt������:�6�� �!�(����Q�:�����V��it"b��d8���G/������R���=ZȨDp���5I2hga�7s����/��In��=x��9^}/cP�<�6����1�t&n�X/m%vr�/;�7+Ln�b��t�r��M?��B�AF����[T/��5�J/���=i<��8<�i��4�
�jtO)�_H.Q'�p�i�s;F���6���Ñ?2le٬���vg���1�SXl� v&�W.��y�I�f~������PZ�J-����?Y=�Tڑ}���c/��Y5����e��y�s���X���d|\�33J��V�t���e~�F�9`u_�������V��8��Rع�����8��8�Ng��u�!Rf��8L]�
ު�E�e���NɅ�i��9�����!�������P�;<o�:�2�Y�b���ߊDtT�|>9��Չm�E\U���u�1��/�NX7E�A�S2L��Į��qa&Gzs��J;#����[��,N�LN,��2s��b��2h����?#�FRS=J�S���X���i���a^������ T7@j�M�Bę걟?U2�=j�#�\��bg�S�W�V 0��(�
��T[[Ք|���Q�Ij���)1_n��b����	G��Pg_s�w9�7��e}����H��b����^����t��v��䥍�d�}��ZM��j�� ƢN,��{.����ɏ�ɦ�쳦��������{�셇jNAE����޾���@���v #��_B�bW;	>�J����M�˓Dz�0rO2�o���o������H��;�7s���c��.Sh��2A2�D��N���Fk�=��*�M�[�����1�w����ۑzG?h��O��E:M�`��m����UK�}CI�Y���&���v���ټ5�(F�arwt�L8Q�F&+������zoFB�q� � x���c���8���k���
�Ȥ3�g��1�sh&; �-:D˳2�h_S&����1\%(a0� ���qR"�\2�2�MY4��(/�F�~�v}c�E��%�ڂ��Q���e�S�rP�\I�8d䳨"�O�?��]	2�$�����D����<�C������ҩ�v�HYz,��Y�8q�����v����!���8�r��Q\4ԉ�jX��+�gst�:�Ze���U��B��V��%g����J�K$h�u��&i ��N��F���i(�P�P�φ��/ ,�g�n�J���e"���B�B�*��B�&�_�$�D���T�OYDY;�f�̎_{��dT?��u��>�yƱO�qYs� ����bF�q���=�$J�1��GD�u6�	��;�+��&��LO�N�����\��>}�q�pR���5������(w�x�,&����Q�/��豆/XP{��x�;�@9���\z˒���O����Sh�j(_�ø����B�Q�PN����(�	O���˸Kp4��(g�~{������v?���:�0���9{��9r{��X�h��T	BG��&� ����\خ%V�����H��0��e4Z��i���1y����u�e߭��E1�9�j�饟������y���a��
���"	2$ g�z� l)��d���P�1e�C(�a$qb�� ��?�!��<�oo��W;g���@����l�~F��X���B{$U��x�6��C�L�����xH���8��0����q`R�?7���O:]�8�(tg�$
6$�����MH(��V�PpF)̵(];j��B�Q��5� )��� ��Fx~�|[���Ұ�@�Qr�Z�2nC�%Ic��]d
�ӿ��*)pEr��q��L&��!��I�O��X:��"ZȮ���7-�*8�Uj�L�ԡ�j��G�=mA�-���C��uSD�2xg#��Y�#���J;��ŧm��K�����2���'�{J�c�ծ=��-����I�ÝHI�x��/������������+���&�!��'l��2�\�J��?��uʁ�R��L��U@�$�^[�T�>fj�����j��P�t�̵a��Omwa,�w�& ��3�7X�6�����zW�x��/�j.f��2�x�D���F
��	�U�P���`7�ef|5	W��x����z�rR�����n��!��~<ϣ���c���;�r�-CJ�ɹa������vW2a�fx�T÷(�'��r����5%~N�1¯�e0�>�,I�h�F_,<$Z���}Ia���N���ZצaQ�Ȝ\F��7t�=!ؒ)F ��h���e4��|����չpp�	�$�Ϥh��9A~����"�܌��e��*�v�e��.�V�L0� ���첝}
�7��Y���.���ׅ���;�
@2�)\��E/-��;��&��6,\c�¿�x������rOi`D���� D� vP1�A_����j�'�Q�>*��+[(O9K��5v�0�V�O@+��ۺHX?�|B�ț�x�$[?�tV[��G��=�O%h��=��R����������7���o�s���1ՉyS��Z\������3�X&+M��4�������I	 p�%�1�S����/��0�M]�Z�i�7�脐"~��KR�w:����u*���<nB�3��+v;x�^1�2z(۩�S�B�� � ��Z��̝w���j�OC�� ܘ:M�!8Ӣ3�@ŋWw��QE���K
hu��<���xh�5��B�M�xn�^��ʲ��FHb�6P�H��ʉ.nh���Y������̸�����2�Adn�D$dy_�y���!;�0��?�WP�P)d�'��H�&%�'�>��X-4��sB6u�Rqn��f G�.%S�Lt��d�~��X��KE���6��bW������ʘ<�����G^��ea�󓣠��U6!~��Վ��Ц�����0FL��?�����O��ľ�b���m;m���T�����!�l Ruj1�-�f�P�a����'g`N�ܢ�DYjFn`��F��l[xϺ��;�*����.!$��D0#�ѓyDA�� sM��s�po�_ �R��-�m�5R�}��R�;~�F���~Y@)�� ˳+�bT��A�t�ƺ�kʉ�
�ͼ�NF��2�ݝ1)ۡQ=�lH����
ђ�q���pk�Ci�&ꣷ�"���-��%�O���5���,��E}D�0�v��T�@d���Y���$���OK���[��CJ�r�Y��=8�v\����-]��Hy���=�=W�akú1q��-�s�m�z>��O�t9.�}u�䅽��������cDPF�.+�b���%z��*̂F}�PCK�Q7�s$��d��_��!&M��d��S3U�C K�����O������/��G�m���3����1m1�V_K*����V����a���)+��c���3�l;�B^�g�!h��V6��R���I���;��~���s�̈	8����g���=�P2�{2���C׼c��[B#�48��}]�I��M��ϥ�
o�^lOT��
m�6u{m1��c:{��1��=���̩�rn��_7�{�r~=փ�ch��'�˴��0
�rJ�j$����%;��-�8ޑ�li.Z�0�c;�y�=7��f�,��CIv7�Rs��21/p����ɪTI����e~��
����B{/�#��wH���*������Y��wK%������Q	�E����#���M����
@8�#y+�A7��/��v�-�Q�` h����Ee�nY�굿v��C�hK��5g%��U��(� !��;��U{ٝץ*\EK�5�Y��O9��-JV(1	]�0i��.��c�nD�\�u���u7S�?�	=��c��Ԝ�2	|���S��E!J�N�xH���,���Uv�H�XR�ׁ\���Z��Z_5 ;hd�$�Z���*�J��Q֥����X�l2�FMv�Yc�t�c��P��\� �~(0�H�`�&��Y(���`R@'�sQ��2�ֵ+O��gx�3��+n�������������l֓IᰫǑ5����S�	����M|�J�}:�7bۆ�9���e�P����*ZD�$�f�]4�9���4y�0�8��a�i�$�ۂ]�e.�z��Us���Vq�܊R<���`Ȥ[>65���@���������.�cX��i�ە��}-؝u6��k�%@s\C㣘���UR4?���W�-����nث��&����R>�"d�5b6 �Vr�,lE�
*͌c,�GSik��Y�D}Vu�$��ۚ�����0G,w!�Np��E�Z?�A,�vBۘ�U�[~�����V�rA����=L�4D�7S�k:n��{]�'�BXԔ�?=����<�jT��ϕs��H����5o�E�Iџ��������"�a��|���sJ�f�X��,�jI ���<oѢ%�� ���b���Ͱ$��٠�a�����X�ޏ��=d"���s�'��H�����]�/������5��j�b2�1�S���R%���N6��vE{��c���9�h�bHh�N_m��7]K{�L%J6,L{IB�L�KCI��dZ:��ǫ<{o0�7�.��;��%^�J:z6_�0�U%�'�\)������ŭލ_���41�LA�'��gu��Cc�jW	\0׌b�+b�J��ىV&�����4�\�Hc�æ�����X����/\<N�^���&ѿ�����M���Sέ�grm�x,��;P�&�z+3�q�S:}������}d>֮PH:v�;*�n%��=-l�7�j'�o.�eKd��հ݋�O�U`A�ʎ���KǕ�G���a�\�==�ro����{Z(wIj���z"_�Z	u�9����o��#�ꃟ�]��������(v��y��C*��֒��5��9z�XB��!�\�?Б"(���涿��SOQ�<��e���ȑ�!����>�Y��P��3�*����am��[_w����rӹ5�YİQI=1������֌}�^�{����L��wɆQ0���HV�	Z�K~^��$z��ͫ��0!H˙]-��R���ue�öߍ�BwІBԛ��mQ���N�����[��>����V��$��#�y��q��[Ǉ&��@��K�i�V7�����r��?g�n�'��B��2L�"�;��r��V�w��[O�9Gs����44��[ǌI���>�,~T� �����N�]ݛ����~�ZR.��DB.>s�R}~��"g.2�u0�>����o�&��v"��<��[�,�}���Z���ܾu8V�F�}`o*5����uͳI��g<��h!Z#��{*�L3vb@����ד_�"�'i���v�xM�.O�i��5b�}z�p�MI~z�;j��ca�p�%����÷Z�x����.��ز˗�T4��ɚ�]���$�8�14h`����N���h��Y8����wB�L�����#�y��c�E�Y��!)FD��/c=��*�1�lX%�>�Mq�oZ���T�EAZfx_�����\���V��r���j~�ߒ$��3��?�^;{$��}T�6�XG��-6.�*T� А����Ъ[��>�����SmA~~��Q�^��_����D�fS"���ިo���)� A��RB�21�����M�a'�ݳ	F�S1�x9_�'����z��xϞp���9җ0H!���JS:��W�o�hk)�u�d�f��T,���5��T�$��خ�2��4�9!G��,��z���I
R��>E���D7НϠ���3�@<�L0k�K;��*`DK�^���I�N?�wn���"Q���'YY� ���я @�P��t�ր�g#�|�?� ���&uᅅ�D��њa�b��>"	�͈���@eK���tdcq�mA[�R|"6Rs�t�C��(,���F�H��\�?I2��fW�p.��c�<N���} �<���zPߥp.�o��Iш��z����稳0��@��Ħ0���}��+O
ZVT=1�G��9�h����S;��J���Q��V0� ��I�|�뉏�4��r������Ӳs����u[��V�5�y$�ٙ� ���[=��)�t����X�vo�:2����5�N ��N�?��u�L� ��>��ܽ택����#�,���\�d�XB���G�7�d�����S��Y�[L�8l�6	
ZT�����4%Y��$�w�{�Ŏ96$���%����1-�4�&*�K���(⡢�
fI��͌��<�އN�2��˺�G��H��T �c%r%��eyCLoN�z7�G>�ZEG-�ԣ߬��Ѵ����.|߸��##�~B�һ�A`�5��3�, 4Ԥ�gP��ʛ�-e(����+�����T���E @aB9�0�� �Ĕ� �����	�w�6z��!��]U�����h��D>��8�գQUиE�GEPL�[���D1���'��KH�������ܹ��I��3��i�}�h{��2i)v䪿[��qྐྵ��)�i�k��Q���-뼣�P�4=�LTn�1�����:ўìD{R�o����сC4�>}��/�J�M�a.!�R��E�e���ƮO�4{��q����������j�P�;����X�����w=~�X
w��<'�%E��X������Y�&r$�՚e^�7�:v@,��pm��۠��Z��'�Nb#��'���Ԥ����)�v6�Bɰ:�����SU�]�d�jP^Wh8��#(\tZ��߉��^/�j�����@����剙C;Ԃo B%
��>����E������d���}=��v9�w9Ƞ#$�;��o�/�QM#�?�שT�����y44
�I5��#.Ò�@�^�:�+��f\�l��~%#D�6�Wv��X����\�'&5���ԑmY=����-
k:�����v�;D���i%�"�V9p��+�0�ؾL�����)��"u'�պᤉG�y,EcJZ�IGc��1���,��V}ՠ G���b�.8A�C�e2=��\@�x�4r�P}�;r�@~�C���%�Y�D��gj~�(�-�D9�y|���� ��Ao'F�`�`.(̃Y��ǐ�k�4wQU��(��*���Ɯ��Jܔ��1e�_���^����q���{��{~�C\�0L�����6�߽[��SS�<�����FE,�R'���x 6/5N���(�W�W,§��(�O��\h�Y6/��h�k���R1��ޯ�uPD�#����K	���.ţ�¯l�ws����ut��R�{��[_��^��2�M���1"�r� G��Mb����_�3�G_[�B�B�
d�jt�B��9���ۅ�#tdH��s6	�����A��Fr�`������a�C&�ِ����03��`��$M�zwY�g%���a��T?�~>6���`NA�k����:k5�s��Y*GP��]���;7u?�^��R`�����*7&�x��t���L}��w�9�>�wFO�-����o��ڸ��T9�-�M@�}0�6�`�7m*DD�v� o}]`ꯈ[]_��J��C�;kp��|���<}�0���r��(Q��X)�Y��R�.�M{�Y�Se\Yʌ8Y�j�]��h8�
�@��Fi�o�������"0(�|f��w|�؄�+���7?/��luQ�xz��E�+�� |�S�Q ��d���l�h�r\C��Q����w,�{�-X����yn���� MLVM�η��O�էsEbBcd�a��]R�K�Hg@O�*�� �+�4��)A�_�{�7���YW����*��#{Կ�l4�Q�ǵ�(��=�A�ߚi�5>��,����B��%�j�	�^v��//�>��x"�
��g�5�������D�i�H�E0���)仹u7���9��ɦU�VU��lG"|��0��a�r��t��������������zʌ�hn_7��,ك"XSĐSl�kɩ&2\��