��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+���]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�O'�yz,�_ ���)ZN�6��dQr�p�x�y�C'�m��H.@'�!ѽ��Ќ����Mڨ��˳0��`q�M�'���2&��Ȯ�W�4��д��|�6�K!b�'mY�`��L����Tr�AW��:��3����'�v�WM��=K*��1<��(t!�1�l�<M.�efvH�\��0V(&��2��j�P�cG���J8�|�ݦ5���'J��I��/���� 9�	q�Ϻ7����5������(����U1v����V���W91ƞ�3^:�)e���'qU)�j7#��ME!A�W���$?}��~I6�L�޾�v��}hK���) ��N�������65�n��ī��7�?|��q�a1@ͫ<W]�M�Q}�?��;�F�G�������E��F��Kz�;@H[�:SegD�2z��B������E�7k�l{r�d��aߪzr�PU���|�>~�!�֚ �ߖU�d6oOg ���	�:���fX�پ�����4��k(�ީ�*n'υn�	N�A��5��Ap&�28+�1�r�W���-�f�KYUs��a����qɛ���*N�Z<�
��l$�`P�M�P}j��@��b�Gx�yS;�,��'��yFB0?K%t�(��ڸ���"��c�8�<y��Ah_�č|~�>+S��hb�����J����.�`���ע�e�D���E�HY�L� `t��� 8�.�`[�ra����~��#�e�ݺ�/��s�	Hf��:�D��������gK��-'��������l�m26�׈ w�R[�?b���� ��=��i��T2é�3���ر� FW@�`�{��w�,�d�R���
�O��<O0t7��-�x!�'{�eQM�u�E������Tnh�w=�qd��^�>Q��a_�#3z�8�]�D?�zV��t0Y,Y�d^TG/��_�<CV��|�ӷ��;M+'z{b�e�ED��-tp;̔�*.	�j�{�Y"�b����-r��.k2�����Q:�A�J�$�����";��*%�����/2��V���YG�H�;�ƺ����+9�Dq�� r��1Q�jp�����t8�K�H��(j�+�{0H����;j4JR�+��W���ȃyPI�^)��{�<�͹��|��1Լ� �64�l���!c���'fa�AE�n��hh�(��<P�Zy(��E`-�0[I0��@��>5 �N@��%��:cj;[==�EM\&e����c���u�`� ���GJz��a|���n����c�UIQ����%3�>{�Kmq��8<
ȸ�M�]��~����8�K�(6j��u�s�t6���[��V����Ԗ��إ�^ul�C��a�4i�3>}�\x[sbTM��P��r<�v�� A�[&"W%�:�+���LY߀�V�������th��� _�J/V�uTD57�k���;|{�����+_/��o{͓��h�۹��"
��O_�\����)�?�)��" ��
��E	e�x�P�U[Cm����r�;C��%p\2*���,Y��l5�u��D�����:��ش�-�x�|g�@s��S| ���w��H$����^F�G/gv�=��Ҝ�K(��%�=�p �f�z�p�D�s�"�n�D�[�EKJ������;�ߒo�#A#�و�u���#�����j.�D��_�P��<�zCgz�M;�Mҷ>��j�pdS�?��m>?����RoK�d���D���!�ܞ�����#J�;w�� ��#vnH;%5��j!�z5�B�n�� ,��Eŋy���bo��|7��B�l!ԃ�<� O�O"E�x�F F�Po�N�t�%+��f������	<9��t���C(5����a����<�h�;��لy*�mw�" 2�]ZbgЁ�A�Y�}p�9~+��f�F%�;��H�y��P< �$��f�����-�/����"����9o���@Y:��S����b�"�Rڶ稙�D����gn���sֵ�G �<�#��%YIX���A�6w�PW����0�@�e�Z�qfq�=��c'�!�}IPOe��Z�%���}�� .���B3��q��R���Z���0?�L�#��L����w/rL�L稽��똰1i�~!� �_ 2\�}OƦ^��5���ˁ�
HI��N�.���f����j�g�~�Ǻ.ķR0�3�$�8�G��,��@06�����VRy���+{p?O�R���!���E��O;�2���R�Y������Lr������!-�$5���U��r� ��኿;�Uz�x�����O��1�Z���_���h%��~W7r�!"��[;K�@�Ǔma�i0S��-c9��Z�ne{���^��Nw�J��]Ke6�V���}�J·�w/]!j�!{���E����Z=�.����r�xx]�o����S3�����;U\^H���B� ����7�8�*-����N�n�L?����y|w(w����h��Zy�GG���#8�P_Ў���s��0��BɫK1�����I ����i��@R��O����ל'�a��5���U����KM{�����^�\�	Y7��ڔ3���=�ښ�B���@*��AhS�!N�h���tA{:
���H�"��AOޛzpp��M��:hB�8��x�z�S\��@�: ��6�ܚ��j���C 4 ��ڡ��}�sƼ��3Z�}�d�zqx<�cK� =�b��'9Of$J���'�n��E�	�L�U��9��赗���ʌ$x���,!�E�F����y,f�`��!����/��n�iG�R_a�%���L \��]�:J�,�d����N���o0��g�G~abd%� V���X�Ҙh�fhRw�u���4_t.��|m�5{% `ֵ$�%�<�����+�B�/m�~�}�bahG��Y����.+g�- ��БD<)�/ٞk\r�8��pʉ�2�/.8��uƙ�Vo�3�ք��n�X�ᆥn�VQ�:��V����{��+�c��<B��/#TA�B1��G!(<�.��{�!��2�'�9�2���4G�Q�*9	"���4����m���;N���F�6�֧�mr��Y콞e��}���*\ұw�Z3�e3��;5�h�����y���p �0���j@ V����v�לBﻟw��S�c
�r`��e�G��&�U���o���ʮ�9�����+���0^�}rv��Id[��]��D�u��� �[�IM�ٝ�4L�CHi
k���yj�.��c�r1`��2���-۳�v�����(�cw^�B �L�f���[����/J��uɰ����m�K%y����rٌ��v�\u�l�R�V��l�Xb��8=7|�{N��B�Gr����:q�#m�ߤ�W�(��^!	t��.�Y���?@�1���X�2�3�j��z���&���5�!��E�Z�=�Z��wQ�g*c�F����4A?�ʊM�����SXZD��c�ws�ؑ�T����ЄF6�s��~W>�m�k��J���R���X���\���gZ]�7a�q6�Y��T(��uR	ؤ���tsf��K�F}���L0e�;�v?��!g��~��WC�>�7j&���;�;�Cè�=��
��#�6�H��t�&]��G}��(c�{�sff���հj�ƥG�Nn�����!r8�4E� � bNjd�ZVhO��z�����D��\8��&��o��j3Ӕ�b�.i��M�w��j��ĹE'�n��w_שe�HX�)���͸�`�����(�N���e^���Hv�yQ+U��:6]�v��G�0��n�uB��]]ُ�21x����<<�).��6��qy��U�03K�����$��+��ɂ���Zo����S_�d~հϳ[�q]{���K/鿏?F��w����_EL��lb�`�`e+�A6��]����~���u��i�<�(��B^�೗��9�C�]��ΰ����	TI�FwzH�>���B�Eh�q���T�a�Q�R�飜����T��nu�W��ݝ��L%��\���*�Jҍ�7bơ@�����|K�!�{�uCz�j^�s��?���n6*`&di�+9�����+�9�I�0��$q-��؋"��E\��D��p8֦� Y��7�����A�� ��*�ӱ��ɥt�qK�d~V�Zw��JՐ�@mk|Ex��I�m��-�9��JH��&^*�9X��G0�'L��-r���I�uČ~��/%������֣��V]V�H�j��D`���²lΞ��O�c�8�M~�ō�m��ªp�,�ϊ�ް��0i�e�x����X��VHz��P�ɜ��yA/�;k��'q���H����.܊�?[��;����ڀeR��կ����X"A���U�ܜ��蜼���qʂ>ߊ~�~��8���1�U&���j�yd0Z�m��ʵ�^6�씝��0t ��U�ɉp��� ѧ�%%7˖c�5�M,�5A�jfUb8������	h��e�<����pȔ���Qf_e� ��y�h���$� H���d�����#ŸV�`V��E�IR�Ӑ5��3ԌK*B�ȆK~;�A�w�_"�g4���Ԯ�I��?�^�
��
ɫ�J"�^�QoX_��Q��Z���c��3y������l8�%��d���w��	�X������rF���w�B��!^��'<���JsCߵMŘ���K? ��Sѽ��(���>���1�&�/��q��v�R�F�7R*�5zŚx��I��K�b��N�\�ْ�q*�C�**}�a������N������f'1V3W��Ψl��Lb��X�[I��Ч�O���'I����3�ue:g��ug���j��R��>��ʌ<5�T�=�SXZc�	��,��-$���"8z��5�{_�$)6����4�ƈB7��W�����V8&�G�3��*��g$Vǌ��M*F#��t�����i'uR�i���"�5���D����{�[w`֩%4����P��w(��^���-�	��0��$v�<��aCݿ
�C)֞U)3"���J&$Zۛ�u�p�.�I��{v`Q��+�j�\P^�����[r�D'���#�L0����/�o�_ɗ����bw�0^�̀�;ʃlv0ı�[���V|ûC�)���؂ǲ'�{¦���/��qUҖ_�B�����i���Dî�:Q]�F���-��`��GS:�¢�*�@gp��uދ����B
V Wf��iZaZ�ɶ�f'�n���ϩ�xP2�ZGtm;�l	��M}x[����~_�+��>b��^Y�BcD�L]Ъ'�0@�����Tׁ��A��DGL`@�7�3:�wL2�(�]��2Et�[� ����U��zϱ������r��%$+z���牔cC=�tI�I��>el�|JC� � �?���-��tm�	����e�Z6P2� [��'� ��r~#̉'�<Is�|�&�h��U~����˜�2@�R/b�po)�s�z^` ��W±�������
���I��2��CeIsK�j���ԭ�#޼[#�B[[�gp;
<�m�y҉~��CJ�o�v�$�w�W> ��=�߫�y�<��Wv�o��U{"6	c;�7��߆�O|0��7�����JS�������"�ͩh	�ò�sx�v�[��� �C ��" W4�
Gs�~�wJ$�~���r�z�h���D�;�D0�ը��ɢ<��4�ш0��9���Rrѡ;�RV౵�dC�x�l����=�H�Zb��i&�|��-�,n��)I�~�D���`uJ1�9{@��M�&n�7B�A�y�Uk;]g�W�4���?�d�7�U�D�`��b<��̒:�H�xp��*{ڝ9C�騱b��c�)s����ĺ��V �����|
&��,_FC^�4�I6�fr<�G>�f`�T�p�������97"�)Yh3՚h�n*5V�˵�E�2��l��պ��4���5W����қ��!���].��Q�}n�O�Yd'�:��I%�Ҕ"Ǝ≚s���ո��4�bC_S���ysԺl��^=D��±hr����Ȱ�߁�V8K��G_��B�����;�+��� "x���a̛�;ڨ�^qD�`�����K��ky�`_Q�����GY-��X)����t�rެ�o^��������>���N8�n�́��[��P����g�K>�!�$;=�AB���ՙeT�梵.�)N&j�Nю�,�k4;B��:�/��G�w��8%��iC�k]3!�\q�|��(�~e�}H	ĩq���cU`B���Du�\����=���v����t�f��d���C&�9[�q2m��g9t���TARRw2<c}���V3r�����5�/�w�a��������h�����W^�GVO�ްPsb?�&��ؓ����nx(�M
aA]!�J`�8���	yY���� 𤯧�ᣲ�I7��	3�O/�#1��^�
L�����{���D��p�h�>f�����e��D��6d��:���.�\�Sڪ'�����N�{����X.��#|�5��]`�l��Y�.��@�߫� ^Rh���	1f�C�1�`�*�	�Ehd�M\����T-�H	�5>-S��NI����>/��<��Գk��񱪨�(�U��(�g�����#&�jaz��i3��o�!zuU����$�P�:�I���(�K�[��P�)8<���2��(�����u��t����	�dHg=K�,ۤª)��'�%xf�}�°Sl�ϲz�h.z�b�#rX$<���洶��sQt���/�)� R�7/	N}��^��+8��2���T'��Oc�g�h�Jy�*-j(7���S��Ժ��6
X��Cr5��6r����UP,&����0t	$=V����7�F[�G�O-��uWS���xSl�+ݲN��֩?���G�������PN4�Er���47�I�|��s$ߖ:���*Oqd�
�<Mqp�