��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P��v�"<ߞ��&'��k%P碶�R�ӣ�sĞ������FY&	a
��#��X��R��E3a��2'��R�@0K^�M�N�����S��u_�ƪ������W�f����>U�`E���NK�g��5����k��ʀ	�+���bT֡l�#��F�ݟ��8�5IS����iɯL{�� ���K�{�ݑ~�o��vh�=���'�d&@�(&I ��=�}�^�̵��l�v��h�7T6��@�����XZߩ���H{]�s� �����P�I�\�9>� ��"�V]^���7J�j�A�	��{P+��;��IVP��m�,�Dʐ�e$�Ø0�@��O����V��U:�������:��^�ͽ^�$v��8&�&�h�E�w}�@���uOQ��W^���A�c�NҲx��+�mQ>�c�	���`�:�����փ��"[�j���X�k���x|5��0�s�`��e��mxW;شA/��
\C�`�p�O�U�ҩW�~^S���G
��<��Kl.�2o���gu,�Cvv�&'n��c�����H��������?㩷����X����`]�/,V����Q�^�3�3�駌�>Z�vElI��eO`I��o)���.5Y�"x1�(ˠ'��rJ���:䫞�l.$.eg*]�]�����IaC�����^5������~a|B�@�9o1��7��7��/W7d�oH����Oݑ��h�K�@.�����]�
����@�߾%h;N�y��\���40���(���>S�#;аw�eZ��˺��e� ;���3	�e��㵺ϳ	�LeSќ������Բ�K�b|�.[��
��Ń�fd���]��7� ���'��J)�i��޹2�I �
�#0��^vGJ��ί�x*��S�ĳ�ԓ��ֈ�`��iث������h&$	�&}?�+Gբ̈�3��1�yG���u��Rg�,��D�~�^���c^;�u�ȭbtX@t�~5Z��60���Q{p��`��(p�m�����ML%��A�ho���7z�*yru�f܍�]]/
dҕc���sGp����^����2��Z��_@� �w,�]��Ǣ+�Νi�
z��"�}d؈g:M��gzWO3���/�>�&�؞t�	[����߶_Wp\�p�-���h�!8fvc�>nG�yae�Y�wꖜ�:c�$�iC�J��lϱZ:��H�
��������[�[ם;��0�����ۋ�Vs0�v�b���?��UBfw�}H�<+s�0�G��O�,����?�"���5��m���XE�܀%e���<mDg��|�+�"fr�����R[L���/f�x+ TS�<fwh�f��^W[�-��q^!D�-rQ������F��h�a=:��D�	x�����S#z<%�>���q�XM�����m��>���RHZLO럏U�N���2�g6e�ߗ�=��u�$���g?�m����t �0�8����x�(� ��Ja�B�%��(@,�K05���RE���t����=uB��EuS�B��a���+&�7����9[~�Eu�|CE	"�n�N�C���E���Q�W_�K���:k�*<��y��Je;Vt袡��)���b��%�ǟ�& �ν0����:E�w��V�<�TPӟ��
�р@N�uP$0W�G7�f�P[:�T�6�\���K�JS���L��j�[�M��4��(����a�Ǐ;�'j:��2����|�@l����ߠ]:���Q����dK�(��4
������=Ԁ%�������j VPZ�,�!��!ݱ�䚉��⩼&B):�dí�Z��n�w�OEV��n�`KNn��O.�'�TKM@���<Kv_�ss��a-�K�D�{�'�,	�A �ե�,�^�l�NB,P@\�A���H�W�I��
�����`܄��3�\<L=�}��^�-t�1��R��=����Xv��C*����ٹ�>�%rG��@�Q�$z��	��&\��qX��'��賏5��tM�e��� �yL������Qxhm�O����!�QZ��$Ͳ��V�97��Y�;�d��gQ�(�~˒�7������Z������(hc�l�a�.F����p�Y΄���.0Ϧ����_��{�xpg�?1��Z��f��^���4x0�B�E���[�.�g�0_�"$��`B_�o���Ǻ�;q��Å͡����շ�W$�O{A2ɲ!���#�eD�?�%��
�d�E��x�XK����vl�c�[�dݧ���Wt��e��4O�}jg)~2ԯ��������KZ�h"=\具���kY:K�� 6V���}�	|7���A�lDF	DF��O, ��Ovھ>	T�B�R4��,�=46NwC�M��ͦ�M�3�G̾6(
R�c`+���l������B����r�n�"�9Wj=�����MA1��k*�v�dl�W��'��ft-Rl}Q	4f��a�b�m,�X%�aZ	!;�����x�GUM�1qe&���SG�Le<�qnB=W�˶�vS.�I�o�X�S���C�=աJ�I� b	ב[TSp��]�3;:��i��ε
^�$�5�&�a�Y�5�(�8tkiI8Z[��>	�8T��*;6��V7�����-v'�������/Z��<}��g2�9�Q���3�j��c̠"�rˈ�+�̶��ښ������k�_�-̬b,&��Ny�m��	�����'�	�D�NG0US��X���>�<�+{a��;n��/Q�8�%��(�Z�2-8����'67���(7)<��	�TSL����s���co^���򳩲�,�ͻA���_Y�tz�d}i� 0�d����0_�Pq��A�֎�	��)^PX޺7�}����
s�#��!G��g��-ȢZTL�8�"1�Fg��obx�Q%$ �f��p/�/��n���XM�n���9��C��:����A�f��]������ˑm�C�W��#P��Op�`"���)+W'���8���~nڌ�X��ja��*�Ea�v%_���xց��ؼ�6�Y�*�M����݈��-��&pE"e�:�&��l�e�Q��ohJ��B�N�#�cnB�>^�u�-�NiL�a �nB�1��6c�	�T�dp3���}5L�̑�7Yu�o��� C�b H�+:�f�OJ���\<mZJBq�/���B�����=d%p�- Y��	rD+���WZ vז�8�a+g&���@cT�A,D	#]>5�g�gA��W���|y�b8ɠ}���/r�O7y	�Rb�A4�������9��&�a`?q*�	�`�ɰ��δ�P/�li$����?o`u��(rŚ�!m_���y�m�?����y@A�p�{�Q��<�vQ��Vs��Č���u�[�ց�^���98�/4��3���ۑ)i�lS��x
E��F	S�Զ<��t$����;��Ҟ��Ԣ��%Yx�B��B����� s-K�ϱ?�J�C��xH࿻9����Ҽh�&E������vQ?�9r�F���u�cDs��l�G�x�i�x?���Wm��*�)ձ8��	=-���	��k����TVI�Y2
K��=��L|�ϟw��0�5�7�O�<�z]��b94�S�f��
`��	���$?���'i��<��;K`.�<�EO�mP��|K�����-ꊮ]���+�z�9�x׈�5̳�Dd������q@���N�)��(�
�y��x������VO�A���ʓ�V�nz�B@R�s�YS}�_�\�r�&*>!"$�aӸ�!��8�����M�O,�|o�{[��þ����`�R���)� �zV�ɛP�)@ƣ�X������������rG�
�qv�K� pN<�[6/���U�h�p�����C���0?Gv�pά�H������w�F��2������Y�A�죚,�16����Y�A}�t�l���˖W-��oۧt��:F`;�ё��5V�6̿��D��m��XÖ�#��ʞ�<��@��e�$��>�^��}��Am:	m�A�X��0��y�A��į�<S4̅���Y���=�Y�0�b�{�k����j�Nv��$��8Y�|E�l�r�Q��[Y�vO/��K|U��G�[-��_�o$"�V)�W�� DL N���d��ƣ��1��gjTН�wm�����O��k�j�\k�_a���f� ~�v�L�t������fe�XT@��	wN[	���^��|������B�3��6]�*9�L��Ѿ�{��m	4i,�A�]c� �y��F(��W�#���#4�
��`(�a'�&���Y�*J �
�F�/T
3v9��Asa������E�ap��E��?�C�13y������b����vv�0�5���8�>��%�>�yC��[m z��#��j���U3`(ѳ����@	�z>�Ր��npʟmJ���MJo��_���,���8�F0��T8v� r~B�����IV��Ŋ�'���{�ANM{�{�Pi���g���Tp@���ɣ"z�wh>�}ޛ^¸�y��^$r:���9X��@{�*剕'"x���`j�ʠM����r5�����3�X��y����b��	SP����{u ��[���k ��y����[��-y��Z�ɚ΃�KB�e�q�p&��.q��.�"ioԳ�Vbs����f[�l 3�Hw� ē��sy��P�op�E%%h�= #��:� �p��б$Rq��BD�?CAǡH�+"�E���Kڶh��N[b���V��AC�,�ݢo�+Mj�Z	������)�z}�!fy��5k���O,��A?�&�j{�v��-�|j(��ׇձO�c�E+�Tԁ��@ZgX���x.�K��]���s�9xWӀ�>��,��d$F~}w�/MX�0�}r�tXn��.7"	9�ʡ;��-U�8|�+w;��Ռ�~\�^"ɔC��_]7a�1P��P#���6jdU9@\lW�%�!��R/*���fq�3�ě�bqrS�1O� ���9�iE��Y[:�$뛜�����B���/L���*��/�,��P���3��r]2��Jwt�L��1���8�L��_[_hU%�j��(gB���Y��?{�	��c;϶
�:a^.��|�d�4���?�=Q]oء #N))f.5](z�*7wDǱ4�#ķ�3�a6V~rq��Q{}��
�A�E@��b+�}L���1֝�Jq9��4�7:1����~��||Rپ�l�Q�P�|�vu��N����,��̦=��߹Ojq��\�~�<$'�Sж��� �]��Dn�E�Un"(r�^;/gR�dͬ5��v�Q�ƻKUV+� LK���7�=e{Y'�q8���ғe�	zh�?L(� �q�����莸�Lݻ/-Al���?�Z}ZOI� ��q�įM���a�%��h	�>���-���bs���ڼKz=� �"C��{a=m��ْP�1��b��;'���="� ��V�|ic�,S�.x�>ku� �Ĕ����`&�uY�ȴ�z~����@���١�G����X8������ʡyH�3����sf����g��Z�^���ge�{�o6+��`@:&6���?�{�M7��8ui�-��'+;q��!̱#�}wAC�S��G�$���F���O���	:�:��J-!�A����U���S��W�|����E�#�e����X�Y����� ��5��D�}�ԥ5��[C\��a𿅡	W�2e���@w'�>����s}��^�z��بG��p5-�nS��.�轘��-�4��),�:�@3&;w������$ >�����d��͚��f1i����ݯ��v���Kb�� ���A~}�Y)e��GʷP�G�8�n���\�b�"�/`��r	�R؟�P!hd�W[!�-���[�*�[�!{�&G�����mqDjtj5���]U�����-�C�Kӵ7�$��^���k��y����,�8�tz���r93��E�䋨��Lb���!�ͨv���q
�T�uwf����5J��������)�°>.Y,���Ԓͨ��]r��Bh� ��>��=T�&���ښǌN ���Y��*GS�-,�o��%5db�w�p>�#���rJ���^�8�2w��\���FK��C_�q��g��Ɋñ���"��T	qwFu7��~!��K�Z�܌R!����2W�W��x*&��}rQmi���j`�1$@"���ՈԢs �O}���0��v�{���ߴ�c�j�jޒ�\�6���颞X�H��'	:z���YG����;���e��'~��7�f��CEq:.f�>d����2'�
��`�A�֯�Z0ӆ�Ķ����Em\T-a��;=-U����vu����u��V�9X'�0T��� �La�:��+r�6����84��z�52�%S\�x�R��*�fw�)�=|w�[;�&�o���[�7��x��!s���Z����ڼu<n�h+Z�#�t@l_�+]M�u�n��K�k�L���{f����D5��c��5��0�e�oSM�)�T�ԗ����.W�X9ߨt�vj����.�q�S�� '�p�Ϋ��O)s�%�1YO����=Yᐽ�����8r�ɞf���%��Vժ�e.���'D�ā��c��@�͒谎����Hc����Q�g�mj�r`�HB&?�"l�@�J�Y�[h�:�뜲\t�	�mt}�%����u�D�ž!|kk�b�@R;4�@���8������;P���{AF0��i��&>Z�fò��e�E�3ٽ*�M��7���JnX��*�	���E P}|�@�����(���+EM��68��X�ك��
������ڊ���[wE��m���q�\]�'i��J�#���<��>��&��LS9A&r@*�l�H��(�����F��������}Vp����-�N=K���&�jU�����S����^\`2�|�P�y�q$���n���\���0a���i����-��*E\\)��e��c��Q�q���#�ԗ?,M��%!���$3�iق��c���0��W�/��0?�<�X4Ν��2t�ƓU���h���`��V��~s�V��+VI���2!�[m�U����]���)n��`=�(�|�?�9���~'���3��ȑ}v���o��4n"��)}���q���%�璟�F1+gb��2� �}�X�|G��҂B��j4�ө�:��dH�p�;s��ȾZ�a�����T������D��ϣo�%�dzuC�Ck�	rHd�C�$�����(��6E�V���nD���R�6~{w-(�H�zm�D.dq���i;��%��շ��V����EFv�S���:>s��6���qnD���I���u�gu��>�ZB"���y}$�Zؐ^T��I� Mn_��5���υ�&Vd�pf�"�r���]Ҕ�"�/~�r SIH�L���qT���ce$��c]���d;���ȷ��Z��E�Lg��U�Uh"#�������E0��7�m�u�/?� v����;�-�|�C��ݧD��p�'/^"�/ �g���F! O���la������K�����*����S��"b�v�g�x������T�w猝���R��ɕ���uHy���O�R���������7w�Q����-�P��� -@A�aF��o����(_�~u��,���S�r�]Sӳ��:Ջ�P�V�V.�6�1�_:��wcQ�}�*��$�<�̓�D`�����SR�@��R������G�l�z�"c7aCx�*l�6�|`̡��r�+_���&���($�仧$�:�k�ph����z�ۉ�����J���a+ �3�O�\m��H5� �Ȅ5�G����5ZoZ/��AI�Z��"�]GK/5�z�eI:Yk$&7&v���$*w�P��Y1*�O �4���7ne�$9�v~�@�n�Vǋ� 0���iM�g�c�yv)[�d���]��]6*�u� ӺM�`C��������j�s�M��f���>7)G�v���/l|#V�e<�f=4/�k��R�S`���b�F�����~�#3R��y�1H�B3O�I�s\F���Nf��P#��&��؟h�\�(���jy��,
�;�|��՜(�ݻ؉�E��I����>R�VQ)\v�C��Nj`YL̽*�;b���9u�h�ڗá�df��{S���������{�UY`*:ߘ<ޛ���I�+ެ�n��{������ǈM7��x�ɜD����oi�� �us�JE�]]m*D���ғ�4�ګ`ГM`Κ��4zw-@�fE���*q&�M �m����NL��쑛�5�x)�=��ڽ�0/�
�i��x��<Y_�aJ��% gpPU�o'4�;�=�d�mR���6�j�͔��u���△{
RZ�r��P$�Go5���0����xޖ��@�R]?����c8)�O�eo��Y���1�P͊q�9���A�-ѱjٗ����>��R�LS�t>�%^���j��'�kջ^�H���F=�;S�yt�}���%*L1�)M��5�R|q�gO{]�jq%��,4��n�����B2P�)/��'^{�4,g��ڭ��_I]	!`lbD�#T؋��	ʞ[��O��a9��{O�(���	:��u�"2yb������'P7S����9��5|� vElo�2�>5 uN0�-Z���Lw��p���פ[W�`����#��|A<�E�֡0��ʠ��&���4�w�d凳w�;��G�޶N0����@*�+�8�>��y �1�
�ݵN�:���9�nщ^�/+��X���F���=�ߩfa�\~�I?Ӈ�K�Y�(u�y���F߰�M��<�� �b�<�@:��t�uG�f�^�s�O���Ǥ���xG��b+ӝ�W��a�T��!jA�.�#�d������hM=X<�Z,�f�j�I�Q��7���|�9y��I�x�\�Tg*���Ω��{�zb`ič�#X�#�ɳ�MB�; >o�SV�����JS�J���>�O83�>{��k��"g�yD��ŧC�N,�1����ԁR)BV�.�-�j���S��gE�'�+��I�E����֭T���{z�������n3I�I����>h���]��a�g�h1Áu���?G�FhA�Z�H������^��Y�yW�!�ܼ�吝���X�K�y�^�CRn\���>����tk����m]#0��_LȕynJ\��|�p�)���n��0�U�P��8�Bu���X�)Ҷ��N9bh�gxs�9��'l��M;��u��BZ��>�j.=�?3�~�|8�j��C}7��������H��n.�	�׏i���a�6�&^��Mp�
�H��s9�p�א� u"�j����#g!�6�g�ļ������i?�e ��^g���as��r��#�--%�z.@p�L.�1�TX��A�aS�3�&�86��!v>�@!�ª�&�k�+A��\��Y]R^����z5lT܅yCVrl��]��)��ϵG(ŭұ�ua?��q�[4^VS�Pٗ�0j�bc�$�k�Jr�Г`��@R��4��JeU�2�*�hxp�kU�p��>���D%����ᚾ�!v5)6釬�Q�09��m�.�~o&�85�~�A�����N]�:#���S+F��NJ��å��+�ա/���(��Mc2�T���~A�,C�	|���ר��A���B}�� ���]K��Y�
17�f��b[��S�lS�4@����4S�D�?�)�b�)T�{Ig�6�뫴(*�BY *�S{�Q�V�O"�s2MF�]"\�ճj:�<��Tv��627ND�P������4��V��V��*�{�����w_�Xsn�/|T��v�����ݢ-3/1���v�K+���J���B����R��V̿L�E/ӂ���}�ZD�X�o=��l�]�x�eq���#�^|�sÍ�u�?DZ�&n'd���"m����|䔈�V�~* ��;⫋�wz�������dI3�ހ|Lu�k�*���zK��+b���|��@�B�_њ�1��xvt��8��s{�P����L�p!�>��K��n�8c6:I����@"q#�'^\��	��J?����qV6,�T�^	[�\z\1��)iTZ)o�}�`�}#nCt^���p�03K��lH��(��E�@����Ζv�s�g �_��_�3�`&�1�ةo�拓��IO�9!�c�&����(0�h��#ώ��QXr�����!�+�s�R	~��'��'�ѩv�{\��e����bU$ww`kVj_���S�7e�)�Mw����V;�mù�J�4��}(�#��P^�Y���������	�T���[�U�����F�6`�"yK�=��8�l�T�-;����@�Y<i����r7	�V�zC�%s����O@�e�ܰ��F���I��`5ߕ
�B����mQ� :�w�3�ol�z��Aa��NÏZ�����w{�����WJ�꒵h�HΙ�&���iwz�F�u`N�)�r���$8q}j�V��޶�}\`C�-{�_�����:��AC=m`Ƹ��9��bVV�Ed�q/�m�?J��T��<�h�m̤P�%�/�o��V�dȬ��|��pL�]�ZYX��.�hk��e��eu4lz�5�"w=�]����<$�Cpt�~��?��њu�p����N4e���Gk�9p{D����)Ps��=̨e�f-pyh�z��薆�=�`�ۜ�lг��O�FO�j2��<��W�Y���J��)�s{��"���g�Z�$Ly�P�}b�$�a�%R��_�+?)2��A$��$��
ħ{��b��y#5�i�� ��D���Ւ�E&#r�Jt��9�����k��̶إ{&A�|l�>�	Oa0�Q�5e UniO���s$��t|[8�Y	�X��x#km�����;�`ׁ�G��1�34�
� ���
�`�:�>¶��8�E���>�SUg>��j�G��o��G��~��f'p�W�1lA�O[�'�0��rH�@��{'�+z��\6Nrcv�$<�[�c�jVz�O�v�Vkí��/�P�հ�h��b�b�r��aF{xȻ{�<��@����q��T�^����y�b��ƉV���MZ�� ��0�%:E�7�OAp���\,��{<o+YgAH�=[�ʩtֹ�P�@��;w�v]u�������&\���� #0D:_a_,a<��.�/��6��L6=s@"���0x������n/!��_���>1\�$�kC7CME0-\1b�^c�3��C��\\2��� c����+�b�"���A#� �A��<J|����^c�}B�C5t���~��"f7:�)�h�p0�t�\u�!�r�y|�!�c�(�@�>���{CEt� ����bZ3�h��~� єR�W�H��gￊ�nў������y�>?*�2mѕ��[p��j?�j�j��7��z94�7b/d��T�
��>i괅t��F=�9�:��;����*ߡ�t���[<e?�Tf�xY{Hـ�]]�/�J��Q�a��A�eyRK�������R��U�2��p��n��Da ��U!���o�4��D`}�Sk�Ny�䵻u�ିh��
c��0L���y��
�̣{�f�8j`�QDZ
�����EP���_yۢ�m��1h=�m�}I�%��I�=l�ch��9�b�g̻�%���Oh<��]���tcOwؾ���h)ڿKk�P\s�F�,9��tpA�#O4( I���K����1⫂����\��6,���alk3��9��	{S7S#�jEL�4S�Xd��X�͟e硬s�&�89�qR_Ae��qP5�b3J����V2�w ,��{o�u�!�k����� ����flBr�f�gk	�rE���v7�:`�	�؇��#f�{��t(�O�hqkJ-��*4V�f��|�'c�������*��3�9_�"��s~����@�"��@JT6��I���q8�liL�UE�C��Uy6���à'����Lm�*����k Xyۊg{����n\�lc�A�T����j��@i�u׍��G裧�\�_G>�4�����e��0Iτ�ö�7�0������������m4T��g���UL�1�+������qa1�z��Ѓ�zJ�Ԋ�e�\H�� "��旋�;��޾�s����� 	�V	�g�|D�ϲ[�O�E���l �Ĵu���7�7�݁��"�0�q��.	O�T%^R+m�	MkSV�@E����N�b�!IY���"}3�X�q�6o���`�*R��{�<��;+��@C3�8��!��5�$��:8B��/���0�n�qÛ�Ì��8Ai���R-��d�_�>w����d8�֚BYs*�S�7�Ԡ���q'L��x��بoqioc���Oi`�����|,;�-�M;����J�JK�ɏ���@#Y���'�2+/\,�7��*�
uY!��YI��# C�Մ����|-�W�܅ 1�H��ج�I�?=h��q����f4�E�� 
��o)&M̑�=�;5�e69��u��t_�^���`���#�&q�_�$�:��� �(`#���Sf��2٬H1z�5��v췇J�l��^��� �"��>���]0oι~���"��(Q7��]E4	1KA$�Q�!�'��l�ɀ��N�>\����
F���@tP��p�$�g�Z�c��^�N�n��2�}
�o��T��7��n��p5d��f(\$�t�]�j��d9v
�ElR�h��$�ܥ��O����Y"hx�57�O���`�����.~N�!�;�2$z @�e�Y��?�X�K��b0���t�НV
}O���]�^+��{H�a�0�\l�WyJ��?�����}�vyH?�f6�����Ў�,�5da�s���]47�����8Yh���Rq�"$5���ۭ�� ������6=��7���㜘k�[��d˅�1���BT��/�<!�F����-t�w)�(cM|�n��gj��]~>����N4��a*�q��x2��������CXnG��l�X~ܠ�8��NE?,�xfn+�Etd��*�㋏d>��ڇk3��{H.4���W4����b���qG��詢:���m���O,f<�1 >\���bR}��uW~�Ԟ��Ċ2�����֙�k����`�x�}����x۲�DJ	,o�S�Z��) �-/�M>3T����(�]Q�rÇO"LCڧtk6Y$�Mv'�1�v�*�_�M������@�$��5ﲕM���Z�)��!�}5ρ��&[w�{(o���i�`X}��v��G֗Q�F`e�$RV!��V��R�I���Z���d��
y�8gr��7[?27�(�a�� �X�$��$�Jf���-h�����Xu� +�5�\�0�렩��ka⤨7h��/��c1��Ҷ(/j1ɻ���bU���t�j@A.h[lqnv���nc��#�Y@�� ��ԋ��Q�V�|;wJ�e��u���d�u��������(��%S�U��!����#�?��l^�W�)��8g����f�3`�$�.,����_�H<󵉨pڰ��r�0�l*��,�ič'������?�"+��Ult[��'"L���(�;XםZ�Zzߙ���KW"�(���:��%���+/��2햑7�܅p��x��	�/έygc�*��\/�l�x��cz����x��"�"�a�c$�I:)^�����RI�2��T�5����B��p�x��?s�~p��j�R
�XReɧ�0u��k3l��-w�����M�I�U�)��<��F��r�ɦ�z]��y�"q���r*���*/gu2��u�8{ܞ�X��3���}�YZٵ+�Pasc1"P��(�
��
e���@%dt{P��ў���z��i��7��qS�ϐ9����\10��d*�̗m���H��^�����ioA� �Q�Cr���~d�_[�u�Z�Py��.��ru�1w_�S�M	�J<D�=,!yr1����Ls*�����E�P�Vt��0��ad7�7���4���Ԉ4�G��J=���ˎ�j������2�"��W��Y?u���6L�Hs��d�E��}�åy��
�zG��.�׏Zm��FB�B/EHcJ7de�si�R�8CSKAƸt��f��0=I�t}M3u����)�yE �e#qܲ+�c�o=��`(ϳ����̄�Q�5�2ʈ
mlt�ޞ9��+�Z&-���Z�>N��ʪ^<A�׫�=aK�]��	:Ӳ ����j�w�WGV�䁕` �`Y̼"��p�Q����
*��u���HķV.������A��;>��ϱ��d}.���y��.V&Ĉ<���G�?G�d�6Z��`��{��14��E���X+^~�V��t :����A`2��$�BgT�׀�ч���HK�i�i�����*t���3�+�D����&�Ë�`�@Ѫ�b����9�#�/�U|��+r�èL�d�Z���EĬ��bR��F����;�Ǭ��k���J�8�j)�4\�*�Gfi ��rU8�Sk�����L�|6'���,Dc:<��,���s���+YJ���w,̿@̊!T�4U���p%9����4*(Ӛ�d�Rvu�k>�  :R����zn�4�Uۿ���W���e���k�Z*�e���`ܲ=yv/��F]81&Z��2U#"3]@���ק������