��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|/K�^!�� �Ϊ�I.F3�h�]D���� �1x�ϓ�k�K]b�ec���9�̑�2�۰�}EW��E�aǧ�b��S��+�/Aė �d��׫�~^^��y�4�4pjTK��~<OS[�EI|�ݾ�wi���tW3|��.�OXhU�3�\�_�7���N�k��W)�$Q�+������FU1���֣>�R������if��'2[ѳ�8A�y���<�Ѫ�7a�y�T!�㹐�o�?�u,�F�sPV�6��q|����Eq4? d�"�^	���W�m���m�^����Z�`(�ZY�;SCu.qM诞`�����&���5$��)�&��SD2d��"�2XWK b�,a���Ga}��ϗ�ٚ�Zu6�X
'*)xHH��A��Ot�� ��D�p/�FD�Öl���^�+���9(��6r��R�c�e,5ۋ/�����]q�PMQQ�k��S8�nM~� x*.�J�2tQ�l�j,��҃S���'Ru�!-�\~��6����.��ó�z� �s'S�F��:��5?����8�����J$�	�|/��r�>瓏¯�jp��E����S�]�ӣ�m��"�r�����]�%�p���}v#�$�%� E%A������y�̗�A�GY�H�G�~�22�a`�ߓ���K�C�v��u�����]��t'��v���HV�05�ӧ��z�Ac9��1���@?�)����6�Ю�Cm�xL<?p��O�&D�ȗ���k.�s�'mv=mg��x�H�_�������˼ӏ��I�]͞����p���{j<F+��\ϲ�^/�1�N���+�@=��tNe�3�,tbk��4<����k��k|��Kip#�t�SH;v�#hK�y���3A�>���u�4���7Tht.g:� � ֽ���k�7�?��;���H����g�p7���?�`��M�ʨ/�/Ewޥ��S�g1�h?�z�b���Kaæ�S�-d*=H�����ĺvJKn����K#I���-�E���J��>�f�z��D$\�_��dY}y�)M�&{0\Z��J�W�*���vJ���`.rD�wt�q*`�i�VSͣ�p>�������P��&{{������)
�?d��7J�Ⱥo�������a����j�	�H����2�	;���e<]JS5���!U�E�zx���@N���H����Zt���ѹ|�[f��>#����O��,�U�����p��d���/M���،��y�o�#ds;`H�#s�T���80g@�����a�n.ӟ��x���ao83���n���p)g��t�0k��CW�����(}R�6�#�;í)�4����՘Ȥi��z'H ݗC�'��d���qE'�M,|pwwEv����*8�@�y5nã	���
|����}wO [�R�!4��>��[������
h�O�<���d�Ɓ�z��� Q.ٱ$�R_JyVͩ-��s�J���\3u"��J�r�|<��9W*l1�����] (\R�]�-��d���=��6��g_���S��خ��5t����1���.�?�R�\�OJ�\P�hP\�}{ZX�;�8�+m)���۬.sPu�z��Ϯx�scsQ}�[��΅~12q� ��zL�K1�ヴ�v	C����,��)=��[?�ǉ���o�c�D�T�3��*���C��� 0�����}@Q#`�T�yiL��;��w�:�����s��᫹�:��q��Y7ȸ
��ͨ�»g^��3Tn\�����1z���!iEiE�������NhP�ڲOI�D�DJ3[����
���N�3��7&�:���X���*����%
F����~����h/��9���H��ZR"�:߻dۀ`^�q��SzY0^r6��Q�Q��_�?
��2Q���;*3��\ۄ�__o#O`��;���;����s��?��p����2��W9���BP]sp��0�*�����3�_�-�nl����q��p�P?�WǌeYkj�KiH��lM�߆�WC;���>.�o�ٻKo:�l�c�5�����D�i�t��.~W�����x>҂h�_�_��Ҥ]��q�8L/d��|fv�}fi��(an�m3���>�}E�ߒ���-�s3�u;~��0Y }G�����L��7R�����|ӥ��P����i����o�c�ܵ�I��1�pN����!(�5��e/wi�H�?��$��$��~��k t�\b�<q�^Ks�����FΆX+CW�Md�7p�%��
'�>@��g�7
��Ԫ}���J�>XЛ��{2���j"�i^.�l2^v��(�YN��)����v�.n�)��K��su� �Ĉ�1z*Cm����=;��dWB�}ZAl]��4�M�`O�\';.`�T	K��B���xs�JN���Y���7ؼ��63�t�D��Yĭ^�kU����x_���R+g�U8{�\q[�gwAv8;{�>JX)�7h;>i�0xތ�2q�ީ�#r>	8cj��_3y:R��;
(�
m�ϼ=��:����N�Zok�3j�.���(��Hu.��zsp~L%�:������T�c����s�!3��].�PB��Y����7N��H�ɢ����,��w���T��hH�{��W��D&������ե&����H�ɯϥ��;u����|�1S��d�7�o���MELYD�!�� ���e��kQ�����M؜�A��}ٹP��`�0T�϶ n�f� . G@3�y���(�'�٭����`���l�xU2m�������w���v��֍������烪о���ߩp{�~�]��N��'��������. L�a�_�3��ЮU�%E	��v\���Mm��`6���Q1�*����u���#���&�o��b�|M�X
�&!�z�+eN����Ҋ��'wS�=S���9n�����٠ȥ�n����#J��X�{`Yg��d;�.v循Q7�`\wd���S���^p�,B�.8�·~�_��t�ʼsZ�
~c��e���$��w���Y��`����МHpzC���T�㙺���I�}}���3.�_#��HX84L>�db<�[�;;ky��u��;��At�g1ܨ�GU�H��o+@���-��pƖ��(���|Z��sD�����80��$i�������������T�h�����SH��2QGb��8TK'QD�����Ϛ�eM�$4�GU��Ē�$�	E�$��&]��y錗��P�F�����?
d�ϟc��F�=û���ݏ��,D���`/z�_ڼ���Ge��RP�}]�o44ο%-��*X22�7�b�TJ�B�'�8�����#���2-�WN����J%�h��s]+������"����VRK�~�U��_��%�,��ȧ=]=�eTUC�l.��9�Y���p���|�~���}.�F�1�6��Mԃ�"�5�֖z����ʩT���9��F���1n���-���L��{lAj�hEXGo���5Ϻh]~g��X�y�K�0 H���4�P��C��]���W�w^���H���Ş	O�*EA�3���U��kt�K�@�!���;�����I��"���A���p�ex8+X<S��m�����~�2���D�˽FR�F<���W��T4� ַ�)r��ȶ�d���ni�	�h4�(pZ"�ez�^-�p<mVٽۋ�7
�X�x��|	K�� ;��t�âo���r�V�z�x���tB�&��pm�� �����Vl��@��=T��=����50He��8�n#�9���S�54
`1<K����|��A��ۜ!K#����qp�c!�s��t�v��o��_�]lu/�i˒-�j�"B'����� S i4rb<DOR��Zos>�Bm��7��7OG5Ƞ�j�|��s`L r�d�=�PP��À�p@.t7��y"�mn�¨�c<�!�;�a�T��7IH�Ŕ��N?�0�v�����e=�[�s���+w8Q��n;���s��j���hF.x�,�����~��Dg��~|���kn�����x�B�4
�p��e>��(�m�Y�pJAϛ;�n�M��j��6�C ��R���.�����ku|��c�k�n�{6�Z���.�r�ާ��iXL׸�3��8�@g��L��": �� ��H>�,��; f���Kb�Z�S֘�М궧41pe4B+w\I\U~{W�1��>0Q[�NJ�ѧ0�*�)5��,)�8sI�%�������n�H��z|�
�@�D,B����aݔ�3������gw�;Z��ﴲ��R�Շ��4.05�v�~as��E:kwLR	&}C�|9n�ܜ����ۋ6y>g�x���`���[F�YI�V�>(y�e�Z�zh�r7<G�­׮i�Υ���Gz]���j�*�|-��q��VpZt�b�~S��<�L��0�Ԡ&/p9��J�'�TŴ��Ѡg�z&49��I�Y�ZOu�D��%��*�p�q1~_7�����Zn�:L{F�Q�?�{��(\��#f ;�6.���^]���H�A�s�^�:Вꋳܡ��Nt�����!���8�>��rT���y;zV���a,��s��Ub�����M�T5�H) ����BF��P�fp@�8�zw�y{��<�%����FԪQ���M\y��hu����t��#��ɣ�^�/^�v�h`-�����8 @�վ5m��+���8I���݉t��U���� sֻAvW��_˴�č�"_�W%-���O�]�̾1_�R�J�j�`���^�M*	l�]�5�?K���9 ���F'��S��崳H���#="s@�������S��^��L��ܚ#�/�#
#n����S^j�?��U���*��Ȟ�? ~�
��t_d���Rs�'s��I[��m���~_[�	2�ӡ��	 �����]����Sm��\�΄N/�P�9��D��r&7$^�靇,���[ǥyg�<����Q���	�c� ԢNuU�}����&�swM����L��!,���#b�U�h�H�tV|�3�v�z�c��qK�/�B��O�)�J��@U�o*b6�ts�q �[6}d�9"�Ǉ��?�̯$�É���i�* �'���'�<|�u!`�W�V���ah�;�jNmve��A�З�Ӻ4�Z�łA:�a�9��'rv��?I��=���E\����Ob�fn�V$��N���׭�v7���Kii{;o<��	��Cs迤��ꩩ��+M�z���y�d�U�9�.�(A1��|���[�!X�{�)/ʵ���~̠�5�gu(��\�OzK�����{Ť��L�Kk ^O��@���W�<��8��d�pq�]�p��]O��e�`QJ�?���9W;|1�ۑ_k�Ld����Rs&ke���S�n�}۩�3w�K�W���Ɓ�"���P�wM&@��A�y-�l��08^1��\�~f��z��_�X���:��+<��R��^L�9�F���@��<U|~� ����·�rϨLK1�P����ŔiH����P�h���S�f��lw��m�����w�<�1��z�����D#��!Ǥ�bEOO��@�\�ok�i��W�_
��A�J��<�P�Ϟ�Wg���kʱAr��)u4Ĭ99�I���]���i���&l!��Q�QhP�1��O�r�y�7bA��l9/��.���A�#c�7;��ݚ��Iwm����Tl���c�w��61婧��C�:N��zi3�Y�{q
��>�1ֹ7�Cu����z���!t�'�$�����K{\��n]8a�w�	7�c��>��E/�c��QnS(8s�͗z��1Z-ƹ#/�
gܧ]��Mr��z�Ύ%���߶:QS�����&���Ep���N|A-��S7Y�=V���)2�J��#��k���&��xJ�6�H�9�H��<�Q�񺪏�0���鶾ߐ�~���=�Ϳ�.���#��5=���X4�i} '�h���~��hEm���Z;P��΀�gB\r5�z���@��[A�?���#��a��q�L���I�,���.vOV},�r��4�<G���n	����Ƞ�g0+��k����yTcp�KA�?�z&C�i0��}��:�6zپSgEe��@y�3%]�@�Ѷ�V�jW�3N�(9C4����Wa����R��RZ�R�3�(��eeY���_��ҹ�[�n��"��z˚�D�c����x �o7Ht_
���9&/o�ޜQ~D��R��$�`І�X������t(/*ve�ǩ�<(��ژ�ĸ�.�3��NG��ۂ<m٥�t�G������O��D#�����%�U�xA�T�ze^ik�����júb"�;���Eכ���Z����㴿�ɯQ�sD\<c���#��~gJN����(/�/cX�Og��(\��Q�uߋ��:*U�F�L�6,���ҠE���ů�)�[c���Qf�P6�~�_��o)�3&i�5�U7�y���p``���'W;�J�)#��>��T�A�#&�R�F�O���e��|o�O�`�*z5��yq��#'T�/�(ZLr��L<����h�*M �����p
H��a!�s9���$�٤���W�rӥ��
�ޑ��I�:�a�9���e���7��q[Ò1k�F=�3����4�bN�w>t2�#�#S�͉��"��I�|q .������qv�� ����y´�8��0TO1�#�r/�!ڊ�}(����NS^̶�p������@�L�*|8)��˞���~�d����ǭ��T*��Jh�E���jB���������g��$���n�bp�S�:滹�Nd�(N�Y��',��ڔD�C" ��j��3������6�q\�S���`,�Gr���!��҆TV	�p�#1�?�CYo.�?�ru�zG���T��'�	��a����9(o�K�+5�C�U!Q�!2������������e���U⛘P^݆��aZ�kn�+�	�(��M��<lE���J���\%&���1KM�h����YM�6l��)���J����@?U�/�&�3�aWP}R���ZJT�bc-?�K��3�~Big���x�Ll��T���������	�4 8�/�dF�c�%�
���̷y#1�(����)��ñ06� d�����T*���-��W�)#Rȱ]������]�<��hWi�esH$�r�1E�������d�I����)/�`�a�y����L5�������H^�9���ǭ2��YCp��3�Jy��ӤW=*!3C��;ٸ�����:�W3�