��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>hs�*�U��Q�����0<���ij5�f=���n��Ŭ�po����-��+J�j��7�0γ#~PF�Ç�n�~\ݥ�����I�'��nn��a���+iB�o�mp��O�C�HnO��H�bМ5<���\J;��r���:h�"0�z���7�=���Hs0���@B�[8 {�e�-w����;���C����=�\�<�f��4�E��}��sh�+�l�V��NB�6(G/����Z��k_�q0|�Rn.�-��?�9v��aPӼ�m�����)�\�ƶ)'ޭw��RSl�e�.��5���2���N�|�����B:�n�5��'Φ�P���s���v{�ӣ�9���D���ÖK�8���	lUhF�`�C6ێ,e�Jn�z���u�Oޞ6�s�~��+�ovۚ��ǒI�_'@����н��n�$oP��ǜvcM��;4T���c��
cL�M�̶�%�^��&���
A^�V����@{-�t�V�V��������^c���_�!�CHn��u0�3��;�I��N\30-�����R�~��8�[	�4؞ɢ��Ҋ<ML3�i���r�5�t��[�~�u|U�Ks[�2��������0�ŉJ7AV!�$�E�����;$qB�5$u�[���f��o��n1P�Dإ��S�X�L3.��h{G�s�r6b�Ն����`��$��������=7/�^o���|.ҙ�	��r���uw�t��_Yy�G�6s��E����
g�㡃v`��q^�����;�)	��\���W���d�'!�R���TjAo�쬂@aѷ
!��<��K�0�����ƒTiO�j.�jS�2�  ���3^���X�'@@9I�����l�݈0߽s��avT��Ʌ�u�t6N�]Qҧ���ףFٱx�.���W�P�!c�"�����[�E�&
��k�͡�</~l�H3�C��%�s��˭FYk΁�g�نضJc��D��K�:�B#!��
�&��E�8��ĩ+��B^؈N0��n��W``������M�Hj��<y.1t.Gj�TD9k��h_0ݹ�̑&��$M�@5�њ�� P�AF��� �n�]��7�dΞV)f-���$�V-��1}!���P7�޲3��z�v"a�R�J�}��I�����is3e���D#�d��������q��-�~@}��j��+�ꯞ!��#����.��Ӆ�$=�y���$��>���|qT��E���l���Ǜ�j}�mn�g��ȤĜ�.�/�{�q�4_G����~w�r�}���q��ͻƆ�X`�C�V��;�M�^�}�����@@p�g��	&�]�`x�����E�ٳ��ő_��3;�s���~�y�љ�*�������X[[8+k��-4�	�D�=,��x�ҵ�~#�ζ��Q���ܿQ��k�}s�q�<p���$7���s5pQWK�X8>������-�(XHerŖKLO	����o2�_������z!6Z��:�ߏ7���YNX����"�Υ1^�J�'�vmY*�)t-��.��F�K�Te����5�.�����������΂�%D+0i�l��X�a]�u0[@����}@F=�)K�Y�q!�\���٧��[�-��n����<t^@<aap��_��6�m��~��<�S|����\�2z͓�=�9��=�.s�Lؗy2��F��m�%W����
o��P@��<�zf���U(zT��;L�J�t_^�<��.*�b��2���y/!Z!�
��!6HDF��F�%��Jg:�ʞ�N�,�����Myw���F��d5f�@ո�8X?}���E��*��x�']�3�Y�4{6	��ub�!��6T�!hs6r;�����v��K���Ck�e����&C> 1���E�u禔��|W3��N���S
�M����6EZ�j��;)ٹ�t��Ę�B��%��ِ]xu�o�	T6��Iا8�=s�)��g��6�`&nB.$,Ej(�xw#����jh�-ʩ������k��-�9�_'�Y.�a	
dY����LدZe�d�hѷ��{`Z.b��'�>r�9�Et�=�HX���b�$�9эcT���m��:�Ou����<9�Yx�~�6�K�����C*^���4��(�>'D-��@epU��]�;L�*��X�CU�\�q��{�-�- =����џ�JN&�g��PG�*���!����Q]*L��]8qB;�l@��Xr$����vcFⅤ�v�׌���P'�st�����N`'%��3��(��޸��$t��#�+̠��&Œ�,�`0�p��A�#�!1Hu�ss��r��v����M�������*��}����3X��	e���'x�K���&�
���b0�>���:0'�<'�sW��65��m]o�,#��J��O�,y�aG'�z��v�X�ފ��O���W�r���ǀ��b>�����H��?��_j�R	��]Q*Oo��	�նx���{�l4G�Ψ���rdB5k7���i�����d��d�B/�����FP�h)2	�
���l�3H�j�x��9ǯ�����n��s�z`cò@Ų���&n�z�t�2*q�&�O�;@���ni&�1{P���2��t�PhF[���T��o�](�J~��;7��	���`ը�����;��r�ʦ���olj��_��:���,���uS��q�BP���ku9}��"����Q��<zLP�Yl�����梆�8��V]�!�	�p��u��Q�:Ga�R�oa!�K9�Ʌ�����^���8���CA�0E�ǥ�=Y�W!E i���<%6�N��[����2}/���w��	�@^IX���0���Cml�R�u��"7��Cp�-�9�uP�?��{MJ�2���1q���1��0�M\@<iop�g����ػ7�� 5��I��2!r�ㅮ3Ǣ�iv;3=�hTƴoQ(e�0��V�ba��Vݭ����}��MGeU.�Q�!����0n�~���	s�@���I�;���I5����MN�0��Ys�M�?H�~u'�~[&Z������p���Pハ�^�)0B��Bˡw�䍉k����Nq
A��|||tFz^�&S�B���O}w* 3ж8,�@�9]�(̻ �v��q5��v�R�TO;���/�4���������j�Vy_��f�?�F��i�6�&̰e!��C+�B��h��U`Z��<�0���2�k+^����g�ދ`s����VJL_�<�<���"�|��D�P6�<��C�D��D�a��4+�}y��U*0�%uk���  ůד����v���ddB���3N}C��
wU���S�������E������.��O���g�b�v l��Z �z$��t=cV�m]@N��%m���D��=y�X�8������n��D�κ+�IU���W�R�:$���4�2�8E3�kd���k�����Z��o6����ҽ0���~���psB����;��P "�#t��Z���=mVw�i�����,��R�)��4��>埨*E]�y  �x�
9._���s���\^̤���9�c  DE.��Ǣ֮�I&�Cx_|�I�`�h}gi���ծ��ū�dw	��h�O�������2���l��_�ʼ����T���[f��~�j'/5�(��ɤl�%I�b��$�#$z>9+��"y-�.H��/(C�@e�q�ELbmK^���3���'ċ���&;#�3�:��D����L4��V},��׬ays�	�p��0�&�U���~�mT3 _/�iR^�/wn���W%k
��k�J�-N�i�8�6��'�bd;�f���v�X���te��.K�ڄ#з��6���TC��N�� �y��)ǹq΀�§@��>����h�|]�����'���s��ћ1�Bd�v,��s�턋����n7]sR�5��
7�,l���:��C�x=[�Z��Ŀ�Ӣ���K���:	�6�	yS~�n-^(���n݉#ڤ���{ڙ#mI�Ѓ��+<��"'�Io�?�P��F�v"�:?Cx���R��ϓ�̨,+׾�zr�|]2ab=�2�Jmq�X��[5�Ϭ�<����'�a���H�ʨ�����S0����m���2K��[�Z���g�5���d�Ѓ�7R�x�}��?6�SV4��9Dv�T�{��F�CIZ�VLg��P�Zs#�c<�q|W�B]^�ˌm��#�j�U6Z��0~�B]���q�d���SC#Z�8����1y�l�r?o]�A�t	�	�aQ�[.��vqc�O���V������WTYbp�}��D�9a��+�lh]z9���R���+��vE�z�����(�a�?����!�pKdnk5߁b������H�k���K�Z/K���DҌ^J0�}`�է���������8=-xX滣4�Dv�C�Pp�S����dI=�pl��#�į$�cy��O��r#,�HZ�տ�Z��}�i'Z7z�CVz]�
��gΜ�}u9�5g�N0������pɱ��,���sI,�FN�"Kb	��|ܰ�\�?�8�&Z��҃nK�I�ۿ�,�5�J�&�5�ck&��/� ��_ ��l+ܐ�X�e�O�o� ��%����`v%in��:�Q��*��o�����!�DX~��V��U �r�A�ƣ��x�拏���-�1��g����ͧ�<�>����FVz\��LwN���d��#������Z�ч_��D��'�N��{�#��
�<��3��:�b�0�k�CW1�u��+2��ڂ1�W
`����8ԏ��դx���?&J<W{�Y�[�*QqY�uf��M�;�8��*�F5���`z8@|�J����l�ـc�'b rg�0���P��!��G�ɑ�C�9i̪�;��u��tЉE�v:m�婾��]b�^9ZQak�Q���c�	�OJ�|��d�zû�w(����>ZL�C\��N�-��t"�#q~�l\U���gI>�ާ�^N.Hh�3���H~�W��B�Oz��$A��$�y��hӍ,!EL^7�/SQ����s�����1��衼�-M2�bgw�}�n�˖���³��+��-̵«v�ҍJ�����U��pIv����7ԟO���IK[�p�=L���+��ٟ��Z�
)4:ĺ8D�����x�*�Vx��Sh�9u.�fl}S]���5��6^`XGs����Tk T#J��K�<"�Y���H�)�'��* /H���e�p�FΕ*��Z+�����2���$j���Q1P1�.��fi�݈�t�)G����B��vD.Ԟo���A)O�  >~ǛK�!DA��08��
2[o�O���B5R�)��uz��l[p�,R�>o?��9��<��(qx��:��S�T�dM�Np'p����fbh�.��<2�҉R��ߩ!s��Iě��13}́�������Pb���Z;�;��x�U7���ޚTD������8H�ttr�ƉSA5&��L�i��9ـ�<i[��Z"]]��ߔ �"���,�m,(���*&�����򺕓�0�=����5�}kI,�P6����M-�ld��ϝ���UI�l?����4�@�˞�=3��"Dȟa�f>�x���y��=���VL;��>@�5f�,��g1���7��?^p5�x�����d��v ���5� R�US!8)��~}�1��[ڿ�cm�@	;�RQq���š����֒��l��1���DF]�jP�������w����e��>4vWn�����j�F����V������+��ޖT��b��K�w�+ow�K5o�+�HH�����A�=�刺5�U#T?��n{��Z^Q="<E��t+�;���)��g��!�Z�ySH�Ѱ_��:�`�~Y+�U�!�É�B��iFƁfb 	$�,��]���e��: ��d�p�&�/�d_��%>���[[��A�����@Q7�P*�<�I��a�dq3�CMQT	�������fI�:��.�=�8�9��v�M�\��m41�K��U%P�~1Ҟ�P��>"	�����F5���\������d�~��S�\�rc���P�Fe�9g��+�=�4!@HF���H����3Yt���;��ߗS�&��=?[8�ի��7�;�UNA��������d�H���R����8Zn�	��d�v��;�(X%���a��T3g���#H-��I�[�H\&"@>@�jtˣ�jD�^�8�4�"�gd�$�yW��ȋ��6|z@2j�Yk��\���/�/~z�����Ҹ��a�e�C���)����byFH;��8�,�5��x̾=	��y�B�0Y��?�x��{��(�y�\^>�é���tWGZz�B	���5���;���s�<�0[�vhZ��ľ���&��ydg�����h����fՖ~�8���|p4S�b�?g���E3݊3��u��$�l�+gu�x{�\����TK~9����P�����6�$��@׾7hk͛��@`�(�����5�Zф�0�>�¦}����z��/i��?q%��~\	�>b �pk�L��$j
G��Ô�Bn-r���#",Yj�]취�Vy�H윀�C]:��D��^��X�g4f �k��!�)��y��)��ќR�-Q5�4h/�ƫ�ӗOO��s��?��2ޢ&իH=���جB�Q5�{.��3�L�U�.A�=�8;��Q�����Izi���7���x��^�FO�)��W.,S�j�=���OZ����o�2���S�~oj�6��Si [D���h^�}es"����Pf0�!�tP�.�P�!|B}���4{B{���� ��0��,ys��۾�OE�7�� ��@)uA)�"X�`��(:�尬Q�A��9��6οU�e��s�U9�����o�#�kL[�2{�
��M��wT�N!<'T� A�O��K�UQ�&HU����	=A:�Hn��U}P�|C�g6�yH�2�ʅ�.ɁO�t��*�O�{拐�P����Lh��/��i�`E{9�L7�-O�����A}N������!��3�B[���}�b9���{�,=T�X�Z/���X�ô�|}�Q7
D�{�J��r�v-ݦ<w}3���	zg���櫥
��$���X-���� ��r���Fx�_���U",?Ҥ�S�P�G�zG����n�	�H���J�Y�������f�3��	2��3z��f.j�1x�g�������S�`��jmo�J��aW��r���������;̥��1���( �E+���g�nl���	�_8�!�:Y��70���w�
�gxwi��H'4�}<@��'��Vt����:d:t���
:�y&��gox��-4��3���d)0�����#�)��:ٹ���ɺ.�{3;n�~�f��[��ه�F��BU�����+Fx�����/�b)�j	y�������i�Py�)��%��~V�X"��*��/�pY*����C�������B�'ܽl�3��8��8�"ni�������&5*�����ru�����J8���P������j�UboiݟV���\�/ڻ�?7)W�fh����@N��耏�����ʩ���r�X�$X��Ke�?����e-��KZ��C�qw�