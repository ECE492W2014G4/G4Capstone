��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P��v�"<ߞ��&'��k%P碶�R�ӣ�sĞ������FY&Ś���#��9�'D�m�c��}[�gG"�ෟ1td�.�-��(�EOdG�7�lU}/bn��JK�|�p<�	�F
D�!�u���s���H��Q����h�{T���`T~^��ʁ��E�fc��5�]��2gQ��n$�}����t2�Z�ο�XPw�p��GS3��ϡht�5���XQ�G-�����.���UךB@d��7R8�IPE���t�>�^.�u;�֬�����&�{��$|��r� y
�,����b�
F��OL��JA�Y�9��\)��+n��k�y����@$�ؕt����qFm��`Zm�j8��j��ŵ�E�_S|�Yʃ�)�	|�/��i9�t��Bzؤ�4HM�T�Ա���S�=:I�E|��@Lx����p���P��~�j�:��,���3x Jj��Uk�//v;�+�'@����mK��Y���S@��ڃ��MXY�l4������5K�I�Է��/k�ܻCz���.K����;z�<������<& *�� ��
,f��6��k�A���d�K�Z�bG���lx����O���T��(2���z���
O�Ɔ"���Y�#t�y����^u"7f�|"��v0,�x�\-�$`-�j�R��15�T�YU�5��3V�� �(Ӭtd�>W�l?RV7�w�)7a$��m^�Q�[��%��O�O;�l���gx�P�0I���T������[��[����I�8ɓ����A�Jm����_�����_9���p��97�:���*Q�<I����M#'`�&��{�.�D�K����E��ަ�� u���?!8,���)�u?'�]7{�?w<�� "�߶�YĩVǹu9��榩f����Y�zY�-@�ǭE���h��)���a쎨���V�OO�m[��v�h���FL�N��Aj�v��w�N����&�����͍�+*h���>SW�֖?�}�]��0���������L���i��M�� }�����m05�yŠ�R)6T�ʒL���m7Gz	�~�*���Z��b?��н������n2��G罎�7b��zF��O�x�{��¯���Q>�qp�UZ]�.���D�!� �5w��ωV�gY��)�cQ國o>V����l��'�E�i�a�'���+��9�ު~f�|���7��Q�(��l�t�����o�}c���nj�S�wu/aۣL��^a���9h��]��E�r�.}�wY�@�f��]	�Zr����%�a���{��K��Lz�P���s�i�GԷG����O8\~�K�wD���.����� �h���Qp�oOO_��':ƣJ���m+KS�1S��i�����:�M�.�������5��:��z?;��qyш�S�
#t`�Z�ȳh@�2�"�,�Y<��Dw]T���55H��Y_[����MH��r�m�l�5��iCYł�~�@8Vz
�~Չ���3^���H3P���g��f�Z�ΏU�B`�f0)l��ٜd�A�;�k��1���Dk/�ң�G8t蠄�Y�
Q�J�'<���B�a!�c辌`������ua7:�a�vM�C��?����"�M�j4Ko���t���;�������՞�j<���X{���]e��@0iaoW�9#�E�����<�4���V�䭴l��B0�Q�c��a�������VZYvl@��K[����g�ER���
��>F���ՙ8�=@k�
+B������𽺴�L
�7,�h`FA����]OA0�ì.��G9����`9��*���.r��`w�n�tjz�8�������l�{w��G���bD`tq�>XZ��\���	�?Sg�Zui�toQ�;��'E�M(g�]���L�B�p�j���`���gO0�W�m����:B�u>8ċ-Jk�;)Jh�������^(�]2:qͰGjYI�f>7�ޫ#�t��qsssa��j ϝ�Ě���m#�F%������H�E�.�s��i�xniZUÁj�K���
�k����f���'3I�C��
�'��͟	���^�U�!��PYMs�)�Ԧ˗]�o�;�x�i7[�͕5i�����]u\�w���&R��N9�`�r=s&���>���&+� V}�z�Qy�}���R\�"ያ�R�����b�ň&5���H&��іp5����ku?����a�k�ճb��ț��AA�O�sf?�=� 8���?L㤻H�� �/��@#��HW}�3��V�z���N�\K���R?������,0I/�.-Ab��-�ͤ䩩��|2��4���<q�����y8D�s���Yt��l#8��V�/�\�ނ_Nc�c4g�~��NZ�9\��Kf���\���3�\2���O�ɋÞ��9����ףH�w6W�-,2�^�:�eg��:b<�Y�8��������-�O�9A#7d�V۽\ڈo'׀��X��8�s��R�	!b���]1��,�|"�%if��n�.�K��1�����w	�௭ ��$�Z��Z��ȽV��"��,Cy�صBԳ]m�!{�b�C���es�Jfŧē��5s'|�E���X�>�X��Ʊ
/G���w�+;���(�l�����҆%���*0�̧��Cc�����}��:[%�J�c�0QEX�@�:'��b鼻Y�<���g���Ȕ�o-E������}4��B���6��C�#t�����7�F�-�n�R�;�D�����hҝ���X��V@�䠛E73�:�V=��s�KP��C
aY����n�"��0�u�<�\�?г�S��z����}ο���x�����������HB���Q.�#�=����}��!��85��ˆ��<p�n"A^�#�� �d����5)�i��p�b7�*��D�DqY�禥1W	���*��r��dV�w���KsoF^JE�d�o'�� ����v�ƻ&��p�5*�S��6V)��P��m=~�]�m\��G�;oI��2w�>O����e�����"<��҂%���>�����jr�E pjE�i>��y����wZW�L�_+��C���o�������I�� 8��[�� [��s��t�����r8݉NN##�#-�Xy���|N� �`�6�}��`�C�n-L�^>�KКr����En9J�X���S�����-lKq�%l�hϨ��wu����U=��,��l���+��5Z��|a���k�2�2G�j�ŷ6��BVJ�����ˍtN=
MJ�� ��9����R޹@��nX�:�%��u*� ��3��g	���Ͽy���r�H�����NU�ߔV��F��=�.�+ M�;C}B�q����3���ޏ ��o�1��Lт��jA�AV�I`8�Q�[i�w/Xj�4�#o��.WA%&�P+��w����材w3�9;�'bKR��)hx��,z6�Ì���
5huKO6cY&����"�+X��Q'��j�k"����]>����Z�X����v*,H7����*6�_Pi.�3oXSs�4ߒv5�m-�Rp[���*o���Y��{��d�����h���&�
$R}��.�臦��Лǟ��;�{A�w:��V`����C���.�M2)$�;��v)���ye�1�11 ��D�6��u|7R��-(�3Fqn�VaZ��3>Ut���o�v���02T�T�c=QW�*�zTj��2wė|U7��(j|ޭ$�>��8mg�΀����bs;��eAĬ2���G�ڗ!�a����3�`�]��E�!�M�0��gZ�텪8����u�=S,���H�W/x��{��8��~B��nU.�ȿCc�|�f�����ߥ;�~�	�PX��]Q���Ӯ�&<����Jͩ�,^2���AT��唃�=%�h��3�?�^���D4�(��?�����,�iC8��� �e�B����-�k�K�ɼ�c�/�H��)2Ay�XpfW�K�r��6|1��A&̷qB�i݉�
��r�I�_��O$=�!z��R��A;ql?�.�Z;�n^��_j�`�����5Ct�vn1�a*b��E�9�����Z�ށ�d��M�0��TX~�����u� ���UH.	Є��4RQMx��[1�@,�;�TXK���}V,`�Q��y�T���K2@�ԛ�6vu��G��^� L���i,C���"f���q|��9��eM��q!����<R�㭰���J���y_����Йhޓ�`�}�<�0��Iž�8��Oq�pZ�|��p>=�t�$5�\���Q/e9�,�f|�WVM�sD��lB>�=��a�n\�A�����J~��Ⱦǒ�4�m��lh9��;��[�Z��_��|}�������]�\�5
�?*y?6�2uf�E�;�!K�l�
HOKh��{�nD?�T�>W2��Z����+�ާ�0�����0m����Kj�Fc���%�~�f�Tʋ��4T�C��U�}b��l	�k�AVa	�8o�`���B����Z��^h
n�}�%��g��3q�����'Ѐ\4u+�Q�x��"�����)eѥ�U�B��}��u�a�o��C�S {��֮�Q=�&J���Q�_o����
 ���T�Y���2Gr۷c�xB>���u�i�Λ�3�D	5���0a��o${���.E�}�G
��V�+픰�Ѐ�Q�tky�������6KL:'H��y���[��3�lU%�.�SE�p2��Ei�u -� �"�YͰ�
Rn�ݾ2L�$���d�!�f��,�ҟn��&���8��7s+������Z�*Ҥcm|C�k׃�P�0$p��W;��Ph�v�����޹��ɠR�wAT��>��hy�0! E-�r� z����:��\TdnQ�f��ƪC	ą�7�L�㭚�&%]-�Ɵ�e'Y�I�/���T��x����5�P�pcTi����s�p{�[� J��Aa�VW���k׸I�������W<ٕm5Z+�L͉�
Oۦ�հ���[�>Uc���&����9��tţ��7�J�K�>��yF�f���3Q;������P��2\Y�f-U��B�Ϲ*����I÷�N�Sj4��VKC,�4����صasc~_�Ab9�2�E����8���g� EX�'-���E���1�#O��2\`Sy"���5�D���fK�j���.�<zd��"v�	t�m�<{�ۨ`�U@��W�Oo0!~qθ���9(�U�-zSr��ĸe��d=pZ�o�m���Q3��H		�� ٞ2C��zj��P�j}�;����eKO�3#��	E5��^ɛ�!XF��R?U��Tcl<�@a�x�Ǚ1�i�9Y��N��d:���A}����!�/r��M���M0�X� 6���o�Z��@�~�UWݲr��§��u�e���@��=�������{_�wGirߪ�l@<D'��+�{����F%�������g�wGM�g�`�q8���A�%�c��ɭ�A���x�<�~��:�le���~���I�Y!��p�Ad$�*Q�3?߰6��9ڒ	֑ �ت�G����/FR�#+B�rʒ�菪�L��j��|�D�G;$��ǐ��Od���Z��������������w��#��v ���8_�Pbju]E��W:Q��^�/����/�;�Q�����~��^E�2B�Nd?k�W>q�(�>�1�j�6t�d�Ъ�s/�y�X)��L����O��S{�,N'鍐���E��Jw/?|[��"8�D;����mB��H vc�)N^��-U��~Ap�԰Ж��գ� R�ӤH\�(���>��S�ȃ�;-����|� QH���b�)�V�����Ef�zh!�6	y�����!Dz��H�fʺfI'�ѫ�5�ksoZ���J1�m�\��?����9�ex���?��.���=�i�WbT�I��C\��B�#� �ފ����MW�1��8~���=�!�<"�cp�+�E��+3� ���ޤ14DZ�?Ö�S��T�,y����E��=��פh
J��-F�N�w~@l\��˕���Ҙ8�{�K�[<:��G��&��nyj�r��/�ý��E.��y���i�=��z��w�>P{-�$GUܡ�ԯn�N2`�T���Aۘ|��N�sZ�""���8b6�8+��(\����Q�Z��ll�ߴl�TQBC�(/_~_�k&�o�� @�D^ٙq�m|	K����c�������&��>��K5����ϯ�4ŕ#mJ���h� p�}ꊽG�+�`�`}�̎�����|�-�D#�B,�
��$�3����J��)Z���)���u���	W m��ԅ�F��o��4�	��I��M�b����
��|��pfT#B��2�[�/�d�Gy�'6.���lh؉٧=J2R/Z蜄�+�·��4S٨eO)��	ɏ�E}(:rEt���-T��"�+m�q5�n�sb�CO�b]�잃�T_� �#`/#3��P�#M�>Όw9-PaOuM��a$��eV�ȩ}��sh�ԅu7 ��L�IC���f�.�!�I!:�Tj���A�Np�;�<<��z������W�]�Lu:$�?�n%=��0�X0�	����	�8G��P��sF��ғՃ�/z����B��1cE[�熢ɉ��,�S	�s�O�k�JFl"����7i�fFO�V����q�2QQ�4nv���Ñ�p�*Դ_+!�`�='-:tj��s#X��+Ǭ��L6��W+6x�ZQP�M`eJqS	0Vz��f�_��8G�]�߃}�C���=��|k��8 Tb��=K[�{�ٸ�2@�{s[i��&M�j}�9���6�K���;�x� �5���8~$��~0uw9�����1�2�(���f�D�3�J�,�	o�ښo{�!�UH�⼄$�#��m����ĨL{�����I�k<-��7���~���;n:\�l�<�n��|K�te�R�/�\����Fm�W�l-D�1��;bg=c�O�c�����[�#1�J����A~+Ś�T:v����C��d�Ҹȕ��\L#�!�
 Jb��,�p�[���p�}b�wg�5$��YH�M�q�wXg�P�����C�u�#^�U'!�3�x7sM����##��c�W�.��|�x�1��do�3.�R��R��G�OбOT_E�p�݀t��Q`�u�-��^���o��fJ�jӯR�q�:��~�w�� �!j���"Û��@�-w����YH��	�E��0ÚG�o%5%�ɂ�@�IǄ�g c��ߦ�ׄ�R��v�?���W6�po��s���\�!dOVB�{&s�� H/���U��o��-��,�e��f� 隱�Aun:@W��xr?�����P��)��;�j�,Q���pz)�%Pň�}I��\"�[��}%P^1�f�Dw�w��,�)܍&�%ke@�X��\��[�q��b9X��{ =�3*ś��7�g0gֲ�����m�.� ���s���U�,�>lN7؜�;!�ˍ�^1P�H�x�3�L��+g���Y?��M�r��XP?�(�Av7�y߯��s�Ƞ9O[���͗�/�PW*����耘(ۢ!����\�qFO)ߕf+fԏ����	��J|�e�<VI3KF��Gm;��x[��l������j��5�/6����4}7�-�_=��+Q
ש�����s��ٚ%��<��zƄP#?Hn��G^��I6�-y���)V��
8��φ��h�ȡ�Ȇk)��+^�j3��E�pu�x	O>��C ���b؟��~ �N3t�{�#F��aȃS��m#��~{IŤ�ȡ��(nw} գZ�o���"3�lV��JT��yԑ�a��P̐��M���/���`Q���͕8���fD?1U��� �3�-�W���y_�Yq㰵^]vGa�����'D�	��K��R�3��7��,ta��<������d	�$q�Hvm�Y�S�X_��e�+̓�m�	��F�ۋ!֠�?�;J�]9õ1�����f�?�h�4���ݩ>S������|��Aٍ/M!1D�(�����$�o���3D�@MD_ �=6��#�uN�]�ǟ�ݜz��i�,��oc�g�F��o�
���NA-�O���E�S��]�9zM��B���]�Bki?4ʝ����s���+�����ƎN�W����X�=�[|<���ub�io�kk����*W	�o�u���cǟb���<G��e��������qZ=�-�#֌4Pn�4���Ǿ�`������g4P
f���L�d���
t���D̀��+ra:��)�X�z���l1\���Wה�����vO�4*��h�)ˮ4�!R\'���������w����ircF���z�Ӊ-NW���h�kܵ��$���H~�x��WT�4���aƝ�'<P��M<&MX�Ɲ�t�K8� �mN��)���궄wg��j�����K�9�}!^��)m�"���oxL��F��v�@ۛ�F`ezs�$VȄejxQ�@G�EZۋ%�O�[�w��~y�a���&�;|^��ؿc����L���)�R����w�z������J<�D��`	�>���D
�i�0J�`ճ��R&/}a��V�!�1[��&qD��T�eR����~����o�����N	��U<�����w�#�=Z����ZL̜��~���(����>�D��;k��5�nnF�ٚ��u��r�+:��Q��)���'M��[_߹��>vѸ毨������eф�;eےl��5���#Gy�X,��p9�VA�W��5c�Dִ=�X0Mŀ�[��ζbC�x�����<�ld���Bs�(�և�R����]"���r�+��WyҰ�����L����H�$r�R5�h�AP%Q���x=e�6:����Kā�r .��AV4(R��c��_ �)�N�������%U�j��[E��[4��;$��c�`B��~��ߥ3�����lԅ@�>�~WԈ�3�N���c=��ph�Pz�;��9*��;�q�ǵ~@��G�MrKo!�����=���8_%~LP�&f��;qH�k�����٤0݌�<��K���w
y��{�L��A1�ɵu����
W��:��&3nL}�u��Ǧ/��f���z�O�h�'d w�#L]hdϣ�x��cSU�fN���0�ыN���|.2p i�``�&��h���S�u��鲎��N� �V���Qָ$��%m�E5it � ���/U�nc����_�5�IߔUv�w�~��{�5� }��u[���1&
����g��O�hy�r#[n5A�<3Wn��Ή�x����`�8���k�L�Ʈ�� f�,��P%�<a�n�a�.<��,��`�����H��wO��o*�сWVo������$�R���:ר�_��8H���gQ�~�̵5j��Ϙ�b潀d<>_�F׭R�r|�M;H��{`���^:z��gm��Q��쉳,ԫk����m�������aiw�����x�v�}�������-+��:�8p���S�K]0R ��F�*D��̱�]b���̍)�4!���OG�0��Hw?���t;N��źm���7ڪv��쨨q������iIP�jO�_TuCX)�����o���(z�R^Pͣ�m���O��	����+�M�����kZ�	�k�z�m���PL�������{Z��5�T`�uٰ^6���}�o�'�[�l�6��"-.��c=5n7��*��	�-6��#9��k$��]v|�N:r��q8��h ���e��4�'�$Ҡ^�+u�%�mT<�D�G�44
`����<�U������uW�NL�e����:����(}�73�m0-��N���B�l���ɢ%�_c9�S�t�s|���Օn�DK<ͽ�����'��ԥ'���v�k9��[
��8�P��k'�����C�!��%\} �#�)@��مn��"V x_+zT��GT��X����,{��CN��G�7˚�!��Ѩ�R���B����iGp�$�[p��Qǥ�p�h�PX��m3���^���-��!r��H��j�����@^�e��b��Ġ#vx�Bx���j�7���=�������<V�d��
��sa���GO�u����<�д��q�I��]��;����������"s��j1{�?Y�w�z�f9�G��}ök��[D�u���N���u�J���>[���9�EZ��>!�3�PK������J��� ���~$4ʁ�j1�8�PA���'���K��a,�	2����c��<�F�x�*kv�zK}&oOј��z��ͧ�rQT�u�8�E{�vu?C�J<y�:�O�r��!�h\���i$����H�	*��Z#��g����.�U�8!�'�rOm��8�������k���W���3V�AN�Ȕ�S���m�>��?���8�"�&�
���zq΂N��Аʥ9�H-�4te3R�^�٢(��#��xUG;�2��RV�0�Eɲk<�'T�8�p`D����O�v(WL���N�t0����~3{GPA���S�D�[�l���B�|�#�/�CZ�,I|��S���W�\_!F$�$��8=R���k�Q���w0E�����x�K��^�.��lGV�D@�����ƕFw��
{['R��S��XP�֮f����+)��#)����0T^��&�<��S�3��E%���	z4���v�t�{mY<Xi9Xzr��ٓ[�Z<;¯�j��v�@cq�(I�@G�̴��w;�U�>Ȋ�]�Z��^>��oL|�ʥ��Z�`�e �(��g����wJ$�zog#��T=���K�O�;\��=oĊ���c��+�zٱ���<�=�UB܅짣�)��~�4n��H��
� ���1���P�(��."ϔA �qt6k�'4i_�e�Q�y?o��+Cb�z	Z�!����9�6,�j3'��Z�<��P�F��$ǲZ)����d;|x-I�V^����~��/��F�^��J�v�V|�FHV|�O���%0�/!�9UȲn��RuP��g��}1��ݨ#��\�W?ÞC��dd�iZ"������s��Hp�D�!��x�,�W�$k7i� ׷]�}R֧��+ mg���Cڏ�`��b�LG �Z2����^?J�2v�A#� j�(^y5�o|0"9�h)�hd1�HA���7�L rwG[Q����!��z~���#U�HQ��}k��B��G�����<���iv�xoo�T��go���EΨ�������G��;����*Zǵ�]�w(����J{wȉ��;ʇ6�fS�)��U�R�6�l�/��<i}�;��PNu�	�1�C�p���|U�'�K�̥R�iӜ¡�2��R�Y���I���fhR�'����.h&�{}���C�B'V�p�$�"<T�ٵu���W�t�߫H,�N��������DC���̍܆M���;� �m;�g5�K�x�ys���s6_� ;��l�����' c�Q�euf�~"��p ��t1�Ƚ�>w���cչ�`{L�M;�}�a��n��3�����ɰ�Sn�SG㚠G��
4~�a���qz_ �,��� 5T2���b%��m�@��.\qh/��e���c��0�K^tSu2��t����y�W� ���4p��.:�#2�KP�U��`\m�?�6e<BAr�T*+,6��NV�uz�������r�LB�4Ȫ���O�YFd�+y0��Ћ���P��*����ݛ�ߺ��x�h}�B	J�
�u�����|~�&3��o����He�j4MV�4�b�C{��T�W:g���R�t,�~����%`į4f旅^��s�j�J�'��ɀ�z�`��M�5�_�C�	<X0_D��a�t9�;��6����h�Z�8o�S g`�d���֕����Mu��?���wY�G�F�ߚ�e<]K}�fL?�U[F���[*q
e�øH�y��quH4��a׃�
��[q�i!��}� Np	�w��&6F�]�J�V5����+�(��C�%zs�|��I��Q��V�x���>��.µCL9.M|�1��p�W��m��?��ٮ�}FUr��.�ı��+���N����� wwQ�-8�ڛ�Bu��Oz<Ð��co����}pY�)�m2���S�j<|�3~WqF$�/n����nٺwj���Ȍ� S̰樛 m�"��J���u�|P�^���7K )�+�[�i{m �w�i{-�hU�0O�ea�,��}+oqz吧�R81\�^A��t'M�u!� \�'�d�1����0S�GS�p�.��B�xh�U%)�*�������=���pz�VW��,����d4� ��3�e:V�)���.����eK<.�:IcO	��y�Փ�VX��Ux������/a�;4,	y_�F~���ȉ�qȱ��H��t��o�LҧJN�P�i�@��w%����KÀ���cg"�6�7�I��E<�?>���g���:	��T7��'7|=~l�!�@w��P�s�%����m+WE����l���LiwK0p ��!����7)`�,N��.�]Wی��D$EՎ�6	�j�r�I�7��ձ�9�T�.�8K�>a��#�m����\��I���$���M������S{�4؜ Dv���� �H>�E���ÆFK�3_J�,�o�s������9>Z_jU\�ؙ$ �h��W骃��q%[��̆�C-���������-u}٪���sTQ��m磣!��-�y�м��A�L�)
�3EY��U=`7T�/�߸�:$��jߕ˓�����=*e��v����!臶�ru�ᄜ,�!wh�T�`��*͹�!s�n�+�ߢ��C��09���������K;l6k���~N�)��"=I����sm�b�%��"_��f�~V-��f�I�KSN�n)	nI@���R��'��jM!�%��tG;Ƥ�ی�"׫Q�W��:���L�$Ac���ψ�^l!�䛴W0��)�G���y��X��E��i�Q9��|iN��ޱ]�X�gd���,� k��.����B�ș�z�5ȝA��G���,�}��(rp~�T#��K�$J��~���Q촎�M���w7c���e��v��lq�m�Lʣ��U�A68�:ޣ����F0������Q¢���[�D�K𺮑�;qD��94%�Y�lM��W����^�q0��'��Y0��Yа�Y��J�˃	��58�.x,aeMI��2dK�g�#e.+���"\ߍC�?T���s�Bv[��wy�w�	�k�3R��@�f��[�G�=�-/3n��~������_%�?�� x�d�r�4�5T9�;_i��\Uj�]����	�H/�&n��.���8&ϼB�Ěk��/&�3�<Y�A�hp�?B�X��MMl"ܖ:�����?8@������͘�և�Σz����<�~�%g��)��0so�D� �&I%~K\y��ً�h��p;��a���7]+���!H;u������>^��,��3"��!W=����_ӤT��CPe�����?�{}�m�J�|V	���7.�<��\�^�8Hk�9�����i�Ո�U�I��4dwc��ka9���� �y��rs�GI��9h�xa��o�Y�ɂ6�fr���DZ6�w�S4N;�zs�k��I�o4�lr-�Ϣy�QOɒ�7��\ d�Yኡ]"���D�ק#���ߡ?��jVϔ~՚2��t!��h�.��Է0��>\�_�Y�M#c����ل˚��hѦ�z�u�y����}达�-�mnN,%ݤ��$��J;��6�a[�N��lI�o��I됻&��2l��i�o��=�|@P-+�ȖGP<q��כ�h�c{̕��䌭����F;��+xt�Z���y����-�n���*»ӳ�{�>c�E��D���5!��A��Y9��S�!��Բ̗�v����2=�I��G��"��ј�Z��6M��|)�z8�툻����Qd�K�_���NdBY���\�s���@$�I�׾�Q}��(j�]t���gH�-�#�r�4#�f�1�%�) �Vp=NW�Orx���ki��ka+ͭ���X&���K-됧����X�\+Fb]N
�����l��ڦ��a�Ӓ�ipw-�^0�O�>n��q���!y$�-���Dy�
���v��/�^]"���@�`�tj�B_>����bf+X��e&�������k��|x�����b,h:$� ���h0s��e���o���{0�X�i��\�ˏB�7�.@�YSG=�hIfF�p5���!-i2t�98@�޹�yh���_7���h�d[�j�ʐ�����t�_b����'�e��	����ynؼȌ���dXO���[�A֪<�M��*�U'��+;�x��Y��U
t����+���H5�#��)���wc�Cg�@7����6O����yi9O�X���4D��"vf}�A�k��t����*Y�pt��i8�X�Z�/��� #���[�ze�!�c��f�"��^	�7[ɂ��hXE�j�f�XY�}�gYW|�#�fկ��mz
��ٰ-��t��K�D���ܦ��e��O"��ʍqI8&R�/�5���4oڗG���N����j�B��Vz{�g:�]����XA�k��)��d�Ocj�G�K(�m@ �t4`�F����o����8����p*k�AM �I��#kP
ɿ�������d�������0q�֏�������6�!�=�$p��#��9���bm�)������I�ːYuU��o(�hd?�0%U%�|/�}���s>����*�arn���Ζg\�׸M��'�/�r����T���Ʊ���2����L
�B�ؤŕ�cN#tkR��wfD#�9J<^ �^%(�{Y��xf�~���"u���6����r�j�I�kY�.s�޲�0m�ʢ��	Ea��೭���H0�܀�Y�Ƈ��]G�Az����ݖ⻠�Y{
A��s��������y3w��M,�n���N�_���m�a��$�&a)"Zb����NnR��[�6A�o �Ne���9�1@�E�x_��G�N���*nM>�d&2a�����iǦ�o��7���M�*^)��*����m{
}O�M
�Ԧ8�pp���V�
xK����*��S��c�n�e&)�?fS�\��E�>�8$�����d=��{-K�-xf��K��Ճ����%�TP��{���8?��ѻ5�YO�^u:h�t�v�dR��i6�j�봐��s����r��C(�ˀ�#�˗Z=��M;�y��a�-��%`龭4�^}#{�[�+��G�8~m�B�H�q�Ea��a� ������3�%�֨��e�^ae��}�h
��y+BP�*�J%f`��(�[x1�����I���j���<��9SVg K'(&���;�4B�5-:�Q�F����&c� 
���h�)m�8��~�#\z�r�� ��	�M6N�T�� �A����Å�C�,����PҞN}���6~My���E/��Ϙ6��0�ԮW��U�B3�B8|e�p8�����4���bK[z�%+�D�ƍvcj�Bo��>fxq���1�/ȒM8J�pB��s�ņ�u!F1y��m:��f�9M���G5�5���?��Y�~'c�S�\�(8ثz�(�� )�������̢j�d�s� �q7��X�P�nO��mp�X�m�]2?��v(A&�؞�z�(��|/�H��_�۹�����lU��.b��N��7J�� 6�����K�����X�OH��񪜛����D��l���7��'����%�$�6�댆��
��fY`;Va:�e  �/� !~�Ffⱐ��ա�!��YUG�g����¹��>.���W��A�
��;j&k�ثq�s�!�$&�i�[rٜ2�*��w_��ԏ(��7��6�;Ȟ���Թ"��G��ùrքg���[�^�{�J`�����>���/�Iץ-@��`���6Կ�q���
��P�ؒ]��C��Ț&s�Pã����sD5�*��L��i�d���r_a_!P�C_�${���?[��ը��P5Ұ{d�+�AK� ��.O)Y��sr�(�1�oc$�� >�t�X»�8h�-P�P��n����Q)	2 �g�>vv-�h�$����Ǝd����$J�福��MJ��9�fL��� �Q
��Ϝ��ڰ�_�t�vq֕��Ch_:���
���h�S�w~Ya����%�MX:4}e(=W��$)��j�K�&RD� ` ��I� s�L!ܷk�<���q��mO�.��tf'mD}�@����b[�p_� r�E�����&��ʖ�$s�����y;6&q%�W��k�^��ij�]]�#�U��l���q���Ll�߱��d���V��^�g�j�i)B��G��ᓰop K,�]ԪA~�^�!��
eX�HrImn��r�?;%Kt$lw��n�ҙ�!�B���K M�����<�` �]Z�Me���I�d+i51�����aL'��
\������C�je�$��I���6k��2��v0�p�a�w8G �j/w��^�ϥ��)k��|�B0S-�I���[��z6��v5���m���� ��հ*��n�ɜX]�1v���.������,9�d5�_�|�x?# E�<,C��ḙ��n�É�E�9<$��8s����R��$��`�XI���j�0�/h�o��:���!���>�6@��W���ĨP�nӼx@�|9����������l�%]�m�hUߩ�9�2����@�-��0�TD�G�(�h8�wxR���j4�2:k)�����ث��(�Q��%z_��ϕh[���jV,�5�%�"jfP���b8?8@������	�R�T����m�jX�僯���3n��JQ"��N���z�1�2D����;���j�T���\�3�ګY���P�O�茮$���7Y�0H�_�Ĥ��K�-��:�5���I�;lT����m�2�b�D H��R�Øsjh_��l���+5A�$7R�6<���TR��!�9��K6_gV���pY�d���4*�%xô��5 &��cQZo>�;���TO��a��L9���t���Ё�W1���0IE\�#��-��WU����,�|>�K��S {�Ix�Q�! z������5҄�,����˶��*?-/:K)�~h��_��=E �c��ps�y
!�K�H ��u��9�������dS�Ƞֶc��
}
�p����Y�su�yCС4�(���C,��Pd�FHN�U��+���m�8 6���3J\�kWg����޸�'�Q=�En5��4�V��%��=��N`�)�t�F�[��K�7�o�M��Ç��0��Sk�@�q����Vz#�E��%�(t@�8ܡv�!����xj(��*����Tk�`U=��n��e�����8��
	�5�=�ꡳ���F>̧O��0����Wp��ӽf��� �b��0�3r�;��o�%/)g{�͍�V�'�ǔ���,�8�"c�cs�Uܜ�8�0�%y(8�E�'rN����D�;h�5�[R~�҃�g1�b�Ǌr@�z���5���8Ҋ�af�k�c�&�N�_kr�^���@/8c�-}ނ㱨2�ԙy���ޗ��B�5ƌ�����":��E>~k�-|��K$M3�&�����S���x\Q�/�X}!�J0���NL~3�K��օEg�g�&^={��ͬԏ-��.M%[ [�Q�Q����-��.I��B��~ho'e�ڱ�������d�)2��e:}�6����PK�C� %����|���K?��~j����ٛp/ P|@��q��Ѵs�u�W%�EW+z�=*:sq���|���|sq?~���d��奝N�s����e���{���3����U�-c_7��q�����&<IQnٗs��Rћ�-Z�F��e9;3�k�>%:�!4����]J���FX�1
>�\�/�C�0��ɓǱvq2�Q�'�o��M*%��Ǔ���n}a�ڴSn����$Vۆ	�`�`�03�b/}�����,�vV��f1<Z��%P!�'P��b �l�>,z�¹]Bk�1�:���f�S�����9LZb�
��#7�ٟ�P6�����\�~z7�z� Ӆ=�m��3�eBjal(��\��ŭ�K:A�	E"I?���79�ƥd~����Z��C�j Z�P�X#m���K�N�}���࡞��ן5�%��8�MI�ѩ�J��%���p�N����r:�}v�s5�ej�粡����L��Y��Ss���>�g�q`)��o��`IBd�<�lG�QJ�ؒ4��L�za�e1�=�Js�F(���k'ub^�ZG� r.�2˭��ie����u�`��o�(i�aR��&E��<��F_Q�����ۃE��}���l~����I4lQ��"�^M8�/(\xX��sj����.�įoY0�F��E�|ڭA����N_��A����� �+-�}�0��[��1r&u�lڹ����qߋ�LV��XCT+�ąt��)��B���"~[Ŕ㘛<��/�n5$u%������\��{�����	)᠋�:��%��F���yy���<H�Ekp"k�ke���?�:�E}W5�K�Y&ǲ/Rk���/��_�ǒ����5�ɰl�]T�.�Ƭ�<+=��� ��������MQ$ yf�����ҁ���,Zw���57�<���).��o� x���Y
v��z�v�;��%��+)����1~�_����&�Xp��M��H� ��B���o�+�
l;JTY{GZ�&9ϋ��*�/��P�^.���B`�e�'UXN��և�{P��\���-oEl�_�+�O:.!���S-�����)ML���Zӕ���K�'d����8�� ��	�CSS�'���mu��(��c��˼��;���Yܣ�=/�S���| q�f����NW�(9��MA����?��I�PՖ�,�]W�j�]|���l��x�Xj�sJȔ8�Lx���]���A��n��h5��Ҫ`:�y��WS�-��|O��PT�ݟc���Jڀb˅�@9E[W�P�9e#@aP�@93�f
���XJ�[�F3s�0|���D/m;��t�K	�O�����X^����M���rt0S&�J4:]5�B�Z������R%�K]�Z�����jJy���d��i�Q����t�^g�\��j�̐�?��m�84�*���S��z��р�LN<<�vQ���x�G�I+���x��*U�Sx�_t9D^w���6�����eUj=���N��wGs����\��-���:eMk�W�z�^�q>�>�g���6��(�wU�+ �����[3�9�����ϖ��@O$�J<��kGU���tS[	�^iC�k�%l$�w����`�f�1	�kOl�&�=x�6���;�KBwH��"=�"����{�_.?��
{C�w=�E�},B�rD^p2�0N)�� g�#�����9Z���͜SJ�*��l+�	
��)�ppt@�\rD`������E0����;�av��wo\\_T8i��>e(�
��A��Oڲ�»��)޴&E�n��r椃;��e�I�U0p�=(FmkJ<3��
2�}�oD9L�f�$��2�n[�=�x\��W!ޅ���<VKjF�
��{��,��;+���M x�����J��j�Bnj���ޠPlC�cD텻�7�߶م!)���a!��R<;�Z�K{D��Q	���g3t�^�"�ֽ��B��1J�T[=0qԼ*��4f�Ev� jY姮ĩ��?��)��E��>j�ۘI��8@pZ|�}X5��tbr*,5~L���r����jW�b")8;�����"�;X]�����BJ-��������2����|j`ţ�C�,=6'������$1������;���)���?��&��j�6A���QY�u���KOhGRVwadQ!]�R-?�������e�Mw� ��b���	E�������p�l��i��J?���p�-ܢ9ܺV�� $���Z�"���j��TCV��,�J�M�IuY��_�н�7 Y�G�kp��,�n�i?�����,:�i��b�GW�(��z.����7� �
F�ٳJ6ܔ?����(/=l�ik@�	����@�-rƿ�|� .�r�p��-��a�擷7ӊچxN��!t!]����Q9�c� @H$�^[��b�����xCGh�����!_RGk��<Z"�4/�W�#s��X!�v���Eʇ\�Bx�-M�Iϫ[�fΆ�P��=t8��c
d�A���DnҢh	�zQ%�g���� r}�,z59p�s�6���G��1���2N��-�"�X��jY�㙕���-��q��Mu�9�g�;eQ:J����_~���>z$O�=Jw�nLj��0���]o� �� t�Ԉ/��^���x�<����V�F�!��B� �'ɽ\ R�~��ӹ�@cf�7#*L���V$1%�����:�����5�ؒ��R��ح��E���(�8�����R���{6?!{����6�jCOE� ��n�r�a��O��:�����8�Y[�x�%7��<H����Jn@RvVN�v?v�C<�y���fzN�*�b|&�3(�_S�>����V��I�=��g@�:0!�^�̎ʑօ��vH��R���Hm}^/��Oݩ�r�	pt݀��B�j�n{-�z�[��T7X�)��������*n?�؝��TޫxHr��.}�$�����a
��z��6J��&�zj��Rnm),ӥRJd�V�ji���Ru23(�����qQ��
���e$�wv�Ui�K���U�{�WZ���KTT#:��p�	���)�,5�¥Jp:iʠ�	NS�0�St��:��̒�aˁT�;7ʟn��}74B6@@G˿�zI(��=�pU 3��`g3zK0!g�}���bB�Q1�5����?[*�=�>����GA��y�zsF��4te���M8��EG�P�lY���W�GGÆ8���c�u�4�K G�刹k��ɓ[ȌW�$T%IF�1�VcMO�'�:2�~y T5���%I��@O1B��m�5AWC�Fx��1%�� O��F��b=V=?�/@Ҵ�W��
p����{Z�^�쿯\���E(��W=�jZ!�V��I�hؗ���5>����SR\:�A��>]�q&�:Y�h:�1�Jlfu�O��r7�?&�����\*X�������3Ee�!���&����w�3â�Q=zq��� ����(��ʵ[9�����d`�6�8\<#Z�E�;_2��;ƬE������E�ƴ���܇J~fV�/��b�d5��{�������wm�T�[��1mK}�ν'XhF���_Ì�<�d���G�A��	Lͳ�S$9C>@r.i���l4�����W;u�ɴbi��������)�G�.�̭���Q����w���>�q�l��S|�j��o����m�:Bn2�t-��J!]O�^�Agn0��wC�`t��^�s�%��CiNc��"���l��9R6Q�+�N\��0�����	(To{K�V<bUS)%�D�ѵ�/h���^�i��sr��"syqؗ�5�Q
W
Bp������Dry9^��L��]L�!�KJ�"~d�\H����4�����G��"-��&=���X��;�^���&����@9g�o��#��!q�'��|�lO�v�j_M?�̢�`�_�]T,hJ�8p�F���֡4�01Y��[׻�`uw�c']��+(��Tpyyt������m�
��� T-4{ T��jg��'�r?����kYH�
pg��n�ϑU�?_j�3���T�B.rLdw���d��3`�yx+�c[�����a�k�M/���Uǭ�n�q����#R��D$��M�
�?<�6ݵ>���Z�f�nY˱'����\�Q*��z�#�z�j���V!�%?�q��%��PA����{k;�k��Zn���ÏL�.��������=�Z�:�@����9��l5����^Z�侜���]\.�|("x����<?��	��2�ZK�ߙ�r�y~J!3��t��Wc�	D��8��+mc���5�y�%CK�ߤ�y�u-��vO"��꾊�)��1��Bu2���4}  �t�*�Ŀ1]��z�5M<��Y��_����, �$��En��q4uN�A�Y����&}^祪�vU��%F؄TP9`;Q��2���Ѵ����-
,{}��+J�Vu�3�ƨ���][��dO��'��Y��a�:�Zeɇ������u3��	���-�C���"v��z�����E.�\)�ajh�ӳ�d����%�mRoH�� �o�J�ɥ�E����p��,����WF��d��Ĝ7W�>�v2yj����{�R�r/V�5�Յ�}���[[��ps��
B�{]������^���Y��}6�B �x�
'�i<������0�K���e�Ղ,��?� ��D�}�˝͇���N*�"�`9�}zb��S#Z�3������Tf��B璮:�[���Ŗ~Q�ʁX�ֱÊ�\S����P�y�A=96$��~6HRl�7��d�/�YѺ�F���Ӹg��"U����!�5��+�.��e�G�1�y1j�GL��HJ%Ȑ�(Csc3Gqt�7ʹ퉩}�0��(��S�:�~W��vw�i���p) ��x�A� �(�M��܃�[t���١.^���Wh����CQ"U�r�ME�V�A�8x���S Y���/}��-@˔$-�;;g��Q.���,�1��P��>�]#�"|�A,Y�?W�9�ա~������@��ꉾZ'��q������ކt �W)�DQ� �;b�7��!|0}���G�+��L��e]M�3��~fK����.��ao)�7���ޔ����]\��|˫h�aq���5>(��,^�'8X�Ť0G�.M:���c4h8om��I�_�"���*v�a�OM8HV�O�R�6JQ7e�T�i����?!O�H�DY'�~�;���ʾ��>�*㸅=��zI"�G��~�Y	��=�J����BONך��+OG�V4�>�'^Y#�钕�/.V� ��@�d��1�9����@�m�%w(��Sz&|�	�1�!�l�	�KX���,��z��4�(W5�^�~��D	d<���!I}��|�����	� -u\C�S�G�Q�$O��WK0*^�F��@�<������zݥT4�U&3��BF+kC��y����ag%�R �P3HŻ���K�	����ܤysK�M>�79:/'%K�6q�����#���t%֑I���ѭM�4|�םZ�+�#ɔ�I=����gyl?5aG��!C�r#��_ˆ�|��p!�<���|�)�&�06B�͙O�G^3����Z���qn�{�s��������m�?���}�Zo�=>�}�[��e�/�!��Z.�<�6�>8��R���3)��@�='����02�Dlx\���m?0�򬜳�X�_�&�=@Of��sۦM����p�Z�4J�T]KB�I �m�m:A��Z����	��V2�ez+��P���
q��ܮ��&G��W��Qn�DS.�C�q$��C�G+@���6^���^_���(ʮۯ��pTD8��t��֐j���u��� {	⺠\ƇW��=N�T%�$����I��l��bת�(Mi2�����3݅8NwL3��p�j�(���b�f�<v����zԠI�����h	�����s��ftXբ�
���E�:2�6=d��X�V���U f�}���
U�eD`9T{����`���\$�3�*ԯS�FgQ��VqTܹ���]@��j��w�t����	�-�ῶz�Y ��Cz9זJ�xg36��_��� j�!�M9PN���-����!?B��fa����X�� 1��g��ULU��22'wl�-Q�f������T@�r��}����c��E��Z逈LPګ��l�
o�mz�����k�H��.1���Yv �tݚ�@�Z���h-e��~Fe� �X�>�nǱآ)��U�d�V����R�X+^^@~��oGHAc
zc���e�_��*�Q�[��f̶���؄�R��[@�+�&j���d�����׬"���s����ɐ�&�<ы��*�P�╤�xS�x(嗝�@�����D��l�F�#��zHԴ˝��͔�{�>x�}�����$��eVL^Gy��F�!�_h5=�$�j\��Xa<���<鳷q�^*��M��vL���V��8.��@�{ȼ|{q1�)�L�)S��Wo��ySij�>Щ"׋��YtV��ia{���+�>�V�;��p�c�d���^��=�~@o�_�L�q�ZWb��n�5�!b�5 �#�S��|��Iu<h
�R��r,�C���r�IE�0:�vXm#��'���m0ɿ�a�qY�����p��c2�����9Z���E��o��9�\g�#���C۸�E���ت���P��n^֮�MEH/n�-��$�a�ĥwݦZ̼P�N��84ڼ�2Z���?U|��)��-��"l���B���cj��YB���j�B���=b\�^"����!��_bu�D0�P�����e� �`3�kgߑ`菬�)ZCY�(`�P�L�
����p�ʲ(���i4l��
������ѫ	�Ԋ*
���8 ���ԩ�pA4�g��yꄳZ`(��lC3ݱeo����RM#��[��LI�R���^W;�I��^��H�w+�z�ǏrG+�r5� ۫�"0zXŅ@'�Kp��_"'"ɜV�L�R�֛N{T�#sl�[����6$I\�%�^挀{�BiVQ�\�o<�W4I�`pz�_�=i�U�KK�Ŀ��pu�*�����CS���8�V��t2��ת���%P���]��E��;Q��I�ǒ	�0�����[j��K�P�n��H�oxv�r,��'7.f<F�@�^��ܑ��Ui�0k��є�mI�\�J����u'Y�H�<�V��Lc�׉HR�����q?N!���$/���R[���KSZ�I�9��`�`�Z��Y�w%k�#"ఒ`�i����A�ż �FZ�Ǻ%k�W�Vj��W�6��ƶ%����i�e=��W{e��7,[���+�P�+!�(Q��L�Vט�i[���qO;]��G��ǭ�V�0P�+�D�v����'55�&�mR6>DѴ��`���`��rk�W���r�_����߀�'��6ɳ�=�}or��f��.�H�����?�o�j��=.2�ߊ�G�;�������%�텺���9wkP�4�����G59�f�>l�>��>��G�G�ox*��F�P��߲O\����v���ۙ��"��E6�Iߠ�O���m��|f�LG�@B�䊴9`�Nݣ-2��Oo�iWI>�t�a-�k��m0U�� xn�(�V���W�
���Aו���1�f�v=������)�y��e����;�k��+�+t�o-#�S�N���}pvlC߶_�=;x�uF�f�J��P�&c�_A(�P�FsE�R#�mvKq�������_���"�<���6�D���u+3APGwf2r<�j�@j��h\�p�i �&1�^h`��PQQ�DpW��'�O�60���Ҷ�ڝ�Ur󆸿�zg�=�}d!�o��n�HJ%L��;�H�2B��BR�KƇ������� ���b�i��~"i�0lE3uP�Ke{d��A^T�Y:�' r��]�wVx�*����aZ:�XO1�sz�^��Ϡ�Vz��xm�Ԑ<�#�W�%K�j���ze�3��u5+͠*��q�q(�ƫJO1��a�u\3���	?�,�${������¡CA5���bV��&��5oyRda%_`A��h$�ڟ��v�Ju��~��WOx��T�ۓɌ�b���h2H;y���t)����5�߿���^���݇�Y3V�f|�1�E����IN��.e��o@�p���B�5m�LH[����r���"�6�o@|���
!e�m�6��[W(μŘ�������Y_�����<�3t�
�4�j�auc����)[�y�X�����H4C��� �`�'#��!�#��b�=2+�ZP������Wg�t8KfVR|�-P���^�N���Ŏ����K��VzR'����0���o�3�<1�����'TP#�!		�W��`�|���N^݂[x�O�����m4�)$�Ψ͒u�5)�6��|�����kS,o/z4�h�d�ȐC��e!������`c��L��]�ݞL0էj` �U�돉)�+�Q��6�+A�H��,��NMt��}] 1e���	s?�h��ۡ�\SB��L��)C�N���ԭ�[�3\�D�?���==(rVQa=jj ��+��̣�I�#߲��k���:/�dtY�I�r�>��n��a���L_����}�4�W�e��
ۚܜ��}��H��),`2�&�M/�7�J)���V�y<���0t]�����E�`�0��ń�:c��vxT�1Ϛ�@�V�7�ŏ=A>�>��� �4$�X�ߦ&�az)$�/4��ҭ�IƱ�wd�(F1;^.��}Yg�/��L��gz�H�>�񐴑{�?buM����FUPO���ن���G"���]!�P:j8G� ��\���Odxݱ�Mf��fU��e�-5�7�tB~8[jFC�J��Q�G�WH�g�wh\S�[�.���K��<E����A���J�����| e��>?���:D{3�T�����LH�:���ڕ���-��
��{0#M-Eê��꤃�}m/兝m.�H��+d<���,��*����ĩ��y澲(x�[��rǇ�n�O�ܱ���]��|�a�h��@kKT�ˡ7��dF���Xc�9�� 4-ĂR�ϗ����"Ȳ���N��!�6 �J$_2:����8��Q3z�1{��J\.��ql�,�}�R0]]�O��3�(̭#97*�T�%��wR��^uBBy�6��o�kiۂ�VKe�Ⱦ.�
����/@�����t��=�=����i����=T�q='���~̖H���ߒ�A��Q��$|�\⃺V����8Y=@s9zo�O?�n8�O��Sd2�*���>�Z�94��>ˊ 2��,b����$V��V����a��̈�BIN���o��P3��g�z��hԞ��&�f�;z ��Gm�*���)[������o�(����	�VS�(�S��~�gʳWC���uR��v��H��x����_]�Dԅ�u�����n#���;(����A��{ad�,��tj��UBa˫��G�� Vj,�Q�4���+��*5�K��pƞu�EU
�@g���s?�g�2�b�^<�1�;�VV�T]_iј��F^!��q��>n��Do^/���eP�~��|�Y�F��ȶXǗ����sQ�+�f�WN�Ĩ��`�\A�9+�gu4��~�s�W��1�,�,�tJ,5_���E|���+�U��a�R�"+/�*x�r�4�L�CkOjΒr�*�����\�3i��'��Ly�
�3d1�8��臂BA��A����,�������2ڳ�$��q9�%vk۱�-o�Lۚ	j�A�	5(�V�/gsՈ�Ӹs�\�D�.Q�^F� ����u ��(�4��gWl%��O<aJ���Aa�:��G@�Kop���~�M��x��S��02����]�<�}��������g��Ώ�ԑML��A�uFax	I��[�a�2�x�k�v+�N⥧����fq4~��������#&�\\�[���G��#>����g����U��8�kI^Vg����Zs�Q�S}�ۊ�&cG�N/���W	��s�O�'7��7:��]ީ�k}�I(���8��	�� �7B���]���V�%1h�p��AJh=���st]!��^sPM%�FV#_����5(%l��l�)}��*"�	n%J*H���7�\qĞc��+�6�%���{w]Gd�䏈;s��=P�43��X[j!�$��.c��U����n�D晲N������1�E���V͈/ G��(����I�P)�m떷jI��Ϥ~����4����\������~�(�b�Q"�4���^�p��	3P�A���ƛL�vr�J�<c��T;�"eb6�܏4���:y��С������b�!6B�[�>j�a�.���aMq��9�f{h�AV`z��+Է�\�D=���M�$�+^B�1s�^-,�Z��<Љ8r'Q�;��p�Э�^i�T(K�VD7F�F䭷��T�P'��/ou0���YkH�Yּ�o5Cq���Ñ���EW�Dl;%>�n�1�4�a�.KDѾ��~;���E��A������me>-|cE�*K��"q��s/�0:���e$B��%�&�Vle�xN�k	ʼ��TY�ʳ9dN/�hG%���r�����i����O�� Qءe4��3���[$�q��� =k�)v�Zuׂkq��Xȱ&R��?kE���k.h�G��b������:�0��DE6`�*�o$A>1�h�8�t��������hGj��"�l�XiL�|�)(��y{:��qI�ٯt�6@��g;|<bќ��Q��]Hà�l�L�B��d��0i4g�A�<�H+��UK�BJ�r
�ps
�[���=ґud�IT���ߍ.�B��(fpgHS���ց�K5��%��������2�mL d>979�����Ħ�%&�^��d�2�HZ����{�h��&g[f�}%�B!�M���@�꿾�[��2��`pt��u���uO>y	j[��Bi�*��VA������
�|��,�GhNҦ�I�au��Ta\�T��	�萻T t>/xR]�=t~{/*ߋsip:�[ ֆ������(C�x ̳|E�A��(o��ȴ��o�aEĂy�w��&�Myr��n^�T�6뚫�9��$���Z�`L� �dq(X�u<qk�(+I`�U���:7��=_a+=�& �ՙ�c=�8>jq�F}3��̋$�^J��Q?����{rJ:$cq�{���U1S���\�:w&���|J�����e�-𮉱���=x�A��=��3��?���G�GJ�m(������'��1x�d�=�z_D>����!�L:���<5Ɋ�ƾ�t�!��:��~��'�o���ŵM?�(r�N��Q�����@��3V�A�
ۻd�ouz�Y��8��q7��b��K��
@Y~hݩ��&[1YЅ��yXi�p�{k�\��Au���q�za-jF��&e�wOr_�Lz8�ٰ�b����C_90d�3�״J�~���'�ta���@5`��QIH��sބ_l��m������I,��W�r7��������|������3��@m�9�G��	�$�&��H�B,����dơB"$b(O�Ŵ������frC�c��K+�0��b:Nf��'����V�����B`��P�;��"���N�O��>�W<�/��P`EP��L!��"��sn�&�
��yr�/�y���Ce���-���+�S,��w(�G��欌��#��j!�*l�
a&&@��ҏHy�����_��`L���aVA=�:����CQ !��4H�l������0/d�4��JR�Q=��	��ѯ�����*6��]���^	�bR�K+"�ɟ��AzP���2�2q]��y�A��4����V��Ǵ��.�L)�.OzP ���4�b���O�õ��H��v�����K�Q�6��=�j���+7�w��v��^�X�Jڋi�����ЩF���9R���j���2���v�i�ym��w��q��.#���g��Et9�o�-�E�7G��憎c�yo%����R���� ��x�K�#AV�p�3GY���~��7����_Fo}���
Viv����2�[�s����f�M>/]4ȇ`�x n�>���w��.T?π�n��vZZ�r���0U��L��U{c�~�˕4�CQL�}# ~З�K��1ի�[2!4w��D��n�np�Iːx��O�n�+�5
]�������2�VFn���+�@�R�Լ���8oO��)]8�%M�b�MAI.�J�d�{XS����e���� �1����B��oeE��R�G�@62f6֡{�^�/hz��><{��g ��o��9�O�G̐���fU{;�N<|Kƣ&[s���)w�f�T����,�[U#W��Xu${	����wm�w_*�S��Ac&�!���5�!�G׎m����u0����n'�� h_�QoIK���N����p�c��jH�j 8,����[�&��J��mYU�J07~� `e+V�r_k;����	U ���^���H IQ�T��T]����^�F4?��!.�����Adz�7>spv#	��� �/Qҩb��R����ɣ�D�j����	�0+�Y)y}�F���z�7~�>`��������&�yX��KH�����7���������ގ�e4Tku��g��+���&��F@�4꘹5����*�9s��8��~h����~��=|�CF�Ճ=��v�����>��D�\��y�L:<��\�?7�{Duc8zP�D�9�'ۯ����0�����R�#s���)��%��%����� meqn��fM����0z���MRT�Gq�r��/Y��D��*H�i��si`"}*|�vT[�������Q������E���[��HqTg\İ����;�jw�:�*A�a,6p|F1��~��w��&A,8Po�k��б�h���zGI|�E�$��aPRV���&�]��J�����:-ewf�$��n���V��$n�T/��}ڌ���D����A�<q�0
�����[l]n���ݭ���a�2n��Q;��J��*���}�)��(��w���}'�D1�E����k0����ق��"�ߧ��>�ןD]����8Md��Q���È�izWy���~H�$l�ɷ������� �q9%*�����xW:v�����MI��\�0݁5�Ϝ�:���Xĳ�*���	�_q����3���/3c�B�.�Xc���\�␩S@'~���"�����<���1�w��GT�%(�a^#��Eԇ����Y0E�K6(=�䃞mR-T���<Ҽ�_;Rok��٥������1e�HY��KJ�1�0��Bq+�b�B[��>�]�q~��i�cB%���G��]��]Яn�Oz�5\~���WW� ��B���0�'p��`d�)q#D���M�f`�6�j�*�E	�lة暑���'}�z��v  ���/!'��%�{��-�lϨ�,@�����EN�u��:H��)+��j/�<�l�������Ue�����_�3D<�I�ڧ۷و�:���U�X�� �|�2��]&4�+3_���ӷ1XonYF�^nt��o}��;�p�{=-]r}�`��L���G,/�p1ux��ܝ �.��l���q�8��CoXj:�5U�9�$m�4�Ƌ=ހ'�D|���~�H�_������!�O�.�iB�&���dF�ޥ�-�8"2S��qO�G(�'��o��c�X���3�XT�������������煣'PR�����CaWa%=R�~�8�|b����64�*������Z2��2�9��<ܽ�LF�6�J����� ̷8��������:r���j{EQo���v�c�)S�Y�z��%�j9y�� d�G#矛z}���J�3���.F�����`��S�J�
�p�q�������썱�OU���ŗ������c�]u#��"���ÿ-��Q��E��,���.���]'_|�.�Ĕ6"�ܦt&L�]|p&Z��!�>ڠ<�_���6ĉ��v|������XKD8������oy�z}�|��ƪڹ���>[��n�ޞ�׭䤕�q#*!Z)����~=χ���ݡ:��6�󬯮<K�gm$�x�("TQ8�y�^ �U;�厪a�ʹHtKs�]%^E������Y�}��8TT<
�ɞ��)�H�I\VQ���/���sX疌>͂Κ�,Y���S����W/|����r�A��
�i��X�	S��Gx�-[ڭ���O���ˊ�t���Bb?�B�4n�К�_ր__�������QTa{' ��yA{i?� 9Q�9��v�@�.)w���)�^�����aX݌�JN�K)���V��[?�v`��#8uV���X����"p"\.�x���FR���� &F4ξ\3*ak�����J�����V���Y�'`������s��Նh4�މ&���?���J� A��A�
�15Lr���"����hl���jJ��uf�x�@�L�A�����Q�Ck`�o��*�W
S�f��9�������:�9�G���a�)Sjfi'�3?>����e��.��r���24�`P�HI%)d��4�W#ꋛ��D]т�c"J.���r���D@z��(rR�����,�[D��޹�_�	^�Q�P�C���7o4]_�����.�$~3ڙk�md/�R�V�����)�߿sU����r�Ef�S޴��^P]?%{vE�
��������&�;'��o}=�6i2&�)����g2X7b	`�5��u:1_(�q�,�� ���~	���`��ds��]���P�� MJ���o}Z�x�߽u�(������VA<��2�Uu���Me�~7b�4�����>R�V��)4;)��$�4�xլ���?�1m?o���@�k��of���ڕ`�}j���G���,!�8�
iU*X�0۱�b���3373��W
P���R�j��Mq��Ӵ�Z��E�)�]���?��8yˑ.���Ǽ&9s��ߕ�P�
��#��"����w��/����3֨"���u?�Lͱ��x��p,�|�����}R��@^��ֽ��<qB�旱H�����l���>ݑq�]��#b�J��KL5h���%ʩ{�>z�,0��B8$LA��|��F��$�=Rj]P�y�Y҆�G�S1\4�L
k!!(}ykJ���j|G;���)z��4��_�|�(Sy�-�zW�=�i<졁�k�{V5�+p��jQY\�E[8������Jf�_^c?~o��q���ˆ��O(@�9�F�ų,jQ(^�?M�Bi��Ҥ� 
<Ƞ���L�aU�� -��M��f9�!��&ͥ�����+�z�'�sg2�R6h�����0���}*A�Gm�
�뾽Y�Ī+ܪ�����DH%�3�!h��R��~�� ;�Ծ$���at�"�>zw���2������~)-�%lkP=�Am�mm�c2u�� G�%�9>��7���p8. �$7�W��b����8���Ŏx�D�4�<����r�o;R
Gq��Y���q>��2�3D�ŖO#z�g�֓�pR�u�6��1����,)Q��� S��rM)�~�g��Ajֲ=8:%�?8A�����_�o�O���c^=|��PI�SX@*4:��.��ߧ���.�H�	ݫ��f��NT��:���O=���O;F�G�(7�=����u�=������k@�޻�:���R�o�ӔIF�������Ԇ�p�/mn�6[h؜_ ji\)��I���V������v �VS�6�eĩqz\��Ǖ����i��@����˧�ˠn��f�=D�
�e�"d��4Ӽ+I|����B��/}q�M#*E���2�4��~S&t�D5�7�X�`�őF�V�E��I��7�:Ц�Te�M��H�껂�H
`,�����Ab4A�+N������m	,��f�9�̷-hC�7J]�~E���fhQ� ���J8!�۲��g�["�?4 ӓ�E�''zӨ�A#)a��^� $t���MT˫MwԱ��e��@��9AL^�M��_�����:��R���Pe�?(K%U>��85W�E��e�(k��3�����=����W�ϐ�Ҁ1=���v�G��D���S�H"),�vR{��6Q���Pq�a�<�g��͒���"�߬~T�p�_���>/��P��@��W�{�g�ů�P����vq�Ҵ���-��щIǗ<C����3k��6�U@q>Z��JJ�nFmi��1�:��A���{љ��pb�)E"v��\:����m�����V��fg	�EՀg��~a���+ٱג���*��ܪ�RϏ�������T)S��M}��B%-�EԿ�+�k
�zʻ����P!a>�:Q{H�O���v���d�i=2x_�[�M�3=���-Wېu�!�ָ��~J���6��5M.!I1���ן��n�7�['L�f��������إ,	+�@�r&��\��������f��0-V��=$	�V���2��+g|cZ���z"f��l��dN�\u�t��C�$��ء$E�4��)d|>����?<�e��h��� �����}���c���౫���b�zl*)�>sT�r�co����TD���_c�*���Df+����³m�pj�ENm`{��P[�?p���u:I�ճǱ��2��1Hdl�"������Zh�@��I��
#`�O����ޖXFM�fW��G@��l8_�����ݱA;�����d��FE�����"���$�~R %�t�N�(@&��(��&�}�L)�q���f ��1���� ��nİ�K[u<8��.��U��W���2$]ߨ�;fbT�O7~#�M�kPVƽ����,���1q�Y��M���r���i���k�&�Gd~��>�*!��
Ct�\�'w�k\2��>%wo�M��� Ծ���H����p� 	H��,;�l�γʶ����������^��Wx�L����H>lǪ|SV�l��Lq����,�n|1�)ku��*H���Mj�iu����	�w���q�<cJd_sک��9�v@ְf�^E���-�=	r�N'ǟ���r�;��K�6%^h,��G5n\�z�ݽl]���2�������x���=9٣�#@�JJ�>T~�-lI��O�����r�Q�͏�9fqT3?���h����3M=�D�Z���a�cCc��%;��w�KA��]��DY{ �����6�F;k��!k���9S������S5�YI��^(ht�J)aBJ�N���
R)+��������/�@�	`����Xˮɤ�@98���-���(��݈Oa*�5���w(NdK��h\GM�o�F:�k%�І����+U�GY��3=���P@�>0+ۘ:؅���o��iV���^0x����\�X	8'�W̦sk�Q�GSj�57Dt��˞PE�&�����=� ����.*����M`NŮ��zA��m7�p���	��V�@�[����r���=R���1���PJ�!�|4R�$�c:�\L���v=���
�r,n��{��L�L�y1�y��P/ee�|�Gkʟ��σ-��j�H�?6���v�[�G��A��-�I#���0k��S*�"��}]�y`�s�.Oe�8t�| �J���2�Cd���1��w��SH��L��a]ň���Oʞ�b����:#pDhG��C�cV���T�i��3�9Ս�.�nΪ�U�~��cx�����P�z<��Y�2�$^Ǖ-�:�����K?���	oN�D�������~t�����.~K��ڣ�}���1�AA�&,˦��|��w������HIz�	�#>��:��/�R�x�����YnWn��kө���5Z�x��7�/X�G#FE�Z��K]W���|���X#iU�!�{&s��^��ޭ��I+r׿t��Bya��$.%��YdA�$��[eI�3y�\�0�wQJ}/�j�?g�uYŉ�H�5�נȈw���U"Ę�iFzR	~�sK1�o#���v�r�(�1�Yo�झp�GK�@Dp�$E�Kf���t=���_E�mW K��~&�۟�%$i��l��&��R ���v=EI�r^������qZ�ھ����,�w1�Ԑ��?�`���\�4N�,��u��W�2��M�"&��V�v��靬ߚ�34���/5�O��u�v�,�Z;f��>_Q�+j�w�o�����4/�$�Yc|��.%���,�7ͻ�J:i܆�
# ?x�f$Ex
���?>5Y#��⾀��M���&?�&��]��3aD�k��BW �q+E�(wx�S��[]��`�z�4*⨥�*��|�`���1vj`�85�SXPNjƯf���¦�J��$}ޖv�r���)�+� A\���x ��Bj�Ԛ�Ky�J�� .s�p�L��´��F���Y,p���5/Q�x,�*j)��DD�N���{�y������glKfH&���?@Kq	D(W���Ob گ$����83�$�U�5��UMN�Ο\?��:qu�7ns�x�~���z%�y��&_��<�9>�SƦ�� D���.���I"a�I��6��K�8�O��Co��K-�1^0��9,���F,�E�;���§�`���U���@h߯rA�O~�ey������d��u?bE:��\	8���
Ҕ8p�mu:��
s+8B�zUw7��ęSÃ:�8J�%R���75,�9Vi���3]�ZǙB�	y5�Qy.�cT`��#�}a�O�N�$rz�ڼ�-��84Xy	7|��C/	V1FKMt���`���D�R`h�TU�N���6����ys#�L�߼�\Q�1m���T�iE��v��q(�$l�Y���o�����+�r��Z/����_�̖�r�a�����#RcRӞ����?�k%G�1i�q�A�i�T�S}��{	������*NW�ο��2WtJ�e�mroofA���Ͻ�.� %XkO�z��!���$k/z��i�q@�)�ք�m-�������8�Cߔ�d���<�����;&.\p��◗�E>��
��sF��2s.� �=(�0/�G�4�hJۯ-��� h&�bQ��4=�K�X��~�44�����cC7��+��Y�-3�[m�ef!m��c�x]{���@�@�{{ـ
��k��2p�
.V9�췅�q���k4؂h��F��89�o6no��C�� Wm�J/9��f[X�!|Q<kbؐԍ��򆩧��
���X-`]�}G�?^��UJ�
��T����oPxn��!O���A�װT{*1��I�Wrj��G�y\���נ-�k/N̲F+%q��>��vD�S՘�v~�f�hOa�� �z�]��H7K70�}[�k���Ex܂��azl�i���uř�t�m�����p�٘���t�EW}&hD 1Z���ht��KC�<Ynl�߾?�(������7�;�m�Sh��EQ�N�"h�/U)�q}�����@p����R�X�Ss���o�/����g�� �oO~�.f��F�8�����3��e}l���í!��խL���ӻt�����z��Üt(��q�dz�"fΧ�m�HF�d瀇�}��z;����9:�2����ja���u��ɕl+����}i�bL��y�<�A���A�-�}�L����8$]����Ż	���8!�
O�J�Ʀl`�f�'�z^�k��>�wG��0aKGhr-n^�EN5� �j��Zrl����w���;-[�"��}�[��n�\y 6!0��I��Hǂy�Se�g�\&�AA�P6��g���%�4&�"�6�v�y�TuCU1������eX�^$�􋱡+�L�-��gxT���󯺠��:8�U�< KXF W/���\���";K2���o� ճ�֚���O�nfC���6_���bAZ�+Sڨ66�y[ M"	\�k�Eʹ=s��ӆ_(���'A(�r������"�f�@�I�,�r|���NQ�W��GR�8�rS���W�������?���w���L$��TJfe�-��!�0j.�[��3(D��|G�Y�r�K�zN���+w��1�n�-w�T�Ig�^�Җ�{IUP��N��7H�O��D�u៟r��N������(�%M�n�P-/��aX�Ʉ�ː��fX�tO��;�s��㑂������x�a{{��4��^�?��|�D���ߋq��v�Q�����DͶu��~l�b;�� � L���Z��s��~��7�]��"�)�?r�?m?���E����&��t���Ŭ%�-kJ�ᜍ�7���Y�R�_�:�Wu/.4�X�-�
 ��m�+%8��:��5եԂ��0��S�Ϧ�PȺ�z\��n�b}�M��K-��9=���v�kkN�����a����!.���zF � F�45�C9g�ꅄ�Ĝ�0�AZ�-̕����b��01�*����pP\�9VN�#��]1,U�0��31�Lb,(|*�n�<S�^�/g��㣭�e0�'"�C�?P��aTUS�΀y�0�붿��ǌP&�Q�Em�!��z<̇=�>EF�=2j��TXT@2^����=�\�X�f��bB��|��<<�@~��q ��M��G�� R�G���NE�|s�qB�5=F�HH�[^.P8��/[�鮆�C��fCT/����ٝ���Q�z��a������-==���8Șڱq���⻋G���XzÁ;]��Q��L$H�KP@T�#T���p���pI��­B��~ϼ��NWXD5�0}ui�օ�.q�u?�9RNW|D��}��)q�td�Uj��ED�$zWÆ��WA����KL��ԥb*��/|�u�O���c>	���c��^Fb�
�w��B�2���~<�F�k�� �l�L�R�	�6OV�a����W���n�|�?�l��G���=�~�����l]��o�~�UV�v���}R]�FB���QY��6�rz�UP� �31]�a��3�(:�hVp�v��M�%	c&��N�Гh�1!��^6�>+cy0�7�7hpEl7��1I��Lu7T$co4;�C�c)�!D�ͨ컾�ʤߎY����׽Ę�m�@�:�:����>�|��})����Kz����V���
�7z�+Tķ�:G�ݑN? e4QU"�꣓Q80敲��k��R�P>pǮ��ճ.b
j�~�	/�H�HDz$O�O��&�g��[a��W�k��'@��/r\�-ʦ	9<au��]�!n�x[)+x��p���_l��:
0�	2���q�W�Ȥ�Y2�u��E��ZC�a��|��X+$��'�J�-J,ye>|��]j��?�2+����owJ�����<�­�V�4v�aε&ѱ�֥���-(���sD��]����;-�Js�%�Mh�z4d�
�7nb4��]�2��������y`���J���<��N���Vx*( ]ʼԌ!s��KdsR2���4d��6����,j�T������Se2�<������f<�s�u~o ��Lk�ŀ�d��ϟ�g�٘w�"8�o���RX���]�� �E���D��