��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|ḱ	I*�n���}וLM��!lА�(��p�&q�;y%�(���)��_��>�>�l}cp�o�6��NO�3�r'{��?�u�>n�� ��<[[0�¿!�csY��[i̺'� %Z���٣X�gG������v��VW5a-I扁k��Η�4�~&W%ns]8ev1�:Sm�&^�RF���B�Ț��G�s8�+6��x;o(D�>+��C�����dP���5��G��+�(XeB��D ���Kh�v�����L��9?���
}:�A=\�-�,#��Р�\|]�ν�SG�h���l������7�A��O��d2M���%ط~L΢,�=9��.t:��O+������e�4��yqM�C�C�G��o��'�_�I��w*�6��~4j0��.�ݯ�+���1$+p4FQ�,2��t�Zv�b\v�%�c:v\l&�vC�D��y��"h�2xVH��ŕ���`V��.A�K�����E�F�O����%���&��$ׅ�m�M&Y�G�ai��=&�x`�ᴩ��;&%��%�`̮<ب<���b;��G�m�K��"_�o�
�	�?#k:Z+���VCe9uu7	x�}��C��`R s�v�Y �&�L��D�ZsI� ���ha�]�Ϩ�b�u�\P���fdz�m��t(�$��l��^�ʅ~pl��P$Ѱ��/t��g�U�o���Ba.a�L�~IɻK����p?��r �3�=�ZVD�dô�F��At$�߁�K{7�9�~T�-?��P��MiƆ��i��D��JshC�yȒ�3������"��v�Q�Va���3�B{r��P
Y�MY-����T�6�K����m�7w�,�<{�P�:d��S���^�]*u���&ߩ�廋�¥�U��;hb�1d�ܝ��!����~E�h���q��_���c����]�A�,��()��ݫ����\��{��X���}��p�fX��RM�yBn�Lv��. B��`W$b�5�"���!ea����A�=���Q/@����:��/n�<��ѬŚ_>����?�0xǨ���ms� ��Ʃ+_9|�$�G|e����9w�́��h�jn�'�����z��-�ܭ�)U��Ճe�;>(��<������+�}Ъ�`��+�8)Ɵm8R��]�$N�%B�(��`v�8�s]����1�(���,ږ���脓�4~����s�:~)��� G'S�b���18Vh������)VY�0����#g�T�~����w2�u��"&}����s'T}��wS�ͭ CH��O8�1?�os�=0�p�}��/E�A�=r'xv������*��E���H{�"u>8�+`:�6�_�"�#��3ӽ���8'ɡ����bo�?D��n@�2� ��ތ ��O�U�g��f�l�\���S���@#"�xyt� ۣ�W���^�|��MQ^
��#���ßG?W5,t�E5>���$�� ̈́/gd�CY��V6l�����ܴ�aJ�l<2@\�T��`��t�`�f�y;�ےpWf�h���K���P	����}�Ro���$.�"��P��\�_�f�zAm�ܩ�`��6�օM�j�`A{\ )�f^"仴bt��$�����'`~�YT�l9�n��r������vTQ{	�ⷵ�l����։���eP2��z�ޜ���/4v���e5����CЄ����t`lZw��;ѫLw�g����i����ЭnХ�r� ���[/Fθ�(.|h�A2�nU�5Z���<�I��̨��~�?Ju�<�(�B<"��o_c��U�}+Ke&_9��t>�,�Z���s�+�k����ô�*&��.�	`Ѳ��y���s%�|׌B2������L�h����ۺH��>,J�[�IGRݗW�}�*i$�N��.F�!B�4�=&��y$�*E��"��^�'/V��6���6��J0qm�h��2��d�������A@Q*�dcņ
̸U珊&t���M�����|���L�V�-���K�b��0ͺ�0s?|+�Ԛ��p9a��}y�i�ܷ���2�Qz��*�0�X���E�������T����R�����r�ݍ����Hb�����0UB��k���i/f9����.�l1��Q�����dg�рޓ>�3�H��� �w�����87��q$�`��G�0�S�>1�T���(�� ��w�s�Ҥ	 ��~�B7�df��S��c�A���r�z����{�ߍBH�ڥ|�,o�Z�K)k�+�a�4��:*}|�qJ���Y��Nwy���m�@i��Śu	4JB���h�\�����xeH55����RP�c�7���S�i�|<���O�9�!릲^�C�&��>7�<��7��{�Qˌ\3�Xh%6���	�L�ک������V��zE=�~��"����qB8�y1���$%��1��q@s�Ά����ڗ�Q������e�J���~�9������G�I���Qc5W?����4$&'t�a�)��[��7|�)�W%I�����P��-1n����`8O�Ʈ�V�� J��xxXh�R��p`P��G̉Ț�-�p��у��+���� 	3��#���
t8Z\E,�$�l�(�5�
xOAcz
 ��]%�B����j��ѨK#�@(p�J��Ѱ�w��j���`D�/��W�9�ˮ��NՑ�4�(~[������TW=��[~L�[�����l�h��vzYPg�N���M�v��\�!h�SB�] ���g[(���	��E�`h�~�˝����8��J�!7>Tnt�&�D*����#�Ҝ:9J�ԅ���e�(��9̭�SK�����y�Q��^U�D�1)W33n�*,�D�.b��A�@ࡑ�w�^刑�ͫWI7�j��-�!U��9��)�=5�0g�=�j\�s] ����V�������k�G���$�e2�|0+@��wO�;&e� K��)V��K�O;���O�Zz�;OV��`^���]bg��d�/��)<[�Ea� w�M�E�`x*#�$e_r�ؼ��6ȡ�#e��?����
ʃ��/�F����m�b�
�)�Z����������]���z�C?W��O������F�����&�e�)bS+�ȏ4VVE�*40���ݍcT��g��m ���BM� R�o�Z�3c��x�H���[Z����W�F��h�V����<vCt��"e=Sh�xm4��ۺ�*6B1,�I'j�t���)����%�pP�ԧ�&
��M>JO:Ϲ�--�8�w�+<wm��kB5qye6
$hU�勉��>L��q�ץ	�D�\y]#?�-a,܋	�ma�iU
a:1�N�!�F�?�y^H���࠺]&�>�}4�ßm-1K�x�w��X�� LG;������e�e������zEe�qr]HDc���=�Ţ�w��$.Y���:�(�*��'��a�6wn2I����0�r��c��!!%왾v�����R���/�WK;��ː%c�;�Br�ղ�eo\V���L��$� h��.ϖ;���Cqi�{B�8m$vE��l ��
,�5՜��I�܌b.j��q�H߅s
�-��Υ�⒞~ip'q(,��A˭
�(*�{yO�7Mw��\�w�dQ��Ip��˟�����I��Z&��o*�K���,W|^(�N��8Ԟ�6u>�6@	��h���z�N[����#ZIzb�@S�+K��-��p�|B�Rŏ9�$����z��'Kλ �-�u��8b�s1N)�Jɮv}ɹj^�7����~_<��g𞻀��܇9�w�����:)!K��Q�F�>n~��R�/�
vt��$�p Y�Q��e"���WS��m��J�0RH`�0%J�5(���9æGY���Ykul�HYH)-@.�DC�px�@)�X$��@[�f�>y'��j����F�u�1G�;�,ml���E�(0��&�ӳq���UʚiU�{��ѧ��!Y�oi�ȹ���GS܂��`b��	�������F;����Q�^��Y��*�\�
e�/�����j��e�y��R�|J�~�K�*{����߬��G�G����-β��?�N�+�>�1�NJ ��_z��V,�T����Ƞk�'f��hp|�~�廬.�f�j�<�O��3��z7�t�K
���������m+��'�O��ށ&];���]P�ZUHTnk.�:x:͞�eй�>ۄ] �ʸ��$Ok97��|N�s�o�@�FA8���)��1���|�vCG�jqh�����O�<�h��)T�=	�'˺����e{��� 9�?�p�̽7��;����ϳ�V�[&�l07F#Η�'N&f�!�t�i�|M���Hī��?F�JP�{��[�QĚ(Q䩒|'ε���PS�-���sM}����f:D ��Mr.SP�� ��b�4���[���gc�(ܫ([�ԣd�GJ�r}+�0�Ƀ̐{-�-�`A�K�M��d���_��c��׌�Xg)���;�d-/�S�����	���-�;��x�qV�S���j����6����paֹ�����v��9�o�o�タ��j��8|ɗ�����0mɘ����E�^~:��p��򈚶�eTe��^�1�u�}�|P�#��kdP�ĘT������Ο�4�~ۙZ	�-�_�'I�Z�z6���K��g�q��EB���U�:�Ͻ�+2��g�+�����H��dtݕg��C�l��J_���\<���98��l��>4���FW�w�xd��er�q�ι/�D�L� �|ꡁ?��:�PV͈�V[��6�q�a�&������w�y��������r��E<��;v"mL�����٩����{�a����~���6l����]��Ŋ6ɪWSJ������G��g�b�5�6��O�s~vZC�j5�Ӱ8A؉f7��5�{
/�Ú��ˇ�9��&��^>��C�U�k�o܀\-զT��^�������5;�Q)�8�+d\&��-�n �� -��򻗳l����Ժ��vrT%ڮeA[�0���*��O�up��2��8] \|�o��B����t��R�zO"?��S]�������~u)�_��[�
P�\>ٗ��v-��JȊ�{*x9���Q�$p����ب,�B�,����:#�mO�z0 0
��rM�F�OX��%���廬�F�6!���xh���qhA3p��jG�H偅�.���-��)������=�L�Ӭ��Y!1��X�ȻT/;�+����m�y^W/ �����&l�A�2�v��I�~&������+= (�~� �5�?`{���Z,%^�%�0x{��Wrz�H�8���Ѻ�׸�:J�d�Me�P�/_n�`?��mrl�i�Z
���s�D4i �
�t��K�M�sn��d�P�B�ƪ�b��h� �o���[�,�W�C3�=%(����f�g�*�|c-���8�RT�k�x�I�i��k��vR�I�?T�߅�l(�?AGy]��gxM+>e	q�]�>C��&j"�Ι���+��\pP�SC�E�?KA��l��ߟx�\3�������&D�+-֌�9K���V��4�늃��y�е2H����{��_Ni	kl�������p^G�kfta��2dA��[�Zn� gQ�0Lﷆ�S���w�]+ ��.���q�b�M�~q�
�[Wo�0�_��#�a2�t�St4���#$Q�I�Xy�L҈�<>�5�Ȭ�D/��MM���9y���f�����a?�_65�>�5� ��g�Ek-��@�[���B���Z�&m�!��Ho-S��Д?9<O��=Ni�	V5�����N��B<�&��km���2�V��fcFE��5.	�ج]���p���D	e{G��0�����dh�nCǙ����Dp�8)��W�q�g��/�~�S@��2�I{�u�r%�d�$4[��鎌֮K�\���E2t|���QcZS�m��T���9���J&'RV�r��'C��51���Y�x��(�?|k�J2��<ۃY5S��g��w���"dg��mg��BP�Ն��=@�U���%u*�
�>Ѳ)(��Y�};�=})0��x0ӼTΌ7��$p"�q�뿪��j�7:	�����q`�5�'�K�]CP�m�����/��o䩫%�x�r�,o�*�(+���N���.��<�4��ul|2�ͧZ�HZ��:�3-�j2�P��� �k�����֟�XДF��"&�s@D(ފ�K9��D
f)jݚ �F��!�T6/��J��3`w�M�b��i>��Jn���Hu8���eA����S<�D��I̀�
���'z}\IȆ��!��i�V�#m����ȥ,ʁ�Es94|c��OiJ*6qW@�({��6 z� �q7�
 ����SU�'Jڶ�ε/�����̳�B|e�I������/�{�e�������q��H����5f]8$�U��}X�����;�HW:��uJ�����H��^^׃R�@���B��u�m�\ 
�l	��uR��6"�Ǘ1M���I��ލ������Xz��A�(~�ֶ¿��@6Zz"S����6T���")���4#UFJ�P
��=� �o�q��b�z����)�:�1p�a�\�7�"���e`%㨚�]��Ns����#S�<~��O�o�V�2rn�������6dq��A׍l�¨�s#b���WI
s[EZI��6*V1O�9�?�@��q��O��g\����	���ͦ2���_e�0;�	ze�n������2�/,�Y���>+ѺL{h�~Q�%2�B���Ǯב�����(�jwUV��89�)�H%d�cI�������0�̤���Ȕѷ��V��=���ADniЭN�W�Y9Jp��~�/Z��"r�bbUu�i���F�:S!���4"?~��Z�}�@gI�����å1���^���uV���j߸�D:�4�x��_���H��ג�@��z@#,�a���`��^�K��KH���BH�t�l�{�]����sc�m��1"��cWK�4�XU+��J��4r���	��F�Ml�\ۦƹ/�n͜�bt1�C�b`*�rW	���<�t��@�� �z�n�������I��Ȩ�F���ZD�+��y�w���V�4�#B��؁�<��W���v�if)7�6E�W��}���D�&8H��`�����O���Kw7UZ%���T��8 r?[�����|�S� 6Wu��YG%{Q��B,:�'|���="z�N�P��F!���o͜r~b���5�*̫��l�[�Ҽz�m�H�=݆h�6�u�-���s�?�\�2�L�L���-�m)�ZM.X9վ$��d�'#��DƟ�5�"��>kʹ"L_�˦�|�2��Nw��ZF�}t2�;���"�+^|��q��}��v�0��x��)��V4+�z޲>Mp�lc�Bvy�8���V�y�y\�������8?;<��\��{�Ґd�0gq�D�R[*����O�&�(Q�����d�*�//#��q]����ӹ�m�&���X�1�3��Z�Z�R���0Ln㪏x�';�={�|�;
=�	/t6�`T�>��JZR��B>����Տ�?����IK�&j�?���\���]��)U������Uo��8@[0�.��[4�m�d�3ײ5�,J�����t��fXlLOڤ��a���KP:{Bl�O�S�m�L-l�y�q�r��z�r���q�j%���]��l)�x�>�a��e��6k;��:�V�P^�{����^߈N�UMi�
�s˃?~N2�3���ɲ���*�=cA�|���r	�GC�m��,қ�y����|��
��� m��{*�3�#Oì&������yϐ\'�Hص{�s�y��l(��i�T�e�� �r'1�Xe�:��*���X�ߜ���ߟ&gq�JҽLw-�!��G��4]B�1��2�G�Y�WN�K�7���!�M�'5c�����_KN�*�Z\�^`�2��Qg��)_Y��������]��7z�-@�T퉶�y�d�3��#/����$g{ƴ�0��o��1y֚��+w'X�D�Ve5y���AZ�$��=����
�\}J9nqE����9v�pm>d�GxI�v�.���{�<�'2���kD���@o��������D���&��pu=�`�4��Lw�v	��ϳ����q����y�ym�z�X�/ˀ�4�՝D�D	�,��LK\|<�A���D���*"ͽ_���w���ߞ�F\v����	?���O3��4��b+)c��\��	�w q�H�PX=V�	�"�tZ����E�	���J�#���i��C`'E���U�B��1�U�ڋ�1�Ӂ���E��l6��t�+R��8ƝUe4�����}�W���F�᠏���í�ܷ�zM#����q��􇽯���J�eɞ����� �a��k��P�mЂ�Ŷ�G�8���A��(�����U�c�j�g1�b�6 9(K��"�w��?J�MM�MZ���QY�yz
i�} _�P�' )���o$/�s��`Z1T:p�ѹxp<0����t��!gfQu�Ϗ�W�3~�%W�I�(%L�����%�A����~p���w�4ŸB�b��^b��.��G\bG�>B	ʘ�V2��<Rt�+'��q��JФ�f�D�4��:�%��e�_��="�wUM>yOW�B�U�w[�W��~Y@�����/�/���jP������{b.4U�^Z��tdC1]��O�� \��'���p�� %��,CR�ZQ��t���ϴ<�Ѳ��/M��c_�ʲR�G�@���_v,�k�~��XS�x%���
�9K���v&a> �^x<�Đ��Tj܆��ݬo��k�H����;��X�zQ��{G�e���ӭ���.#�O&!��Z��J7�V�'ۺ�`1�c;��jWdI��2��R�d8S}"LC��g�֖�Sk��l�xA���+���B��n^Kڡ��D21r��]a���ᛡ��X�q��%��ǁT����R�%�4��z�%�@��5�plL�X��&'�؋Z�rV�yS f������h#r�%��D�Xၥ�#d���#��o��P��T�v����M��b��.��3viH췸��B�J�Q�O�_
"xU���g�|nI�]h�_�8��Z��ɲ�Q|fn��� �լ>��zb[���>Y�����|��rN�Ol�/3ţ��P��d��2�w^�A\P�J��tT�WFl��b3\���q�7�BO��`�����AS�����@g,�xҴS����0�gea��o��DH{�1���{o��c���h�7 ��C��Eg��Z���U��N��i��%��W�t�k�9�Un��0�g��<���t�qP7����^�*ؒ�zC�.�RSz�$��^�������i�u%qB�5&�+}e%x�@����nz'�,����";#W��3�~W,���g�CR��0E����X�R<��Q�=4Z<�z��V��G�6K��j@�)�1<�EȦu}2��p�b��V'A�u�i 9����#j�5��lI��P���)P�zw?wQ^֤�F��jvr���
�cx�<j�s�.����ٿM�3G�to�=���bv7����@U�O��W�b�CP�������Q����%U�i.�ф�^T���MlmFO�f��/N-e�o"nn���w�}C]x�L)��2���w�<OlNI�Nr7
E�&�e�5�*��i��_GD���(���V��y�����N���BTώD��,?o�����YN��C(߄���3�,%=�U�_s�e�0�M�y]��$��*��9���v㺫
�u�x���iɣ���4n6�g�{�45f-��)�훍�C.�+���-�k6�^�{���i1!I��\�z%2�y�&��@T�7��Їr2�'��r����&�}|������V��2�m��B��ZzV;o��yd�0;������������w$Cy��R'���=KO9��'xl�U1�����G�����;64K�sw�ʶ��;ZX��#��F��b�CDSrX������ωс�����ߋ�-lɂ!� ���mk'm��<�dlnY�[�b���?Ӑ��Bz58�����To�(�����$̰MU<���4�>HR$��3��>ɵ#R��0x����ʹ�L����\��<Cu]H��$C/��3�����Tg����s?>5�9��k�̑z���#��!i��q��)!�^gE�w���7.��[]"��'�s�}�����`���6���*'%�W%�),'��f��<���v�� ��FNC�� 1Ё i�"�j�R#l�3�ЭHb���B�-�mބQ��8h^+/�`����|��&(�|�LҳlQJ�7cʑ��� mBl�����eZ�c�	݇�2���G�6���h�Wb2�W\=9�Z2�!��Pf幅����y�ɤ�F�;2��upe�Y�����,�4��li�8���yꮱ���ٚ|�g>yQ�Aq9�5�O������`׌�Tu�BO��b�i���.+0��2�(��@���_�'e�3�m�x�q�z���}�W�.�;���9��f�q��N��M/�7k6��8w*�5v0'@�P8�
�u3����>͊$i����~�� ԅ��yoѢlUW�dk��a�9nN1��;&V�����A��~D�Rb��"�s�U�u8ox �-����F�_�4K䊕H�R�������,���$��l�M*�S�U���9$dy�;�U͡CF�=�\R7v-�Kە�'`?߁�} R�ܝ����^��5�S�'|W��7�w����%���?'yhme�#Փ��vOF�� �P�$&����ܾ�B�����>�cw��ַ�Y�@������
h@���\��=6�e`*�Ou����Z����P��\����9�� �d��o���ۂ�4��f�]��J���U�U��h�2 V�������IG�)�?%޳�wW9r�8���>i�6�>����O�C*/ȼ���[�e��6:�p��@zb������{4�Amp��j����\��T����������O�o�󩂼�D���2�!�T�#A��V.�����j3%�	L42#Ec2N�c����:�R��z��,���'�vL�Ƒ�tV�'�3ֱ!��D�ӝ�C��4�r��cs�A������z;�F�ҭ`A.�C���d*�H9-9;TA������#'���������{4j�RU��B�����1'���]N�� �ï�͋�L�h��j_ALx�3t0| ���|Ȍ�����H�yT��͈�|�<vq�,�LB���v=�R\*^F��i*"��@ݘ5�`��H�t���ۧ��UʾB��%dY��" H�ҭ����\����w7��R�rϐ�D/��R�;	�mޫ��m��lҾ-���������
]Ϩ�=�w˓�lRa�x�EX&p�������ޕU�s�S�M}�������muN��dd�G�أVE)����^t0�	qOGtoKn�B�2�<y 5#^Ǟ��Gg�L	}�כ�G����ۄB��y$�T[04��޹���s�0�̑��Y���f�֫�Ђn��R�Ϊ�(���`2��n�\E��Q%(B���kl�L����s�b}�?Z��O�U�6�2�<ظU]�]�-�P��Ys������d�ɦ���P�=_�0,�T�J}�[������O��l�t��-j`-B�S^q���J%�ӕ�E��݆�H��|1!�/��D���n�'��e������$U�֩�<�`�`��J�C��ndh�-�MN��xw�iP���M*C}�jm��P���9%����"�V�`���6�2f��#�K�z�!L.�1�,x0���5��k��I�� P��o:@��Ǩ��|���O�4��6���桜�J䂛ƙb�O^"s-i%���)E=�ʼ�|<E���Vr�=Ӭ��_�$������<���軇���n�DZ=~�$$P���푿e��; ,�pjT�k/9C��ī�T�w=;UfA��VE����\Mp� �$xB�A|��ڶ��Ε����gHOe;5�����Q�\Vmg����Y��SV�]i@��Zy^9�Bi�z3*d&٢�#�&��T�^w���{J����Y��}e�&(I���w6_��6��c�Ӱ�D5-b���h>���^�]w2��Iƍɉ�*<��ჷ��H\|�����4Ǖ� 5��] h��v�:犥�E���ho��:����Ze�OA%�׸�(3��S֔�����C��ц}��������x%�X��#D��E>c���>P/[ɣ�3�X�Fݡ��T��y�aƽ��^m�����:mX�X͟()�(}��y�����=�-r�u�{���;��y51���H�	S�� �B5��w�u��Tl
4"/��5p�y��g��]���}�g�q��:��6�T����@r�l�:�"���WT������PD��������X���l�'��Э8"�Lc������b����.�b]�X�LBxSG�Zܬ��U��$�,�*���S�>���� x���Au�-�0���'���8�Dd�ր�J<$�'6��jHܷ/�AH�u�߸C��Y6���r������[�hp[t�U��a�6����O:�����K��W�S�R���*��#'���C;lK#$b���Y�d�8�ӽ?Ȉr��0����<�:��Z
L#�"�y^Z��2I�W鍭��&����v)pmw�^���#���?�]�#k]�r��k�����\ar��6?�և���ي��Օ���S�Q]�+����2Q_�C�KG�R���A�qҪv�B�;ԶT� ��$Ӫ��}��g�����p���A�F���hm�W,�%Č���zK)ذ9'����4�[10,ڡ�կ{!��fa>�{��<�pߚ���N%O�|Gm�q��]bX��#qb�h1%RS�s��vފ��ɪ���[����z���ʡI�C��\�:A��{
�F��"��+y��2	�y���1
d�o����A!�TM%?� �z=ÓS7n�`Zm
]�G��]�QY�X�n�I_6��1S���KCΒ��Q�/�c�,�3�����x���x4��c�:}dx�=tM������Ԣ�%�W�4���M%�t�@��YZ�V�^6)z�߃�0)���ȸzo�Y�fT�O᣿A
.�t��Ws& ���/̲vXѕ�z�z�m�U�a?�H��r�����l�p����	[L�Mf�yq=
��ɷ���rW�Z�H�A��9�D�m6ȓ��\�v��wNd�F]t���OS�C��||�d�RmXX��z��&u]tr:�s��=U��g��|�z��a�9��C)�����x�|O�|fx�+��ã����B'Ż�,�4ݲ�Ou�u����ڑ����9un���$U�DwaN�T${���ʥ�וq��}I.G�ͻv����f�t:s��$z䳂9e[P�Hk�t��'�ȋ���iҲUl�
f����������$!%�p�(RR]5uw��,2*'Ș�A����S"�EAJ4��8�G����Z?[3���i�9mGEO��+M_�[$Yt���qR��
�g�����}���+�{O��܉�f��(�^�D;�(-��#���)��q�g��6�_�����ئ��(8��f�=���Y��C�Ln* q����3��\�׊g�Ӷ:�)Q���P�3K�,_�����0��W�{E��R��#����9�/)�9�5]be�"�@�e#�V#ҥ�3� �7Z�����Cn�g �b��#�����1����>��vy��;B�-͸j��`�/[�%3�0�EQG`nc�J
.
�S�mz00�d�#Ӕ��9��(b���-��αF�9Dv�񜝪��ƿގms��*�50?Kn˥]d��xtnc��H���L`ݿH���G�Q! o�k�����4��ݦ��w��g\�/b���Z�z�lC4��:�m1�W������-";����-J+`�t�� �	�~�w�}vGKIr��
����z��|���*��n�� ���,�A�u�̛ҊuD�c9����������xL8ts.�����Ρ<�xR7�����u���n��}���lK���!���_�G���\A{e<b���OX�����d%����l8`"�?.�qfӎθzBx���@=��IA��>����X���$,��/^�qzIO����c�Us@ѱ���ZK�����J^9��aa������s[��7*���dq�t@�f�_р LN��x��$�g6�o�7�Bt킌���U���)�V�[<����p����F�(>�(QaL��NIz��y��>�ɨ�����q0�0��@���6��1c�d�|�����|�D�ڻ��YHK�R#�yWts&x�Y����@~�T���p�{�d���?``F�!���8���2�q��r~�K��L����c`m:�7�"�%5U�
 ;��Hܳ@��]���N��[��`NS����ZÒ�k<Z?E$1p)=��p���c����N�f��B��<ג?P�L�Ԇ�����^;7��37�;R]���RG׎Te�-���ba9J�7'��Up��j�ͻG���:��m,�/W��^�}^��m��"���g)�ד ��x�W�u����G5s��rq��>�	,J��T�-�!&&q���v�!F���uW�24֏iE~D��uX�Ŧ��k�Q�7�[.�5
�����D��gn1m�wU�!��ī>��S���Cd��ܦ*�5��	
ݥs�rLV �25χ��⻏�NE�d��^[b��@f�
1D�	ȶ����J�� B3�/���q33U�MG{m��,�|g�9j���ЕR���Vq]�{ JPP$׵$'�o���S #נ訶�*���a�}(����1C��y�����0��0!#��އ" b�kK<�p�}��A�����-e�&�t�B�ƽЪlS������3*��M��J���J#��у��yd �4�%��G�%��X�|��g����ez۾��l�R�͙�Nϖ���s�����)���I#�ɻ�o��F�qaj]`�bc(k�ķl���L�S��9j_i!Q�{xNuJ#po�p���:�����IƇ( gl�`P���
�O�wR��;�D���*������5��a@g�o��~խ������l>��&����A�ewLF�����_�D����΄;�-v:W�-��K����s���t�iV�3�rߦG�9n����GY�S���ŏ�u�г��;���.�`���F;/t���ZNBbwhyiGP=��s�[��k��'�Q��ߜ䴝�!��-�`�;�������/jl3��uG. ���d���j���b!	^r��?�ȜL�O�2Izp	����hρ<�2#M�N1 fB��9T����t���r�����֏��9��U�-�Ǟ�H+��f���c_Bo�����x�j�M�?� �O��Ƃ�a@S>��Q��gݘ�Z��ɾ.���C�3Z�~��y��׳U��lZ̯x�S��7e�9Ҹ���i� �걟%�B��z��i#�9_�S��v������Y'\E&YO��Bp٪7N�*w,���?7.5f�G�zK�� ֚��~
���䣃���K��y�a����$o��w��Aꚃ΃i�m����]'
�w�f��/�~t�(Đ4b4�a*�~�����-��N�1��i���/�S���[��h����i�Pm�v����7�*�1x��� �+T��$2IJ�F�SU��p.�d�=(C��e�|c�<�bB,��77Г1X��gn�*�k��?`��0e�0LA&���>8|�)Cct=�t�:��X��$"dkU�2^��e�$%�����c�X�����EI.���$�7�ơ}%I���&M��Q��;%wo�V�T����.�f�Dm&��4�nKT�뗬O��&�X�n���`S�/�9vf����S��El��S��O_P�+�L@��ayj���P�M�{�jӾ~�|���^�ˮ���1��q [SF*U�k{��~,»AD�\ �}u���D��<�[^�=�S�Sj��$�%πa��k��66kz2�S*o+9�a���/����<!i�j��1�\�,X�DK=�Zv�����Dsr�24��E�I��3��%3k�2&���x��)�\>�S���+,��j���5���ۜ�Խ7�J~�d���M霞x���)��խ�7�j���A ]�m��c!)y�c E�F$ғP�U��\�w�|J���Ǖr-nn�'Pܖk}��Ͱ�Ow����\����<>#����mW*��~? +�H�	5}ay<NR�ui�P�{�{�#~���[��
K෥(�+E�U� d��!I�&;	p���b���v̻"FV�	�D��#��ba��:��"軸�qH��jp�$��{?��6�U#��>����]�z�TJZ�L�@�!Ӛ>������i9-�X<�˒#����\^�"��������D�Ws�S�2��(8��������×�9'��� �y��C��-pC�
ݴ&A�$^���Di��=�I��Q��M�PG&S"�匒m��oD\
[������OD][��8\�M��^�V�����FEg�Z�n?�l�Ѥ'Ȝ����?w.G��'�J!��+G�'�a?#��IY^���f��ryJA._ۂ��Ň���@���a
�,���>�A�����Fą��`��}�C&��-�{�\cۺ[:�f�xط��ެ���&e�r��9:|�m_��u�m���7O-Xk��ξ��\s=���3�
K�S+����-䤲��(�ċ�FH�HM��TQ#U�G�Wp0���6���M���)f����$�<�Gz-snW ��!�Hx��B)�N:ʈ	�"n���=�h2���!�y���It�*��Uؾ�A�g��"&�=��$��|�~R1)�g����C�77�M��/�˛�����x����`/���Y]����_o�Q�|��Z��P�c|�����a���ѷ��i�aC-vxF;��6�g�4>qDx��ǪcM�/���X�|Z�q�Q��t_�@t�G>e�3淼�}�MJ�E���Mh��*���#�	�*�7�^=FIFI� ��'��������Q01�=����K	��W�I�k�4f��UÄ�*�3�2I����M�{�j�!Zy�R_���K�3L���lOZRz5h�D�+�6�F�":���(�[�����0�ol��W��*;r9��N�z���,s�SK�3V�p��V	H#���Bz�Ų�+�N���S6��9�6�H^�C������딶�X�F4���oG�p�2H�R:I���ѓ3Ѿ�����J.�ZqB�n{6{��d�#�Q�0&�91�p�1h�9�Km�7�UL�"���L�+CHS=��������M %����)��$�wb�� �w�C۰�g�)���c}U�ɽ��Ct�xx`��7�����P�yN93����$��^Y����J�G�U�:�ċx��On��? \�u6�7��
���=��>=i��.p����^_���0kj�.�D�kYD�s�h�m�G蓅�D��ݺ��C�bC�pM �EB�o��������In�D���!�!@n�<������z�QTJ��g�#�m�b74��KMF灒?�B㔍Ü���nX(!���8Q�-���k%��N�U����U+�a\�����������X��B���u�#�6�yl٤�S���M�~�!}6�'���}��1��]�Y��e}B�jd�;��S-����߾H����R���7ȓ�O�D��+ڷ��;2����~%��1�*9�b�=�-
��{K���s�ٝ���_��=oL0���/�獼�����.�-#Mۿ�`K#��4�����pSS��]�ԍ����Y����sy�>Ѥ�V4�,j��Bv �M�����)��k��E���B�I�1=�����[�pP�3Y�9�s��㏗�յ]uk�X �v���wVc��qJE�Q]eu���~��n���ԃ�4=������[�}�I%V%=R!��V�'ʊ���P���Y
�w��������:�J�1@�}�^O�O�9�Ho���¹�j�e���	�������݆��P�P�������[��L��%�N�Z쬡~ZR��<���Cjkb�n>�Bp��F��>��s�0�B���z�C�@���[	ۮ/Y�|6��F�W��X��?�:P��R�F��`�)�ˠ)a��^/���9������x`O9�{�"KHv��h��<���H,�S%��U�����I��N��q�b��sm�P�%�:��pوɼ�`�E$�:��!�^�12�ŭj����]^�+�m0j��WMj�3ǧ�w彪��ъ�� B��<Y6U-YħR>W	���qC�����j��(���i����'�xO(C��I��2^����^��I�=�):�nwF+��/��[�B�?�?Wd ���W*{��+�����ձy�����։��d"�n1v�dc�����G]TNV���<'��8D�,����k(�C�U|�y9��m}H�y?�b�l�p/�D��%d(;}È�����WXɒ����&x�P�;�|��B�ٜ��qk �Ϯ1�'=�fd ��Vg�J
��=�H��	�&�L�`f�7�����+iz@���7q1� `�0�t�s��q�z��"�˩��`^.b �Kh
\�
�(�nA<d��k�ZK`�T@D��H�❃�
�F�)��*kAk<Eh{m�p0�Sf���{Ōm��� ����҅���$���тp|�(ogp�\�Pv�@з X6��&���X5�ީz�V��R8pT� ��g�ߺ�?��t
7�&����̆k\�50����͐�X��Fŏu�]�$U$#�1��X��>�.��]��^r����Nԁ�lmY��u�ip��۟������O���P6�X9��
��4�#N��
��P�`k����eR��f�/�Ӡ^��J��=���g�]\K�� ������hZ{��A�/�� �����~K�3a@�@�d�G�s椳%���� 
 �5���L�w�����������+�堖~�CE]�	����h���"�e<r# ڇf��!���d�&<��{.��_u�,��E��}΅�>�̕c��;�9�=<�R_K)�-ۍ	Cg�<�ik�֋���I-��x�45��u��^1QR�A�(�Z�S�*�ŝ��L�@ф��#��C|��GH`';��]̵�/8�8�Y���f�W�[�i���7��q ���ٞ��RY�-1�\�,�ۮ����Ѕ�ř�"����=WQ��/L��1�-�:*�ʗ�� G�A�}`���ʊ`\$u��A�����؛/!l$bT"��t6'�V��F�o����4؞��C�h?�ڷ�%"+H�n���sP�ea���h�����,�ᒐ�)eF���Z�D��_q�0�r<�V� �k���,w(d��V�ϥ�Eà��Y�\$�pg���-4xy%��q�T��~+W{��x�9�\0|���N��6��x�,]�WT���|CX�5�@�}^��Y�y�Cst��x��?f��&�7]G!��1���ĥ��<�K�{)]�-�(�GE�:c��m���D�ÏԅP�33�<�&��tߐoJj�Cm��{[�=��:K��a���p����[�s�PÅWǲ.Ԉt��f���������d[g��LG]�K��3ўd?T�&$yO8itw��a��s�0M���ઇ͇�h��)�!>��@U��A}=��Y5�}�ݽ�v�����\М
�K@��H��3t����(��ۂ�����>�����n�z`���J*f{Ɓ`���R�V�s+���Ɇhq��3��pi@�J#ч�QW-�л��m[�0*=C���Q�V*͘UA�&���f	Ǘ}e�H�M���*P���酛�*�����%��ԕZ�2�򗀈���Y���NF��4?4�5;�� +�nu�sC'��6s����O�/���=�w؉m&X �ʂ��є���F�!Y�X��M�W��Ej[l�Ģ}@}"5�GK|�kI���C�"%;pJ0��9�������s�v�Ua�P"��,y�+Þ�������x���Y����P�˜t^�"ġD�}�%gf�3�j�+�E��3��z�8K^�Q}X�b����t_Ӛ!OE����>��u���(��$�|
/z~�X���W� �'�FNg��`�D�h���n�$?�HM�*���ksڑrZ������գ�ճ�)����޺�e�!]�3��P��r#�%�}���� F��~��gS���۫F��~nY��y����2s�df��w�[��/^kЂ1.�����Ɨ�(K�:9'�&#�?�	�-N�l��1������$.��3��T�*zs���[^ǿ7,�75*��%;����(���������^��s>�t��~�}��ut�P��>|��F2*	K���8��������OY�ː	H��h�p[Ե3�N�2@�[��� �|/E����.�����\eW:~�CFnH���Dzd i�X]�bJ�*oW�ebP��YJ�|�I�B:�SX-�[)����Z{:V��}4�X�c���=/o�n/(̧���Sy����돳��G���>��?�ׂ�y��aw�R�#���K%�6^�wT�>H�2>מ�k��q�7�~}Z�&��ٔ%�H�aM&a�xR_/�DmL�TP�����h)�U_F������#�T�7�=� /r}4^`m>��F���:,kk��֨�j`��jP���*\9W�h��2��L>�]�,Rc���>h@�5�D9���<�%op������P-5��s�Ѕt�n�����J��W]7q��6J���<%�n4�t�4}�C��̩s�V���$��"P=X�0:v�$�%�#c/"+�+�G�d�Ä�7w��l��,�&x��+"�api8V�}e��%��8=$�ګ>+5���^��I��D��j濍o�����������0Z�\��ߊ
����\U�h�6�>���̰����dw��C�p7�͏�<P5{�@�d�f��$�)���9%�⴬lOGܘ��@�٤c3Y'j�XCz����~�G�o2`^�ƫ�����::~��߼���EA{q����=	��I�^k�40�
d75��+%��NO���n҉�t3T��R&G8o���W��P��ml�G�"ċ��qw�cε���p�?��_֕���B�Ȳv0���;:2�X�UĖc�U֦N8��
�g[C�[.��ձt-�����_�44�M��P���$z�����#�DvYU����.. �c�2-�7 p�)�F58M�H��<�Ӛ��
m�f`z�� r���p]�7�2�:#�)����B�ˉ�w�!�Bu������F,�=wN/)j՞��ϰ�m�M�tz�P�2S���7���
9S���=��^hY~���q�#�!6W\��}�x�g�r6�l[fΎR	���Y������x�8�8c�����"�y�w�!�� ���*�7��I��S}����ĴyJ*�)��]��Vf?`D�w�3Wz��B�75��ws���^�\qʯ����g�����A���D�H�.�Z����O�P��9��	�_!^U�U�"I��񡅠D���$����搶y�Z���/;��jg݊I�pʲ��z��n�fv�~�6�oR(��HAx�4 å�����jz�����/J3�
�z��=�o��Ţ�>�
��B��.:��6�#�|SG�#��"��5��3��4xB٘���uBP�K����$�\i�z����1YinPN�������vj�'}p�h�i�ձ�)��C��ܳ����|�Sn�\sw�8����Ϣts���U�f=�m�?��pE؞��s\7�g�5T������'&}h��a�ᛅ豓{^fE�Pz�!|
)U���������/�͠��ՉF�Xr�?l�l�S,c6��9��rj�M\�$#�ں��&�ߜ�^�q�L�m@1�Q95�{l�S��0R�~��&�r+��k�lcVC�����_KGq���hq
�0