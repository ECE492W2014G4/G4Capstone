��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|�&���ڴzk^�2�t�tC��)�/���KL:�kD3���1Y,�d1	��Rv���)�g#��5�fŽâA�|Z^���,~t
��/�1����,�ơ��:y��q��u��f���c� Q��:oe��ɬH�3UH�vF���=f�r�:��dї��;jT|��C����C��7�]�x��vN2�9����]��ɬ������x�og����;�έ�u��C�&��0��qN�RG��0��R �	!���런K����9�h�I-��Ƒ��x1��],I���!٢�H������ٛ��R�O�X�-qi�>b<sKP���ZQ�{V�[*�~8��;~B��֎Š5Ȯ;��m�����x%̗o�^�4O�H9���� �����A��6�^�Op(ΣOjϹd��r���0�:��p�K@�++*�"1��} EZYP�����? ��G��-��x��G|?��e���&(3#��%���sc3L>�yW��0nꬍ����,�s��ɛif����u|��4E��*���ŀ��;�[�
}�:09}�
��d�#f��R�I��^���,���N1��l��u(�G�_���\\	��i�����@/�K��Amѷ�M<�жX��?m��ޮ>���o_�<<}7��[�����A��E�	N��ߟ��V�0�0�<;��/�Y{�W�,�Q�]e"=�p����L?I.�ģ�x��%l*�ȸӃϺ��@�(�y��O̦����J�Hi��+�J�i;Z�-)�E�%h�����{��1)a\a�9�$�Ă���D�:�D�sz�~�L��P%�Zt�?��ǲPS,�]�FY$�56���A��P�S5���iل���N��E�B�� �-KJ���5�>��]Knק���)Q��?���&��Xs]���2��A������EX(�C�G��^�m�jZ��®�;�,bl���Mշ�fr{���8�s;��|2��b���2yZ'��g��E�v�ͷ�{ś���vU?Y��A+�w�O����=z�͟4tZ�. ��\��P:D�_8���1�|t#Ji��-{��_�K��@z;�9�B�(qY$k��9dÉ��v��&>����M
���#��6lo�-�����w6��r�K��UC��p��!��K7F��H�qP�5�"ºh���7ȕ�媃�u��x��t{�~t)�U#-B�p�θ	6�!y�����mU<<��E��QO���M��G
��'V͸���@9�h-W�f8D1�]��!�<HSMJ��*Xُ|��� �&^�J�VK9��8���&z><V�N^2�A�Y�D�v�љYz�E����f���q�ޑ��H������~������,1 ��{�hs�f�'�uj�f�i�����~�����e��r��P���4��@XLOo��t&�
b(i�L�/�ȩQc-�	fhZ�%M�S�d�=W5n��.�"�g�M�~��M����מ����j�xG�j-��e��ΡOH�Ҥ�y���Ʌ�7W'rx�B(_�T��Q��?KΗ�������TĨ?4�h�V٩_}��B�oLsPP�0���oQ�i�Kx�eU���:<��} ��d�W����j�P��L`��)���|V��a��}�5nA� 7I��eE�1SZ	mEi!��M�o�T-�Ű3���m�/��b���v��{'��w�L��e�3�I����Y�N7c��TIk����~�ӅSb�������}��;T�ՉCg80��>XJ_EuY�@vާ�QBS1�Cit��O��L�L�5��J��}aM㦘�W��ޞ�T�3��F�=U����|j���e����T�9��<6��}��"M+�i���]J���
hɮ�(c�.��y\Z�z4`��xi���}��?Q�R116B��/i4�;)~$�ϰ�y}���8@�3��Xc ���ǅ���M�+�:�b�W]!��7���-� ,�pG3��&>���Yk�����nQM���ʏ��VlY�>�U����U����d�nv(��2Ly�ȐF�E�O9,P��$t��=$lA����!C�>b�>Y__
۸��a��Ks�te��ړo4ȧ/h[����Jr/Q��޴���u��T��ܒD_P�樇��laE{�Xk	9O[ЮkP�m��7�/4�����k�Sa-� ��<iQө�J9+ڐ�?�����h0Lڕ�ꮾ@��?8VF��4�I�P�[R�&xפ'ܒC}���p���v�؛t>���9�K3FZ=Z��'�[�ɯp�m���b�9������]�����F���^�'T#��nM�	h@F�;�~l9���(֠[�ȕ�ږW���虨����>QM�N�ʚЈf<�f����-7l�Y�ܾ�@i^�u;�||���Y��֊���\�͹�0�97��_�'g$�(���TQ�O�i!7�4�0�׆�jV�f(~�Q�P�	��Y���y���l5�VM�(�
�����r�@�|Xt��2 SҐ���'���c\��s;��PX�u���M����7����#�fbq���b��'�G�aq�y���ʁ��']�?�ɟ��-|�^t���Z ҈�$!�Č�
�3�
K��Iu
��Y9�Hq|�\����3X<F)݆����e'8�=��ط���X�P~ځY+M ��<��ΕD���� ��	����?A��!��|�p:M�7C	Ȩ?|�@�+�N�y�R*DFu��<{+��P9��W����8�h�ki�Ο�)|���2�P��ui"�5j4��w����g��7���q��x1���E�f�Ęw~iY�'fiQ�*c�58���l��e���&hC����a�����V!���T�-��� ����>�+W��c�A�L�j��h�P�{��/E��Ug�p:����=5P�)QJ0�0'*���a�53T�Ƭ���Vr)�,�W�a��YI8��&u��Jt��T���\�8\౷�h���4(���Y�g�;���޾O�ؼ(��֤}�:�1�OK�1;c9/o� ������v+/f��BU�:���-|cv!у6�]kQ	��q��
�X��a ��e��.��`�g����4�=�A�m0��e�)�w��	a��P�g��uY\�Ҙ�L:�Q1���`�OZ��ۻ}��V�,N"LWj�(S���5�Llm�N���T�mM�ľ���+c�`�p5�5�~$)u� ��"op���/�{��X]��G!�3��K�ഺVc;�f0��A��b<&ڬ�+���$�U�4
��oX1M3)�<L�rِ��a�sb�[���Ws �m�(:����C&���	O�+<�`Wi@��cGڶ�X�b�����4�V#jr���s�N*�.[p�'R�v�`9��I��v���q�H�n�X����%q�y0d�����ڪ���F/s������b��$���!�$^a,�݌ܜ�CZ�Jl!'��+`4�{���}������6��Jd�8��+�	�`) T��K���~.�bg�s[J�탯�H�0�,ϭ�
����:~X��n��r9'�#daŌ�. NC��)�q5:��h�v�ϙqV��P�A�o����^��f��J�^?\���bR"N+��
��"�lM	OOyr�FmdG4��3S1�O �R3b�<Q*�'\5��Xu�o`����ΰ����>wl4G 
�yO	ީ�-��s�@�;p���j���e� �5F�����F�HF,��X�)�D��\�?�=�q�cj�c&^��my;�S��f��_#O�)
P(��>ՁVI�ɻM�Ո��~j?).���c�uDzL.Q}�:9�M�OȘ�*�݉<8i
+.�X�߱fD�fM-^-���FN"k� q����3�w�{>�@����-����!��~NǛoΕYt�m�*��Tz��-˭���%2�Y3�«m��b֤���o
�@��!���7�9X+�:댩�&qh��soQ�I���	Ժ�	2
���e`Ŗ�DR�^�AU�W����tN�ă�biZIb+(p�r�X�}q;���L��"�S�<X��C>U2�~���Cr��[>��;ڶ��	޲b>���T��|j���p4$��4|���qF��\��aʐ�q4�K2M�M�yn��[S��x{|ǝ�pn�o̵�;��	Lh�
	�?�i�������`ْ��'"�訾.~�~�8P���	��0R4�j �hg8J�e�h� ��A�e���)���5�9�g7Z���*��\Ǯ2U��>pП�Lp[�tfyusuv�[���_�붰3)��x+92��wu�ς2Q����h�:M��%�aN)��U	�{�(>��5�}u������|e�� (E���.��.���ҕz|���9}��T}#������Ċ�$_���Ѳ\?*ߑ��0�[w壗�Q�xZ˝έ���l����t��Q�j.�����T kD&�������h�Td`g����R���݇��u��:Z��@�^��0Up��7�7���O�X���򻥠�YA����jɭx�kZ��ec�ɢY��,� -ے�U�#�pD�q
��)&VO	�2��C���u��(Ɯs����1���_8�6�&_Ưɤ|
|2����3����E�8�Xg^0&���@A���/�;�q�)��<wdȮ��Jq����c.��z�]���R.�1��]��p��Ь�u��(R(���1>2`f�:3��ZTz��R	T���*E��62�qD�Ȁ�}�;8��l��͇�ƫ���i�"��BY"58e���e"*�;���Ox�_&��i�5+��*��%^Je�l�ƣ̵����_�T�-C��Y�յ�y6���7iG���Zԙ�f"�v�p��"��ǟ�B�2'�xCL#���0�mO�0� ���o\�=;�D��z��k}���d} �:�$�e-��x�P���kr�@�>:�ΝRJ����sR�#�H���C�v��-<��Vܐ[�/���*�$,<��Ğ�D�&�
,p�ܞ��k��e�3�D�p�T���4���d$<o3�Jw��VƗ���lJ�հ�C�$z�����S�`j������}sjS��zX�����1��1BMΗuy
AZ�Y0\��o���k.�8a&�O-���e��=�R�T����%���U�:�h��$����Ð�`|8����IDW�g�h}����c5ưL��3���j㖣����z�T�"󂡂�L����>�m�����\����!� ��Men�n?��.�g���P	yXQ\="�j�;�za�����\��bQn�ƿ�,�����IO��C��zr� ��'_���:���a��B8�K���衐|9���:S��|��� EU�srd�o���;���H\"&o�(-��0���d�Ŕ`5A�E��W�T�0'<�\^'��nA��>��S0�re|�<��ȃ�ޫ
��^��ĺ����S��-��[C'�Ё&�����)��^ip
X�l#�b�V�,SK <.�8f~�Y�3b9Ũ��S3���3=��_�C�����ǆ
�c$h0o����6�R�E}j}�����Fį�߬���^:���,E�n�_}Q1ir��I���ɤ��+�RLq��:���L~Iǻ��P5S%m�ܠ4����X��M�4ŗw,ׂK8c���&�
�yy�)��߄��J[�=�<���<�m���;*B��PʄpJy��������_����xf��:�˘ܱ/��6��j�nv��5��Ȍmf]�������Q�����$�P�f�am�U��8��0��.��K���~� ���&L�^"���'f���]��+)�	h���մZ���p@��>���en�s=yKi����u��NqͻTM�&��nR� �R�H���k&����Hv�v� �V�b���m�*s�Qj�_��l����c�N���<��LS���@��q�g���b��f��U`{�0�D��Y���L�}/�I�E�&�_�]���!��[L����P -�;.�T+����p/=9�q��a̚yʲZ�-T�DH���1~E�h�ι�E6.Ye\����'����;�Z����и��Q/B��sϖ/�N[�R{�d�e�<��cb�x( S%M�]s���`��^J�^s��T<�?AC�ђ[>�@���=�q;����x�nf