��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]
�x����Vu\�P��Xz����z��g���F��[�W���b�T4�n�^�[��`厸n2���@�-��y����1W��T��j3����1��1�W!Dy���z$+�ۚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P��v�"<ߞ��&'��k%P碶�R�ӣ�sĞ������FY&<��� H���+�S���A1�JEI��NRcΩ��wNp�J00!��Gk�B��Ճ	ID���_�N���1�4!
Hiߙ�+�!�Y�?�MQh�A3�Ӯ�*��%������E��,�wd���:���	J�c���IV�dΑX��tJG���?��Qk�r�t�q�7Ⱥd��M�T�"64�QREs�I�W�D�D�JP�y�tR���>ͺ���[X�	�}٠�W�:��A� �݄�,�4@�{ս�K{�E��D�6�e�s?U�f䝲����E����$&�$���0�B���KG��B,� �J�n:�@_�/�R7LPC��`RD���0eJ4�Ԣ��Pl_Gr}���.��u�(a�=�5���sc�#�sS�t�oZy�JΔ�[=X�o7�I2g	�@eba��S�BW��������e�֮��$C���~C-�ם�Qث�(>5&�4��h?�2�[[V�O�j�&���Z-��Eq��Xz���������7B�w6M�8��W��LO�y�y�%���HQOӯ���ų�xW�H!.IHк�n�pc��P��X��=�_���r�� ���
�)�	z�I9L4�T"̗��V;�����O,���D��>d߱	Q�JN����?e�i�Y���m�߼�ZlV~�>ޯ�Iv�L��/A��y� ��ؗ�֜à!m�͉Zh�`��}���u�܏���!^�`:$����/�!4f�=;0j+z$N<KC�CK�'�9�%��r{��y�;]� ����I�7鼱1��2fh�ح�?����(=2����v�%���O�&��ɘ�F�X�q��u�Vo����Y�G�9x1-Qxo��%Q h >K
sW9?�J Ao�O`�q1-0M��yR���+�&E������(f�LhlQ�o/�kS_[�TÒz�_��j=����D��Zi}�wp^1���K�lJV䬚�t�޶|�%|�͞
UfO��o�0[����Z�=���#� a ȶa0�`�B��ɮ�G�P@�Ø+����2�-K�t N��qv����7��p�/[?eK�3�ɏW��A1h*A�R����<�0B��ջ,�b�=�Y�
-�a`�2����r�"��1FDz��h���լywxW�@jwm���,����+[N��d�D���>@���,�J/@:��S�9�ƌ��(v��K���y$ �R
Ժ9��m�z)��V̒��u��L��>o��u�mU?_�ڝ�gc2�N�,�*L}oѦ`)�3<h~�(�{�x��eL�Nj_"˺lڱ���D���E�!�t����U�A>z�����v�r�����������'�}V��a&�%�z�R�l�=Z���%=}{*�[$N��Mr'L�B<�V�J?�D��Y��z���tjt� �Dlf�Sj|M���L�6��՘���Y����=��Or#0�a�`ŕ��Rq����[�EM�D�q��b���v���H��;^�ہ�����8��	�?�lt7�O[x=�t���]B�]�yU��*V��p������:	��, �Q�I?�z�l��Ɨ0 BXN���GG�^��H��~O�PQ~�5FU���;��ٖ��l ��D���ё�ZM�p1�A�0�U��}jƳ��Жv��qYo��8��L�����������(/ٞ �E����1m;u�_�����E���ţ�[D�v�m@�?��t�J��T��9,���N\[��~�W#�o~�scی���KR䃦��]��%j��#���&��k �y\����	���.Q_7��X�9Q2��+������I����G*��1�q��P�8>-4V���z�%7(V�$B&R�]?��%���U��?��izʽwt֎@@�ԿZ�HgS.�?�+���Ж���_���bI:¤ݓ�-/�A)�[/�Ǻ�(�Q��- ��KF�j��LBf�I��V2u|�	��sۊW9��y����^/yX'�m�{����H�{��_�~6>�YQ}�l�y�}z��"��)%Fk��.�~=�?��$w�x!hv^���"�tD�<brR�Pp%�Y����1]j��W�<����&���Bh��K�|pw��
��'�����ƻQpm�������A��꾷~���X�U�~�"W��Yu�]���.��-x�������C��%}4�!�>�kz��TFT�#�p��YY�N�
�f��͖d�ѩ�cۈ	"ߟ�^��+�V�ɳ��o�"����\��~��\�`AT^��)���'d EL�g��fm4��?��'��G}�p�H8\�afe�K�V{R���������.��"f�t���"�vH+S�#��b O0Oٌ���/�\�֎@�Nl�k�	���py��zfF#'`�lJ� J�;�9i��%4��67z�}A^�d,�1w0lev���չ�6�==���f��R�op� �ҿ�|0���6Č���ޯ�l��Fu�/�o+���#<h��j3�o�.��f��*:H~m��q�2�x=D ����[-��U{g�e�Lꃏ?<��2�y�Tz����j��T��Hv��_���=�h�/��}0��.}ZD�u��f�i�D2]��)��K?�o�Jl��:�=��eO"&��K�[w�#��!�dt��x����/�+��w���దȥ�C'�ԧa��t:�Cmf	ۥ�Ju���-�<���Ϸ:��$���A�M�S����l���}'�8uК����Lh��H��[�`8-���9��y�%,�E�b��LFG����6yyF� ʜq �p1�?��Ha���>}Z���ϊ#%e�U-)O��@��	'V]dy�n�G]�^�D�;�ɞ��b��b��og[=�J�C"�yx��b�ۅY�76!�pYIw�������R�\�{q󭯵ɬ��	'M2��O��V���n6������a��H�<�(
i�=�y{��XbwjБ������T���/�u֥#�{l9���Ã���`Ӝ��5$^�j��ͮC���b.��TC�֠��S���/�oǑ0�ς�K��+���#g���=�!�i]C���_ڲL�@94��4�@�}eJ&ܿ�����e��! M�A�t�^M�zW���kNw��E7^]�����v0��"�w�9�*��3�$�hy�ui��E��P@��0*� y��uk*���p}zTe�AC%���9!̃���ģ������{[*��0�	��=Z�� '��y��\��*�'�ϴ!��y�Ë#y�X�?�Xk��H�G�d�����	��g`p�)e��I��J�,���Ä]��}F#��h��ңߋ��<;F�FK�Smz�ԧ�+6��l{=QA�]���:L�����Ԩ*�?��Q���%nm rի!�<V�T��P�2U
��z��JTN*#��ALQGR�I0�f�8~�vLS$��otG�(Ү~ؕ�2}���X*rNQ�(e��g�[�9kP�a�'q
�VJ=gu(��	Z�O�u�l�����՜�=W���c�(�L�`���ع?���� �T�j
c"[X�:��� ϭ/��|�����R���Oߏ�-;��O#�� }��r9h<ZU~�f�pizAڀ�V�uUOpB��׉�$�Ok"��%�S73QWL&�b:�����i�����.
�	| i(4� K@ݪ1T���E�P��ޗ�kɑ\ΪA^�~m#X�.b��ax˿��gԮ��8�1�$cL����l^�:���|�C�����!�y$��jE�9W��H�$�z�k�*Lc�0r����������ub�5�j1��0�=��%X�2��b����Oq?�(��,�]�3���$b�l����]:�W�ΚN-{����<��\	�^'���%�Ρ��x(�<-jx�Ne�g���~y~9�Q%��[�T�5�yf��3���y"�pws6�@Â�f	Tu��5�cEn��+��*�;�e�1`N�	[ĭ��c����n���?�4��"�ç:���Fl�'L��.�>eTa!R�1-���e_�'fŇ���ظ9��b�R&�3> �7��S��CX?��-�ju��ls&���8i��W���:+�nwUք�j��<���H*�F����J�f��E(�ξCU��_�h-u�h��.ֽ�î���
}OA�d�L.�Q��t�|a����96
3�S.��鷳ծ������{�&��-��Gy�G
���yþA����U4��-r"���]%�����	�:d�W��xK9�������Q*�jR��Y����*�����^H���m>b�!,�ǌ9�H�s~l�Q+p��O�������|3N�y}�I����պ���jN�l�������$zޛ��H`�mذ�@�g�H��]g|�#CU��|=�f���9����-et����8#\�
j���t�V�t���A`�Q����QE��%矆������0����R+���w�v� {��I)s+�ː��~T8��zd
|:T~�jƊ	ݳ�ϩ�5(��ї�;1G�+�J���Gz#T��3M�&t jqGl���.�c�˓_�N,;x\͐lT���s���G�^�ǙE�@*N0�0H܉�@�OE"}�UȨ�/(�:����5��5!��Dӵ�w1 �.�9�F�@�^��(�W,�U���U�9��/�z�d	�W΀�蒱B<	fEmXMqm��%�a����rϷ>����@�h�+k�n�-q	ei�����|:1�?��$a"����_�,0��p��x��js�2�DF������b�'
8qK�;��^��f���= 4x�����&ؗ�G�0�u,"4��k���x����f3�29�9��%R�o�"�?�� `���������V�=Ile��λ��k�����*�lU��-pR�n)��.�ag['e�z9$
U�wڛ}�z1��3F��Z�q�����@.�X4�_u@3���̗F2FȎ�.n1�o}�t�M��p��.�1�y� 踫���v��BY{��Њ��E}�g�(�ğ�6�B�˂Ɔ`�K�)�%�'/(�����!�UrF��˳:���G9�r�~קtQ�u2�n4����ol�ᬝ��|bR���F���4��]�ԝli���E׎�J�<ח�]~��ޚ�ڽ�84����*�\1�gp{�ȉ[��;�?|��69(S���<��K2��@Zd���jg� ȸ�T
0� ^�Y�9���I6����d��Q�8H)BfuH� �0�����jUCB� eEz�������Q�N5+Zo�9����oC:�RT�����m��0����~�7ڛd9���0N�!��p�x���0^�W޴j_.�
j��#6ֲG:A{L9�	� ?��5�G͞|��H�$1�((�y��uAy��[�f@>�����X4�Z+~Jzu�L��g���rf�� �M?=��,���6֤hu'��&�f�ފŃ�d�?�6:o\��X�vS��o���"`����a��'�۫�4+j��[Ay=��Y���,_@�
�Fz�G�CO^�����:���,�O�үP��8�S+��7�N�=�&q���6�	���<� EF�J�I9��4���n���OZ�L���!�:��!�P�Kj ܈�N&��s&#��vM/�|"T|��;�ܵ`���|X�?�w>{R��i|��3��)9y�5�}��x��y����/��)`ধ�?��`�B3��	3�g��	�@i����m7kp{gV���}pKL-�t�!��^|t0����2��yzc~�1���?LN3C��.f���|�i��ݪ�¢�����+fW�@<F����ʾ��@�'�ԇ��I�qɤ&�z����Ὅ��(�>�Ҫ��;��r���e�� ��u}�d��s!]�,��`\3��_�����`�[x?���+�o'$����k�L���Tw�5\��A�'Y-��~���Y�C�}6�HE{d�ٲ��jYZ���#yoa�:�
W��S{9�T,�@��c��hJHu*=��jH��0kV��k.��[�D�Cb]��5��ߞ�����u+LU(��J�#�r����_�(��ϦV�)'+m�>Եs@A&o-�X `d�_���i�ۄ@
HF�o\l:�;{����1�(�|���~�&U�𜁸���f|0�eȢ.p�L&�Ȳ��x�#L��02�e�ͼ5%��2�ʫ�+�{j�h��<g�6M ��eC�<�kB\���N����]����s�&='G;���/������3��҆�h��ɝm��d7�wW+3�`�<c��y�0�dN�P�g�N�zE΅T���9n�ψ�Ƶ5o]�V���#��;�[P}��Rx[�� ҳ�Z.��a����h�#�+/���	V�5 ٜ5(��1}d�_)�y����E�w;���M����\Ӷ��q�H����V�f�u����G�aȦ�I_rY�9�'�I�xi��N�����D����A��Q_�P;N�eܐ�	�!]����)(�q�i���CPvi<Bf�M�Q��J�4�~�Ql����[ޖ����?:�M(߰}3�4O�F��s�Om��s���1�	�K�o�y��u&��S`������B5;�Yo�6���~���#E����1�����9
I�B�Jg���RBb]o��OXx�Fo��o r�%����8K�<:��4�h�1#j��e%��&%��	(ift����S� >����%I�4�y2��;�q(k��W�U���-��t��x-V|��f=p7�U�p�C�\�����yS�J�|m�����E���e8ąY7���L��k;x�Ų|>��/�Nï��0�zA�!z:�_"��BI��D}W�2��.���[�{@s�oK�Q���ӀִM"LT��&��,��gee�%�Sl[=����ػ����A���{C����`�D�r��S�!�ݡ6ӗ�бX�S���~Vۊ�4235���5r;y�24p��7�_S�a�vܘ�0�nJ<�o���5~-Up���E�Xߚl��ĵ�{Ad�����B�� Y%�O(���H��7�B�8��������c2A�� �M�}���=�A�+Y<H�UR9g_�|}����E�ZX�\�u�6�o�����gV9M9%�#��_����T����^.�%
'z�r�EJ���L���|xH����@��d�R:	�كй.J����*��Jsj�r2C5���v%��Ԙy4^�v(S@�F�P�E�'j��?Ǫ�&k��gp�Vs���x�ϻ�!���,���	Y֌�Ϯ,d�Od"��~=��	��"a�gpy���1�$�� ���{�:*���m�w��e��:��<J�N���\��*v s�U�~���� c ~�~��v���HI�<���h22�rǻ�g��3��8�BMqv���
{׌��8؟w�+!Z��<zx�8���@�ʖc3c���g�OQ����ě*�A�E������
��B���yl���'����i����'(AQ������߲tJw ��U�m_��¥.b�����=�T�t�A�od�\:yMݭ,E�,tG<�/���+��SD�<34����1=I������	�Gm|��2���~���R�f���&}���x#�G��U-�?aiu���Fg�r0$�C� �2�ْ���"���f��xKM��4@��c�-3�X�FB�<b�D��^�����A�X���h�Ĳ$Pg"E �ئ��A��&z����:�48��P&������Ѱ%�B��7H�f��کr�����K�'���
Ķ"S�au�wY�;d��G#i@�`-&\�53:��z����|ȹo��U&�2I���>���1?�S�|K�m\��S�d������-_�Ȥ> 9l�HQ55.΍h�ۺ� h����IX`���*���r<����͝aZ@�<<x�K�$1b�5s�)o*����QF�|�n�6�׹��V�V�Gj矴889
�ݲ,x���C^��4|te.8�>p��;yg�Ћ��d�
_<b64AJh׵�k��[;FxКf%����G qS�������&3�7��H�C�_ch�f��0<P��������o����E�}��FUro]��� �p���G䮇�S\R�� ��mCɀI��]�4uǈP�^�=�J��^�k�^v!? O���L�-b2��.��K�?[����BaØj��!������W�ۙy�b�(A-�~'L��>�n<k�g.�W�CR5�JP��|i���2���7"α'���SٌN(�?j��Q���`ˣ�n�����o�8@�\o+lE��կ��z7�������=2_�Y��e��e,Y� ��k���6��U&C� i�/����7�+�8ք���|��fz����Ј�r#��<�����X��?��B�2�ֳ�(�3O+�!�4��$L����9�
���C�
�BdsC,!!�������}�uy'��>?|��Q3����Y��4�Il����F]b���Ȕ\@YZ���uf6�!�Q�B=J����Q�Yc�J;��V�]c�D�#����l�f��������Rr�0�?�R�߾߂Du��2���A��S����6���CM3O�-'`�*	��gF���lBM�q����u���/.�Ҫ����L��L#�<�T0�9O�[j��kې�;=�����!������d�F�Cx�>Fxv�L ����`}G zlh��~+�I�!�d��{��k+�gl�6��a�X����h�|�5k�i��h����Y���x��F����p5�`<�%I���奪�N!��^ʥ�vs��< 	`���K����y6wn.?��s!��K�@ʹ�R�>VbN�W�z"B.����i���,W=��a������1Í�E�����ߚ4������ܯ��J��M�On�I�BX��Л�%L�=NZfF��ȶ�ga�4�~�0�Y{S�c���\����8��P��<%x���g����(��90Q�Y ?f�ەʾ
��G<^���o���4[�cz�� 尮��Ar��4�$!��S4��(��2��u@���!1�%u�y�u�x�Ȥ� [�3u��k���cʏA5z ^�sO����Tg�7����38��uD(��+@�f�.��r(�Q�|��y�<3�!���k�9 F��40SH�*��[��캓���]@P�$|m慗KS�Z��6�?��>�j�1o�9����м����S<�>
����c�_�5j}X�h(>Ck���)�%�]l��T���%��JPl(-�2x��֝r*f��9����u��0)�j��3�M�f��Hyٔ;������(���"�tV�@1Z�q��}�K�7��"k�Y]1���[6�K��v��d��p�Ce�*,`dx@�_l6��\IɁkʚ��>�|���WZ^�S��8��&��W�o3��?K�ك��1C"T��ՅN\�B���c#�E����f�%Ϡ���dB�6���+kt���e��x��u�A����9Y�NÓ�1�8$�o�(ib,��hgwB����$#?���O[ԤN~�!�
4��:���%|Ko�KHZEmDD���T#qD���3m�U���}{l�7��.O���k�H#�y�F�sC�QYř�_�k��F�6���� 	�n�dR��J�U߾�Q�D���ZF�?��x鍚��y�6/�lAg�>��;��bWXe�L����f9}#��.(:|i�����Z�6��Q��g��WICDkb¼����<�6t�FcN��$*[���S�y�H�*�u^��z�����C���"(�I�@���b �a���y��Gթ�+�/����!VU�a�
��"�O���m^����NЁ��s�d+?�g8y�UT��Gp�ZW۳��qU؈�[	�/3�gS���S-��m����������N0�U�TB�;EL�c`�� ��61`��Ӡ���O�}o�
��?XvV��V���`~���؄=)�ln(=��3N��*_T��*����ϛ��	��A���̚��;���&n�(����zL$]@����[<�d�r�az(�jܞJ�&��j�E|8���}QPF���
'��f�*���:aNz/���)��C�S��a]���̤�[��z����NL8�f�׿��|#q�qm��,ì �����RSŶ]�0������~��>\��l�&;olE0�}4��O�4�;��zo��E���`��^����ȁ)A-ޖˣ�mT��b��k-J̘*7XJ:�u��Y��=G%�v�\cS~���mU%E6#�E(!`��@s�.Us����Y�������.�җO~Ц+��O����$aܨ�"p��tR�5=b�վ��d���P(ܥ��pYj'��)<�t����vF,���hk�n�F&�1�9�j�� �!�dz����=\��˻ܞ�7��L���R[�:�wZop����@��}��;܍��Q$�����.u���<3V]�*� ���Df�����[fow�8d�`� �k'�}X¸�+�D��|�]9���BX��R�����mU�_�G�v�������Z��u9��8�b�]��H%��L��0��{@�N��U��(J=c�����q�*c�����0G���s(��pD@R����<P&tc3ꚼ�+'TT㈆G����W@��UH��%���w�z��m����i�ې�|hQh_qI�Є�9Ÿ�^�L����׌5�Svv�x���E���]NH� �c�����s,�~��e���e 2>;x���#�f�JA1��Ӈ�ɟ�*~R���`31��$��ge�AtZ0��Blv�uYA�BU��[aAA\aP�[)�D�yf|v�����=��4��+�?.�N���HyŅ�f���DΪAOO�E����Ck!PQQếpj�z�ţ�i��T���[�����5�1�6&�¼��GIf�Ǭ'$g�B��FR���5�P�~�a�Q�|�����.��
̹��پ��}��BAͥ�P���5/!��UQs��Ҏ���j����W��8j��ى��o�T���tf��g�Y6��}���ˣXuҡ�ֈ츋�RW�J�~m��ԎNq����y�M��q~�^D-�K��%w�na�"�_�IGj�^���~�a���m( �"=X�����F�?OE�m�w5+��	I��_ۙ:��꼚V�J�'|��YdO�UaB�n(p��M6l�3J�muD�Z�c�%;ס1�����70=98(;3WLp���xNJ�xH�)3sQ�_���*���>D� �Ni@�Ē@³�[���<�?�.h�j-�u�O0j�5,���ŵ�Zs<�(�~ \vS���6k	���	M�0&������@z������qQ�1��#��s�@���'�!
U�4|�+ͷz���^�	�1�f��L U�{A	�=;�ٓ�����P5dNzŰ�j��ᴦ���*$�z({~���ӣ��W��%��:���S."`-+��yr߰�=&o�B=��k軮��O�k����m�6�Q7�O�X	'N����fxX�=o��n+M-<�8��R��2J�-ķ1�_�P|�h��jͲC� m9-�mb�����
�Ό��P�Iu_��F}O!���pP��t�L9�jO����p���I�]@��0 [
$��hV�����}��|�;�եWm
�9�V�1x]3�w�����j0!��p�PQ(��u��@�*�}}��EP�[}׏F�f)�M���j���p��h����!f:�]��$i,�B�	�g�|�%��/�F�{�y��ʯ{5k��#f����^a��C*Ot-;��[r'sĀѪ���ت4#3��u��F��Ni�i��N�n����NA;�f$����6�H��C�	f\�Q�c��Ъb�tcc��1س���"�28�:&5�<�	�bzF=4J���$*���~�z �� ߿�ls+�Z��W��
mg��(�/f���K��g���e�U�)1��B�_���Et-�Vlj�dd���	���Q��?�AyQê~��ϥ�/0WmF'S#*��"Ʒ�	�Ye7��EX��0��]i������<T�	�k�:����H1���_�+���f	��?�o�D �?��9"��E1�_���1�N�@�?�ܝ���g8C-ژ×ܘ��T�g1��oz�;�`T#��M�҅��i�������jͿ�G��������~�o\�A�9s�H�2K�Bg�^��!A�i>pQ�P	I�au����#�J �,�?TM<lO��p��H�S�X�8����0!�xQP^+��JC5əV�@y;�9V�����l���i$�F�Y�Y��*�[G�ɡ[֦Q/N�7mw-��5)�؍��2}�.�0�]��CI��./A�N���}��� ��_�V����L-��6�y����e�3�{���6XP�QYy��`�I����'�'�P��P�����|�t A~��\��-�!Jt��u'=�"Ը�b6DZ���h]�� Q�)�f��@M�"��b�����栽�z�����:�l�jRz��}�Z�1jfc/���%1��Wu�`���9�Þ7�x{@�o�e�M*ߧMZH$�2����S̭��`�a�9e"y[�#� #���(��U�C<|W�
g�ǹ��K'~"�۹%�i���s]�l�:�b�|Q��c�p�f����U.�n�σ.�'T/�~�d��Y4���\Hc[=�a�1�O�ǂ�||�(�ڮ��#CC��#��ܡ���Mi{hκ܊������@<���3«웷�-w���,�p��<������$��UY.er��=��L���G���&N��X���:(Lm+�Ym0{4�)����<|z3\%����il:5Y�{�X着��P�40�Ov��c���/�� c�m&�5<�D�@H*��x9H`�X���@���h9Sr
��^tbMXK,b��`����M��\l���*�z��$�G>��J����� Y6i��䎽�:�����ݬ���ū�9}�oha>/��wg� nXCs�]R�N��MK�1��)�^JO�X���f����6�M�r�r�"��SF0$+��{d�:�8
�Fr:3���s,�(��{�t^l�����~ж����@�4��Sc�c�Q՝���w{�E���|�A��%�ag����'V0�Ǖs'��^yƝq�����~���
�0l<>��^�j��j�:��.D��V����(/�'��si �Z}#r�p��bꏼ�x�:����r�����Q�<~fF�_SYg��_eՁ�|�a������2BTb���G���'�wb_ek��_��r���"5l��J��yہ=l�o���?R��������p�����Rr�*4D,��Ua�}0�OixNe�^�'zbf{e���^L+����.�UZ����b*.�&�(yh<��W?�b�V�AGnSr�_�ł �z�\=lm�"�4;��;�b�9/;&��o��p#32�������������[e}���H,V�G�y8GK^9�s���8s��5����.���CQRsj�_і����-��Pz~E��R۞;�Ϋ$gm]% �@^(7��X�k�MNX{�7��~���KhRܹ0+\����W��XvB�`�l��v�s�@3m]�tލ\����ʏ�`���*Ę�V��l�&�
�1�N�b߯���K[�t�N0נ�şSy��%�h�M�ds&VJ��[��Nd��.Ֆr��o���7�5D-�?8����z��ѕM&�Xݕ��4�J�j?=0+{�o�q��"���l���7l�K�R>J��7��2.����6�<���-��Z�7�H���po��0� ms�!q�����nl�>��Z.���F�ϰ�b�#���D��C��yG	�5<U���m� *�����D��)pI��ɂ�z�X�.B�ujQ�˝��/i53 �T4�nN4�<� ��ԕI�����`��`��<���]���H�B��$��Dv�[M�H.K�yt��i���9��Z��4K��k�d���X d�(p2�	H�w�㴔��|;g'���w�3G>r�_^�mJf� �<M���2�ѱlҬ�L4C4�x$	F`GO�^*˧��!E��$��Mܿ��hK�c�D��U׼��[S��E��ⶒ�	MVVL�:��0�� ���r3�{+Y���쪰U�d鯯 ��(_0�G�D4�H��T��3�c�Q�D�{Y{1�ߦ�	7oa���gD����('��6�V�e�]� C�Ќ�+�T'i&��~)���я	豰��4ʕ@���l짪�*�Ն�'+K�r�l~ڝ���V�Cjq.��i��r+"��J
	�r�����}�j���
v�W�rR�6}$�Í�M�l`5h�E��P�F���E��Q,���7��!�'�����xW����Z��[�7֌(��m�<=|���)f�zlF$��7f����������M����!N#{���F����Z�2@��h�gRr̥�e�Z��fY�3��Dn>�llC�����u�������%��yc0vb6�(�j����mc����!S���T��ҫ�����e�Sg���q<�>'����[Q~G�VyK��v�=^$RR��3��X��zee"������}��*��=I���%qн�t��]�Ѭb�'�v����XQ��F>�BWXr�	��B3�z�(�,nQ�MRJ-F��tg���OA$F��#���J�R��������u�}�wp_�*-ϻEPf���?��B��G��zş��]q��zqA�k��8�ʩh�'C����hZ�-�N�uRAH���҉iœ�NpL�s5�1+c�B�b�ίj��`2�w+�,һIV���T�">��36_ƪ�I�k*\�N�e�d1����>k�\���� �����<A=;ƿ�ĸc<����j�V�h��7t��i��;hc�n�?3��W�s����=i*f�2=k)o���=�g"3��B���N~���.r�'?���:��F0�RP� .<_02�]�L�����>L�v���{�!�:�����휍��BkI�3�&0�MҼ�X��bݱ�jp�na U���\�ȭ6�"���k��?��jd�_������R<�_�!EH0t���>����B�c�� 0��A��E�0��7B�z�1,(��F�d�o��up:ĞZlZ�<Ov�z�Pk�`������`C����[ԭ9�k�<p6[>Q����v@��c�J+��G`obF�t�)����F`"�A�����tUl_+����Z�<�K\N����(ȿU'��@\�����d�:�TpΜ[�$m�_�*M�ʉ����L|���<�F�&TkB�����K������w��^�m���G��ۓ W�YOI��5��:>S��}���-�q��fD�Ϙ����D9����
ֆ�O�Nj�a��ӭv�!V4;� ؕfw`�R�v��CO&.<yo��X�N%��s��JG:@�;4-�i�b�uS�a����H�:��`=���U󛉄�jer��&�2���/�>1S��8�az�!�Bњ3۠�:A:�,�.������w��"��(�cCY�CQ���dF�b��኶?!�7�.���7�,��"Q�?��V:h?�xV������������'�j�pd�`A���H�!�k���(�M�5C�l�ϱ�-H�mw�gX�r��p�u+�~!�!�Ϸ�ėt�����"�PՄ�������)c��G����ieWX���;��j&��G�#e4I֤\�W6d�ۿOH��%8x̤��	<-�j��P�8٬�QF�(�3Ȯo��Ǭ�B#�`t��U�"�����v���}�=�NԆ	��7k�P�4~s��5�U ����˲�䚚��i@1�BT���A��7�a;5�b]��z�����1�WF)#�4W=M��X�z`�]�: @X�N�K·�OJƟ�3l�ߋ	I��F���)�DԂ$���D�	Y?Co�z��P�-Y��Pw��}�fL�Z�g���p�N��ߪ�{�Hg2Bqؔ��.�[�+��1p��Q�I��`�
�_�~�F>+1�����.$w_��r�� ]T�Us>diy�T��N�|`�9j��72�UU����-�f�J��Ԕ�1qe�U���&�$ 0�m�i��!ѽi~(�{GH�.c=�փ{���C�/T)x@-��d��X��#�ٸl��?��rn'Eo�N���Iȸe��
���k��� ��� ��2��ġ�"!'7ͨ	��<Թڷſ7����:�W���}�iL�Ө�R� �~�>�5=Ve>�X�+ �g�:��0�\R@[4�P�tk��8-!M�S5	9+u[�yP�r���K0��dѢ/����BcC��Aiܣ��-�����X���|�R��oMP��)md���Z!͎����=��DS�)��L,x0T��>I���6�h��J�b�N/ɋ �c���Wf]~��}x+���,v5���W��C�g ������J7��:C)�A%��Jh�3'��c�f?��/���vQ2�fsL�DM"\駻t_4�cS�0 ��,|㬴�$��5}O�n��&�I"�w��H�[��-�1�/�j�G����J�V�)h�������1gjkĹ6J�=ܣ������UQQ�
���/�	m���vwB�	~�'��F!���fI�U;2�Ĉ^��L�[ͧ͒��;�� 1�y�^}�ޚ�����.W�j�I`U�K&�#"��P�G�W9�tײ=�����"~�Sds,�|��E�(��é����b���0Z�/����l"�hW �j����iڈ��N�Oԃ"��]�4^�DˇT�ɋ$�r�:����(�M2� �F;�������%��Rx)�I�l�V/�iv3
��l��b4�DӺ��H���d�?V��Z���tJh�P�?�#���0E�I��Vfj�h�����F�9��~s@F7�Ч{����|1��?�}���K���Q+���ܼ@b��* ;|,��盙����?[®�AS���?��يȅ�@�4�Y����%�,A'�>8��%[��d��?�7s`��l����1)����	�cn�l��)1]qY�5,�p��ʒ�"mH��gf�zƣ��or+�S�XD��c�ty<��K�Y�6����#+�T�:F���	�|�b̸�փlQ�z5_Y�>&.��rh�>�cA5���7{�� ��<�?Kd�AK+.15Yy���|��9�L���{R��v�����������j��#0�ZE���ԗ�B�y�cV� �Ȋqj=(#����\<Z3�  	�鄷%DPO��V�'���gW�_
�d���Z�����6n%w(1�}�?�ɢ�<���,I�3�����X�k�����f����ӓ\���:��գ��EPKh�sńI����&�--ܼ��u�R(NJ�T��gӘ�����yTa���'�,v����Ϗ2xb٥��0ڌ����:I�c�L�2���yd(J��pQ77�ߨ��o�P/�d���P�����v��B���}y�����K��Ʈ.�J�'���B1�wz���J�����#��S���4�朧\ʚxpΪ|:�2J���9Z��7nh�����rKP����ҕe�vI3���K�3���8��A���S3�M�q4��)Kyܐ��Tҩ�D�R�՗��j'7[���t������6C�9m����K���G$/k�E�%�-ٷ����f�2�if��l��(g�� ŝi���6�����y"t5�2�U`������0l�$�����-���^�@�^�5��|6�|�S���++�+W��Y(�R�xv�oP2�&�V1�E��2-�L�vMz�535?�s�g�Y������x�O���O���y��Y�@���J����sM1Ш��[���c:y*3�`��-��g{�6K��-��־&0B��'��r�"�4J��=0��W޿WG���#B�x��3��7$�0���S�F�d�I�9xAൻ[��J��^�[</�e�L�Dt������LU�)`�^(Y��J*}�j��{If� <��a���#$[���[�� ����<3~�@�bQU�5�4#�X�iK/�Q��@'t �Hn�)�l80�z^��əX��^$T�SM� ��Jv��b�}F2�i�W�k�6��?�@ZWw[˛c�D�1�Z<ǜ��L�F('�mW�!��_�*tqy4�W��%���ͻ@�  �8JN���P